// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.13.0.56.2
// Netlist written on Tue Sep 10 11:08:38 2024
//
// Verilog Description of module top
//

module top (clk_25mhz, rx_serial, rf_in, diff_out, pwm_out, pwm_out_p, 
            pwm_out_n, led) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(37[8:11])
    input clk_25mhz;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(38[22:31])
    input rx_serial;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(39[22:31])
    input rf_in;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(40[22:27])
    output diff_out;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(41[22:30])
    output pwm_out;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(42[22:29])
    output [3:0]pwm_out_p;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(43[22:31])
    output [3:0]pwm_out_n;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(44[22:31])
    output [7:0]led;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(45[22:25])
    
    wire clk_25mhz_c /* synthesis is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(38[22:31])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(61[34:43])
    wire cic_sine_clk /* synthesis SET_AS_NETWORK=cic_sine_clk, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(78[33:45])
    
    wire GND_net, VCC_net, rx_serial_c, rf_in_c, diff_out_c, pwm_out_c, 
        pwm_out_p_c, led_0_6, led_0_5, led_0_4, led_0_3, led_0_2, 
        led_0_1, led_0_0;
    wire [63:0]\phase_increment[1] ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(64[33:48])
    wire [63:0]\phase_increment[0] ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(64[33:48])
    wire [12:0]lo_sinewave;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(69[33:44])
    wire [12:0]lo_cosinewave;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(70[33:46])
    wire [11:0]mix_sinewave;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(73[33:45])
    wire [11:0]mix_cosinewave;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(74[33:47])
    wire [11:0]cic_sine_out;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(77[33:45])
    wire [11:0]cic_cosine_out;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(79[33:47])
    wire [7:0]cic_gain;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(81[33:41])
    wire [11:0]amdemod_out;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(84[33:44])
    
    wire rx_data_valid;
    wire [7:0]rx_byte;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(88[33:40])
    
    wire rx_data_valid1;
    wire [7:0]rx_byte1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(90[33:41])
    
    wire n17684;
    wire [7:0]cic_gain_7__N_544;
    wire [63:0]phase_increment_1__63__N_16;
    wire [63:0]phase_accumulator_adj_6545;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(23[33:50])
    wire [63:0]phase_increment_1__63__N_17;
    wire [63:0]phase_increment_1__63__N_18;
    wire [63:0]phase_increment_1__63__N_19;
    wire [63:0]phase_increment_1__63__N_20;
    wire [63:0]phase_increment_1__63__N_21;
    
    wire n17683, n17682, n17681, n17680, n17679, n17678, n17677, 
        n17676, n17675, n17674, n17673, n17672, n17671, n17670, 
        n17669, n17668, n17662, n17661, n17660, n17659, n17658, 
        n17657, n17656, n17655, n17654, n17653, n17652, n17651, 
        n17650, n17649, n17648, n17647, n17646, n17645, n17644, 
        n17643, n17642, n17641, n17640, n17639, n17638, n17637, 
        n17636, n17635, n17634, n17633, n17632, n17631, n17629, 
        n17628, n17627, n17626, n17625, n17624, n17623, n17622, 
        n17621, n17620, n17327, n17326, n17325, n17324, n17323, 
        n19627, n17321, n17320, n17319, n17318, n17317, n17316, 
        n17315, n17314, n17313, n17312, n17311, n17310, n17309, 
        n17308, n17307, n17306, n17305, n17304, n17299, n17298, 
        n17297, n17296, n17295, n17294, n17293, n17292, n17291, 
        n17290, n17289, n17288, n17287, n17286, n17285, n17284, 
        n17283, n17282, n17277, n17276, n17275, n17274, n17273, 
        n17272, n17271, n17270, n17269, n17268, n17267, n17266, 
        n17265, n17264, n17263, n17262, n17619, n19606, n19605;
    wire [11:0]sine_table_value;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(17[32:48])
    
    wire n1480;
    wire [11:0]cosine_table_value;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(21[32:50])
    
    wire n90, n87, n84, n81, n78, n75, n72, n69, n66, n63, 
        n60, n57, n54, n19792, n141, n141_adj_3522, n1601, n17618, 
        n17617, n1616, n1626, n1632, n1635, n17910, n19626, n17909, 
        n19625, n17908, n17616, n19603, n1554, n1475, n19436, 
        n1494, n37, n1491;
    wire [71:0]integrator_tmp;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(60[35:49])
    wire [71:0]integrator_d_tmp;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(60[51:67])
    wire [71:0]integrator1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(61[35:46])
    wire [71:0]integrator2;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(61[48:59])
    wire [71:0]integrator3;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(61[61:72])
    wire [71:0]integrator4;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(61[74:85])
    wire [71:0]integrator5;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(61[87:98])
    wire [71:0]comb6;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[35:40])
    wire [71:0]comb_d6;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[42:49])
    wire [71:0]comb7;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[51:56])
    wire [71:0]comb_d7;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[58:65])
    wire [71:0]comb8;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[67:72])
    wire [71:0]comb_d8;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[74:81])
    wire [71:0]comb9;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[83:88])
    wire [71:0]comb_d9;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[90:97])
    
    wire n19624;
    wire [11:0]count;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(65[35:40])
    wire [71:0]integrator1_71__N_960;
    wire [71:0]integrator2_71__N_1032;
    wire [71:0]integrator3_71__N_1104;
    wire [71:0]integrator4_71__N_1176;
    wire [71:0]integrator5_71__N_1248;
    
    wire n17615, n17614, n17613, n17612, n17611, n17610, n17609, 
        n17608, n17607, n17606;
    wire [71:0]comb6_71__N_1993;
    wire [71:0]comb7_71__N_2065;
    wire [71:0]comb8_71__N_2137;
    wire [71:0]comb9_71__N_2209;
    
    wire n19602, n19601, n19435, cout, n183, n180, n177, n174;
    wire [71:0]integrator_tmp_adj_6556;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(60[35:49])
    wire [71:0]integrator_d_tmp_adj_6557;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(60[51:67])
    wire [71:0]integrator1_adj_6558;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(61[35:46])
    wire [71:0]integrator2_adj_6559;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(61[48:59])
    wire [71:0]integrator3_adj_6560;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(61[61:72])
    wire [71:0]integrator4_adj_6561;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(61[74:85])
    wire [71:0]integrator5_adj_6562;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(61[87:98])
    wire [71:0]comb6_adj_6563;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[35:40])
    wire [71:0]comb_d6_adj_6564;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[42:49])
    wire [71:0]comb7_adj_6565;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[51:56])
    wire [71:0]comb_d7_adj_6566;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[58:65])
    wire [71:0]comb8_adj_6567;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[67:72])
    wire [71:0]comb_d8_adj_6568;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[74:81])
    wire [71:0]comb9_adj_6569;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[83:88])
    wire [71:0]comb_d9_adj_6570;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[90:97])
    wire [71:0]comb10_adj_6571;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[99:105])
    
    wire n1428;
    wire [11:0]count_adj_6572;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(65[35:40])
    wire [71:0]integrator1_71__N_960_adj_6573;
    wire [71:0]integrator2_71__N_1032_adj_6574;
    wire [71:0]integrator3_71__N_1104_adj_6575;
    wire [71:0]integrator4_71__N_1176_adj_6576;
    wire [71:0]integrator5_71__N_1248_adj_6577;
    
    wire n17605, n17604, n17603, n17602, n17601, n17600, n17599, 
        n17598, n17597, n17596, n171, n168, n165, n162, n159, 
        n156, n153, n150, n147, n144, n141_adj_4975, n138, n135, 
        n132, n129, n126, n123, n120, n117, n114, n111, n108, 
        n105, n102;
    wire [71:0]comb6_71__N_1993_adj_6589;
    wire [71:0]comb7_71__N_2065_adj_6590;
    wire [71:0]comb8_71__N_2137_adj_6591;
    wire [71:0]comb9_71__N_2209_adj_6592;
    
    wire n17448, n17261, n17260, n17259, n17258, n17257, n17256, 
        n17255, n17254, n17253, n17251, n17250, n17249, n17248, 
        n17247, n99, n96, n93, n90_adj_5264, n87_adj_5265, n84_adj_5266, 
        n81_adj_5267, n78_adj_5268, cout_adj_5269, n61, n58, n55, 
        n52, n49, n46, n43, n40, n37_adj_5270, n34, n31, n28, 
        cout_adj_5271, n1416, n17246, n17245;
    wire [25:0]square_sum;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(18[26:36])
    wire [23:0]i_squared;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(22[34:43])
    wire [23:0]q_squared;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(27[34:43])
    
    wire n17906;
    wire [14:0]amdemod_out_d_11__N_2358;
    
    wire n36, n35, n34_adj_5272, n33, n32, n31_adj_5273, n30, 
        n29, n28_adj_5274, n27, n26, n25, n24;
    wire [14:0]amdemod_out_d_11__N_2365;
    
    wire n17447, n17595, n17594, n17593, n17592, n17591, n17590, 
        n17589, n17588, n17587, n17586, amdemod_out_d_11__N_2363, 
        amdemod_out_d_11__N_2501, amdemod_out_d_11__N_2504, amdemod_out_d_11__N_2507, 
        amdemod_out_d_11__N_2510, amdemod_out_d_11__N_2513, amdemod_out_d_11__N_2516, 
        n17244, n17243;
    wire [14:0]amdemod_out_d_11__N_2370;
    
    wire n17242, n17241;
    wire [14:0]amdemod_out_d_11__N_2369;
    
    wire n23, n22, n21, n20, n19, n18, n17, n16, n15, n14, 
        n13, n12, n11, n16248, n16247, n16246, n16245, n16244, 
        n16239, n16238, n16237, n16236, n16235, n16234, amdemod_out_d_11__N_2564, 
        amdemod_out_d_11__N_2567, amdemod_out_d_11__N_2570, amdemod_out_d_11__N_2573, 
        amdemod_out_d_11__N_2576, amdemod_out_d_11__N_2579, amdemod_out_d_11__N_2582, 
        amdemod_out_d_11__N_2585, amdemod_out_d_11__N_2588, amdemod_out_d_11__N_2591, 
        amdemod_out_d_11__N_2594, amdemod_out_d_11__N_2597, amdemod_out_d_11__N_2600;
    wire [14:0]amdemod_out_d_11__N_2380;
    wire [14:0]amdemod_out_d_11__N_2379;
    
    wire n10, n9, n8, n7, n6, n5, n4, n3, n2, amdemod_out_d_11__N_2642, 
        amdemod_out_d_11__N_2645, amdemod_out_d_11__N_2648, amdemod_out_d_11__N_2651, 
        amdemod_out_d_11__N_2654, amdemod_out_d_11__N_2657, amdemod_out_d_11__N_2660, 
        amdemod_out_d_11__N_2663, amdemod_out_d_11__N_2666, amdemod_out_d_11__N_2669, 
        amdemod_out_d_11__N_2672, amdemod_out_d_11__N_2675, amdemod_out_d_11__N_2678;
    wire [14:0]amdemod_out_d_11__N_2390;
    wire [14:0]amdemod_out_d_11__N_2389;
    
    wire amdemod_out_d_11__N_2720, amdemod_out_d_11__N_2723, amdemod_out_d_11__N_2726, 
        amdemod_out_d_11__N_2729, amdemod_out_d_11__N_2732, amdemod_out_d_11__N_2735, 
        amdemod_out_d_11__N_2738, amdemod_out_d_11__N_2741, amdemod_out_d_11__N_2744, 
        amdemod_out_d_11__N_2747, amdemod_out_d_11__N_2750, amdemod_out_d_11__N_2753, 
        amdemod_out_d_11__N_2756;
    wire [14:0]amdemod_out_d_11__N_2400;
    wire [14:0]amdemod_out_d_11__N_2399;
    
    wire amdemod_out_d_11__N_2798, amdemod_out_d_11__N_2801, amdemod_out_d_11__N_2804, 
        amdemod_out_d_11__N_2807, amdemod_out_d_11__N_2810, amdemod_out_d_11__N_2813, 
        amdemod_out_d_11__N_2816, amdemod_out_d_11__N_2819, amdemod_out_d_11__N_2822, 
        amdemod_out_d_11__N_2825, amdemod_out_d_11__N_2828, amdemod_out_d_11__N_2831, 
        amdemod_out_d_11__N_2834;
    wire [14:0]amdemod_out_d_11__N_2410;
    wire [14:0]amdemod_out_d_11__N_2409;
    wire [9:0]count_adj_6635;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(43[25:30])
    wire [11:0]data_in_reg;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(44[25:36])
    
    wire n17585;
    wire [31:0]data_in_reg_11__N_2898;
    
    wire n17584, n17583, n17582, n17446, n17445, n19434, n1465, 
        n17581, n17579, n17578, n17577, n17576, n17575, n17574, 
        n17573, n17572, n19433, n17571, n17570, n17569, n17568, 
        n17567, n17566, n17565, n17564, n17563, n17562, n19587, 
        n19586, n1447, n17444, n1444, n19863, n19862, n1441, n17560, 
        n17559, n17558, n17557, n17556, n17555, n17554, n17553, 
        n17552, n17240, n17239, n17238, n17551, n17550, n17549, 
        n17548, n17547, n17237, n17236, n17235, n17234, n17229, 
        n17228, n17227, n17226, n17225, n17224, n17223, n17222, 
        n17221, n17220, n17219, n17218, n1438, n17443, n19765, 
        n19764, n1488, n19762, n17442, n17441, n17905, n19585, 
        n19582, n17440, n19581, n17439, n17438, n17437, n19799, 
        n17436, n19440, n19857, n17435, n17434, n17433, n19579, 
        n17432, n1729, n1726, n1723, n1720, n1715, n17431, n17430, 
        n17429, n17427, n17426, n82, n17425, n17424, n17423, n17422, 
        n19432, n17421, n17420, n1823, n1820, n1817, n1814, n1809, 
        n1804, n1794, n174_adj_5285, n1945, n1935, n8_adj_5286, 
        n1917, n1914, n1908, n1898, n1541, n1538, n1535, n1532, 
        n1527, n1522, n2058, n2055, n2052, n2049, n2044, n2039, 
        n135_adj_5287, n2029, n19578, n19295, n198, n17419, n2011, 
        n2008, n19577, n19576, n61_adj_5288, n62, n63_adj_5289, 
        n64, n65, n66_adj_5290, n67, n68, n70, n19575, n17418, 
        n17904, n17903, n17417, n17902, n17546, n1648, n17416, 
        n17901, n171_adj_5291, n1710, n1700, n309, n138_adj_5292, 
        n306, n1776, n1773, n1770, n1767, n1762, n1757, n17415, 
        n1747, n1883, n204, n300, n17414, n19426, n17413, n17412, 
        n17411, n1836, n1512, n1433, n1485, n2002, n17410, n1992, 
        n315, n1977, n1964, n1961, n1958, n1955, n1950, n19856, 
        n2076, n2086, n2091, n2096, n2099, n2102, n2105, n2118, 
        cout_adj_5293, n2133, n2143, n2149, n2152, n189, n2165, 
        n2180, n2190, n2196, n2199, n186, n2212, n2227, n2237, 
        n19553, n2243, n2246, n85, n7_adj_5294, n19431, n2259, 
        n2274, n17409, n2284, n2290, n2293, n183_adj_5295, n2311, 
        n2321, n118, n2326, n2331, n2334, n2337, n2340, cout_adj_5296, 
        n76, n2353, n2368, n2378, n2384, n2387, n258, n2400, 
        n2415, n2425, n19604, n2431, n2434, n201, n249, n2452, 
        n2462, n2467, n2472, n2475, n2478, n2481, n243, n2499, 
        n17545, n2509, n264, n2514, n2519, n2522, n2525, n2528, 
        n156_adj_5297, n2541, n273, n2556, n2566, n2572, n2575, 
        n213, n2588, n195, n2603, n2613, n17217, n2619, n6_adj_5298, 
        n2622, n276, n26_adj_5299, n2635, n5_adj_5300, n2650, n4_adj_5301, 
        n2660, n19682, n2666, n2669, n153_adj_5302, n228, n2682, 
        n2697, n2707, n19679, n2713, n2716, n267, n2729, n2744, 
        n174_adj_5303, n2754, n19828, n2760, n17408, n2763, n3_adj_5304, 
        n210, n17216, n237, n2776, n132_adj_5305, n2823, n2838, 
        n2848, n16233, n2854, n171_adj_5306, n2857, n246, n2870, 
        n17544, n17407, n159_adj_5307, n19827, n240, n2917, n17543, 
        n231, n2932, n2942, n19721, n2948, n2951, n165_adj_5308, 
        n2964, n17215, n162_adj_5309, n2979, n219, n17406, n2989, 
        n19718, n2995, n2998, n97, n207, n3016, n17214, n3026, 
        n3031, n222, n3036, n3039, n3042, n3045, n45, n36_adj_5310, 
        n3058, n3073, n3083, n3089, n3092, n225, n270, n3105, 
        n106, n132_adj_5311, n3120, n3130, n19419, n3136, n3139, 
        n3152, n303, n17213, n3167, n129_adj_5312, n3177, n3183, 
        n3186, n192, n3199, n297, n3214, n3224, n3230, n108_adj_5313, 
        n3233, cout_adj_5314, n3246, n120_adj_5315, n19478, n255, 
        n3293, n3308, n117_adj_5316, n3318, n3324, n3327, n3345, 
        n312, n91, n3355, n3360, n3365, n3368, n3371, n3374, 
        n162_adj_5317, n3392, cout_adj_5318, n3402, n103, n3407, 
        n3412, n3415, n3418, n105_adj_5319, n3421, n147_adj_5320, 
        n17212, n159_adj_5321, n94, n19662, n234, n3486, n3496, 
        n3501, n3506, n3509, n3512, n3515, n19430, n3528, n84_adj_5322, 
        n19700, n3580, n3590, n216, n3595, n81_adj_5323, n3600, 
        n79, n3603, n3606, n3609, n183_adj_5324, n88, n3622, n321, 
        n3637, n3647, n3653, n3656, n180_adj_5325, n177_adj_5326, 
        n3674, n17405, n3684, n3689, n3694, n3697, n3700, n3703, 
        n17900, n279, n3716, n18645, n17404, n17403, n282, n17402, 
        n3768, n17401, n3778, n252, cout_adj_5327, n3783, n3788, 
        n3791, n3794, n3797, n19302, n17400, n3815, n17399, n3825, 
        n3830, n3835, n3838, n3841, n3844, cout_adj_5328, n17398, 
        n3862, n3872, n3877, n3882, n3885, n3888, n3891, n294, 
        n3904, n17397, n3919, n3929, n3935, n3938, n112, n115, 
        n3951, n17396, n3966, n3976, n19763, n3982, n3985, n109, 
        n3998, n19760, n19447, n150_adj_5329, n19301, n17539, n4050, 
        n4060, n4065, n4070, n4073, n4076, n4079, n78_adj_5330, 
        n19300, n4097, n17395, n4107, n4112, n4117, n4120, n4123, 
        n4126, n318, n90_adj_5331, n4139, n4154, n17207, n4164, 
        n19429, n4170, n144_adj_5332, n4173, n114_adj_5333, n96_adj_5334, 
        n102_adj_5335, n87_adj_5336, n4186, n93_adj_5337, n4201, n4211, 
        n4217, n4220, n126_adj_5338, n100, n111_adj_5339, n285, 
        n99_adj_5340, n180_adj_5341, n288, n19761, n4248, n17538, 
        n4258, n4264, n4267, n123_adj_5342, n17206, n135_adj_5343, 
        n291, n147_adj_5344, n4295, n19299, n4305, n4308, n4311, 
        n4314, n138_adj_5345, n150_adj_5346, n165_adj_5347, n17537, 
        n4342, n19555, n4355, n4358, n4361, n144_adj_5348, n153_adj_5349, 
        n19554, n168_adj_5350, n177_adj_5351, n19552, n156_adj_5352, 
        n261, n168_adj_5353, n2_adj_5354, n19551, n19825, n19824, 
        n9_adj_5355, n10_adj_5356, n11_adj_5357, n12_adj_5358, n13_adj_5359, 
        n14_adj_5360, n15_adj_5361, n16_adj_5362, n17_adj_5363, n18_adj_5364, 
        n19_adj_5365, n20_adj_5366, n21_adj_5367, n22_adj_5368, n23_adj_5369, 
        n24_adj_5370, n25_adj_5371, n26_adj_5372, n27_adj_5373, n28_adj_5374, 
        n29_adj_5375, n30_adj_5376, n31_adj_5377, n32_adj_5378, n33_adj_5379, 
        n34_adj_5380, n35_adj_5381, n36_adj_5382, n37_adj_5383, n19823, 
        n19822, n2_adj_5384, n3_adj_5385, n4_adj_5386, n5_adj_5387, 
        n6_adj_5388, n7_adj_5389, n8_adj_5390, n9_adj_5391, n10_adj_5392, 
        n11_adj_5393, n12_adj_5394, n13_adj_5395, n14_adj_5396, n15_adj_5397, 
        n16_adj_5398, n17_adj_5399, n18_adj_5400, n19_adj_5401, n20_adj_5402, 
        n21_adj_5403, n22_adj_5404, n23_adj_5405, n24_adj_5406, n25_adj_5407, 
        n26_adj_5408, n27_adj_5409, n28_adj_5410, n29_adj_5411, n30_adj_5412, 
        n31_adj_5413, n32_adj_5414, n33_adj_5415, n34_adj_5416, n35_adj_5417, 
        n36_adj_5418, n37_adj_5419, n2_adj_5420, n3_adj_5421, n4_adj_5422, 
        n5_adj_5423, n6_adj_5424, n7_adj_5425, n8_adj_5426, n9_adj_5427, 
        n10_adj_5428, n11_adj_5429, n12_adj_5430, n13_adj_5431, n14_adj_5432, 
        n15_adj_5433, n16_adj_5434, n17_adj_5435, n18_adj_5436, n19_adj_5437, 
        n20_adj_5438, n21_adj_5439, n22_adj_5440, n23_adj_5441, n24_adj_5442, 
        n25_adj_5443, n26_adj_5444, n27_adj_5445, n28_adj_5446, n29_adj_5447, 
        n30_adj_5448, n31_adj_5449, n32_adj_5450, n33_adj_5451, n34_adj_5452, 
        n35_adj_5453, n36_adj_5454, n37_adj_5455, n19550, n19543, 
        n19542, n2_adj_5456, n3_adj_5457, n4_adj_5458, n5_adj_5459, 
        n6_adj_5460, n7_adj_5461, n8_adj_5462, n9_adj_5463, n10_adj_5464, 
        n11_adj_5465, n12_adj_5466, n13_adj_5467, n14_adj_5468, n15_adj_5469, 
        n16_adj_5470, n17_adj_5471, n18_adj_5472, n19_adj_5473, n20_adj_5474, 
        n21_adj_5475, n22_adj_5476, n23_adj_5477, n24_adj_5478, n25_adj_5479, 
        n26_adj_5480, n27_adj_5481, n28_adj_5482, n29_adj_5483, n30_adj_5484, 
        n31_adj_5485, n32_adj_5486, n33_adj_5487, n34_adj_5488, n35_adj_5489, 
        n36_adj_5490, n37_adj_5491, n19541, n2_adj_5492, n3_adj_5493, 
        n4_adj_5494, n5_adj_5495, n6_adj_5496, n7_adj_5497, n8_adj_5498, 
        n9_adj_5499, n10_adj_5500, n11_adj_5501, n12_adj_5502, n13_adj_5503, 
        n14_adj_5504, n15_adj_5505, n16_adj_5506, n17_adj_5507, n18_adj_5508, 
        n19_adj_5509, n20_adj_5510, n21_adj_5511, n22_adj_5512, n23_adj_5513, 
        n24_adj_5514, n25_adj_5515, n26_adj_5516, n27_adj_5517, n28_adj_5518, 
        n29_adj_5519, n30_adj_5520, n31_adj_5521, n32_adj_5522, n33_adj_5523, 
        n34_adj_5524, n35_adj_5525, n36_adj_5526, n37_adj_5527, n2_adj_5528, 
        n3_adj_5529, n4_adj_5530, n5_adj_5531, n6_adj_5532, n7_adj_5533, 
        n8_adj_5534, n9_adj_5535, n10_adj_5536, n11_adj_5537, n12_adj_5538, 
        n13_adj_5539, n14_adj_5540, n15_adj_5541, n16_adj_5542, n17_adj_5543, 
        n18_adj_5544, n19_adj_5545, n20_adj_5546, n21_adj_5547, n22_adj_5548, 
        n23_adj_5549, n24_adj_5550, n25_adj_5551, n26_adj_5552, n27_adj_5553, 
        n28_adj_5554, n29_adj_5555, n30_adj_5556, n31_adj_5557, n32_adj_5558, 
        n33_adj_5559, n34_adj_5560, n35_adj_5561, n36_adj_5562, n37_adj_5563, 
        n2_adj_5564, n3_adj_5565, n4_adj_5566, n5_adj_5567, n6_adj_5568, 
        n7_adj_5569, n8_adj_5570, n9_adj_5571, n10_adj_5572, n11_adj_5573, 
        n12_adj_5574, n13_adj_5575, n14_adj_5576, n15_adj_5577, n16_adj_5578, 
        n17_adj_5579, n18_adj_5580, n19_adj_5581, n20_adj_5582, n21_adj_5583, 
        n22_adj_5584, n23_adj_5585, n24_adj_5586, n25_adj_5587, n26_adj_5588, 
        n27_adj_5589, n28_adj_5590, n29_adj_5591, n30_adj_5592, n31_adj_5593, 
        n32_adj_5594, n33_adj_5595, n34_adj_5596, n35_adj_5597, n36_adj_5598, 
        n37_adj_5599, n19737, n19736, n19735, n19807, n17394, n17393, 
        n17392, n17391, n17390, n17389, n17388, n17387, n17386, 
        n17385, n17205, n126_adj_5600, n123_adj_5601, n17204, n120_adj_5602, 
        n117_adj_5603, n17203, n17383, n17382, n17381, n17380, n17379, 
        n17378, n114_adj_5604, n17377, n17376, n17375, n16232, n111_adj_5605, 
        n108_adj_5606, n105_adj_5607, n102_adj_5608, n99_adj_5609, n96_adj_5610, 
        n93_adj_5611, n19734, n19733, n19526, n78_adj_5612, n81_adj_5613, 
        n84_adj_5614, n87_adj_5615, n90_adj_5616, n93_adj_5617, n96_adj_5618, 
        n99_adj_5619, n102_adj_5620, n105_adj_5621, n108_adj_5622, n111_adj_5623, 
        n114_adj_5624, n117_adj_5625, n120_adj_5626, n19525, cout_adj_5627, 
        n78_adj_5628, n81_adj_5629, n84_adj_5630, n87_adj_5631, n90_adj_5632, 
        n93_adj_5633, n96_adj_5634, n99_adj_5635, n102_adj_5636, n105_adj_5637, 
        n108_adj_5638, n111_adj_5639, n114_adj_5640, n117_adj_5641, 
        n120_adj_5642, n123_adj_5643, n126_adj_5644, n129_adj_5645, 
        n132_adj_5646, n135_adj_5647, n138_adj_5648, n141_adj_5649, 
        n144_adj_5650, n147_adj_5651, n150_adj_5652, n153_adj_5653, 
        n156_adj_5654, n159_adj_5655, n162_adj_5656, n165_adj_5657, 
        n168_adj_5658, n171_adj_5659, n174_adj_5660, n177_adj_5661, 
        n180_adj_5662, n183_adj_5663, n36_adj_5664, n42, n45_adj_5665, 
        n48, n51, n54_adj_5666, n57_adj_5667, n60_adj_5668, n63_adj_5669, 
        n66_adj_5670, n69_adj_5671, n72_adj_5672, n75_adj_5673, n78_adj_5674, 
        n78_adj_5675, n81_adj_5676, n84_adj_5677, n87_adj_5678, n90_adj_5679, 
        n93_adj_5680, n96_adj_5681, n99_adj_5682, n102_adj_5683, n105_adj_5684, 
        n108_adj_5685, n111_adj_5686, n114_adj_5687, n117_adj_5688, 
        n120_adj_5689, n123_adj_5690, n126_adj_5691, n129_adj_5692, 
        n132_adj_5693, n135_adj_5694, n138_adj_5695, n141_adj_5696, 
        n144_adj_5697, n147_adj_5698, n150_adj_5699, n153_adj_5700, 
        n156_adj_5701, n159_adj_5702, n162_adj_5703, n165_adj_5704, 
        n168_adj_5705, n171_adj_5706, n174_adj_5707, n177_adj_5708, 
        n180_adj_5709, n183_adj_5710, n36_adj_5711, n42_adj_5712, n45_adj_5713, 
        n48_adj_5714, n51_adj_5715, n54_adj_5716, n57_adj_5717, n60_adj_5718, 
        n63_adj_5719, n66_adj_5720, n69_adj_5721, n72_adj_5722, n75_adj_5723, 
        n78_adj_5724, n78_adj_5725, n81_adj_5726, n84_adj_5727, n87_adj_5728, 
        n90_adj_5729, n93_adj_5730, n96_adj_5731, n99_adj_5732, n102_adj_5733, 
        n105_adj_5734, n108_adj_5735, n111_adj_5736, n114_adj_5737, 
        n117_adj_5738, n120_adj_5739, n123_adj_5740, n126_adj_5741, 
        n129_adj_5742, n132_adj_5743, n135_adj_5744, n138_adj_5745, 
        n141_adj_5746, n144_adj_5747, n147_adj_5748, n150_adj_5749, 
        n153_adj_5750, n156_adj_5751, n159_adj_5752, n162_adj_5753, 
        n165_adj_5754, n168_adj_5755, n171_adj_5756, n174_adj_5757, 
        n177_adj_5758, n180_adj_5759, n183_adj_5760, n78_adj_5761, n81_adj_5762, 
        n84_adj_5763, n87_adj_5764, n90_adj_5765, n93_adj_5766, n96_adj_5767, 
        n99_adj_5768, n102_adj_5769, n105_adj_5770, n108_adj_5771, n111_adj_5772, 
        n114_adj_5773, n117_adj_5774, n120_adj_5775, n123_adj_5776, 
        n126_adj_5777, n129_adj_5778, n132_adj_5779, n135_adj_5780, 
        n138_adj_5781, n141_adj_5782, n144_adj_5783, n147_adj_5784, 
        n150_adj_5785, n153_adj_5786, n156_adj_5787, n159_adj_5788, 
        n162_adj_5789, n165_adj_5790, n168_adj_5791, n171_adj_5792, 
        n174_adj_5793, n177_adj_5794, n180_adj_5795, n183_adj_5796, 
        n36_adj_5797, n42_adj_5798, n45_adj_5799, n48_adj_5800, n51_adj_5801, 
        n54_adj_5802, n57_adj_5803, n60_adj_5804, n63_adj_5805, n66_adj_5806, 
        n69_adj_5807, n72_adj_5808, n75_adj_5809, n78_adj_5810, n36_adj_5811, 
        n42_adj_5812, n45_adj_5813, n48_adj_5814, n51_adj_5815, n54_adj_5816, 
        n57_adj_5817, n60_adj_5818, n63_adj_5819, n66_adj_5820, n69_adj_5821, 
        n72_adj_5822, n75_adj_5823, n78_adj_5824, n78_adj_5825, n81_adj_5826, 
        n84_adj_5827, n87_adj_5828, n90_adj_5829, n93_adj_5830, n96_adj_5831, 
        n99_adj_5832, n102_adj_5833, n105_adj_5834, n108_adj_5835, n111_adj_5836, 
        n114_adj_5837, n117_adj_5838, n120_adj_5839, n19524, cout_adj_5840, 
        n36_adj_5841, n42_adj_5842, n45_adj_5843, n48_adj_5844, n51_adj_5845, 
        n54_adj_5846, n57_adj_5847, n60_adj_5848, n63_adj_5849, n66_adj_5850, 
        n69_adj_5851, n72_adj_5852, n75_adj_5853, n78_adj_5854, n78_adj_5855, 
        n81_adj_5856, n84_adj_5857, n87_adj_5858, n90_adj_5859, n93_adj_5860, 
        n96_adj_5861, n99_adj_5862, n102_adj_5863, n105_adj_5864, n108_adj_5865, 
        n111_adj_5866, n114_adj_5867, n117_adj_5868, n120_adj_5869, 
        n123_adj_5870, n126_adj_5871, n129_adj_5872, n132_adj_5873, 
        n135_adj_5874, n138_adj_5875, n141_adj_5876, n144_adj_5877, 
        n147_adj_5878, n150_adj_5879, n153_adj_5880, n156_adj_5881, 
        n159_adj_5882, n162_adj_5883, n165_adj_5884, n168_adj_5885, 
        n171_adj_5886, n174_adj_5887, n177_adj_5888, n180_adj_5889, 
        n183_adj_5890, cout_adj_5891, n78_adj_5892, n81_adj_5893, n84_adj_5894, 
        n87_adj_5895, n90_adj_5896, n93_adj_5897, n96_adj_5898, n99_adj_5899, 
        n102_adj_5900, n105_adj_5901, n108_adj_5902, n111_adj_5903, 
        n114_adj_5904, n117_adj_5905, n120_adj_5906, n123_adj_5907, 
        n126_adj_5908, n129_adj_5909, n132_adj_5910, n135_adj_5911, 
        n138_adj_5912, n141_adj_5913, n144_adj_5914, n147_adj_5915, 
        n150_adj_5916, n153_adj_5917, n156_adj_5918, n159_adj_5919, 
        n162_adj_5920, n165_adj_5921, n168_adj_5922, n171_adj_5923, 
        n174_adj_5924, n177_adj_5925, n180_adj_5926, n183_adj_5927, 
        n78_adj_5928, n81_adj_5929, n84_adj_5930, n87_adj_5931, n90_adj_5932, 
        n93_adj_5933, n96_adj_5934, n99_adj_5935, n102_adj_5936, n105_adj_5937, 
        n108_adj_5938, n111_adj_5939, n114_adj_5940, n117_adj_5941, 
        n120_adj_5942, n123_adj_5943, n126_adj_5944, n129_adj_5945, 
        n132_adj_5946, n135_adj_5947, n138_adj_5948, n141_adj_5949, 
        n144_adj_5950, n147_adj_5951, n150_adj_5952, n153_adj_5953, 
        n156_adj_5954, n159_adj_5955, n162_adj_5956, n165_adj_5957, 
        n168_adj_5958, n171_adj_5959, n174_adj_5960, n177_adj_5961, 
        n180_adj_5962, n183_adj_5963, n78_adj_5964, n81_adj_5965, n84_adj_5966, 
        n87_adj_5967, n90_adj_5968, n93_adj_5969, n96_adj_5970, n99_adj_5971, 
        n102_adj_5972, n105_adj_5973, n108_adj_5974, n111_adj_5975, 
        n114_adj_5976, n117_adj_5977, n120_adj_5978, n123_adj_5979, 
        n126_adj_5980, n129_adj_5981, n132_adj_5982, n135_adj_5983, 
        n138_adj_5984, n141_adj_5985, n144_adj_5986, n147_adj_5987, 
        n150_adj_5988, n153_adj_5989, n156_adj_5990, n159_adj_5991, 
        n162_adj_5992, n165_adj_5993, n168_adj_5994, n171_adj_5995, 
        n174_adj_5996, n177_adj_5997, n180_adj_5998, n183_adj_5999, 
        n78_adj_6000, n81_adj_6001, n84_adj_6002, n87_adj_6003, n90_adj_6004, 
        n93_adj_6005, n96_adj_6006, n99_adj_6007, n102_adj_6008, n105_adj_6009, 
        n108_adj_6010, n111_adj_6011, n114_adj_6012, n117_adj_6013, 
        n120_adj_6014, n123_adj_6015, n126_adj_6016, n129_adj_6017, 
        n132_adj_6018, n135_adj_6019, n138_adj_6020, n141_adj_6021, 
        n144_adj_6022, n147_adj_6023, n150_adj_6024, n153_adj_6025, 
        n156_adj_6026, n159_adj_6027, n162_adj_6028, n165_adj_6029, 
        n168_adj_6030, n171_adj_6031, n174_adj_6032, n177_adj_6033, 
        n180_adj_6034, n183_adj_6035, n34_adj_6036, n40_adj_6037, n43_adj_6038, 
        n46_adj_6039, n49_adj_6040, n52_adj_6041, n55_adj_6042, n58_adj_6043, 
        n61_adj_6044, n64_adj_6045, n67_adj_6046, n70_adj_6047, n73, 
        n76_adj_6048, n34_adj_6049, n40_adj_6050, n43_adj_6051, n46_adj_6052, 
        n49_adj_6053, n52_adj_6054, n55_adj_6055, n58_adj_6056, n61_adj_6057, 
        n64_adj_6058, n67_adj_6059, n70_adj_6060, n73_adj_6061, n76_adj_6062, 
        n34_adj_6063, n40_adj_6064, n43_adj_6065, n46_adj_6066, n49_adj_6067, 
        n52_adj_6068, n55_adj_6069, n58_adj_6070, n61_adj_6071, n64_adj_6072, 
        n67_adj_6073, n70_adj_6074, n73_adj_6075, n76_adj_6076, n34_adj_6077, 
        n40_adj_6078, n43_adj_6079, n46_adj_6080, n49_adj_6081, n52_adj_6082, 
        n55_adj_6083, n58_adj_6084, n61_adj_6085, n64_adj_6086, n67_adj_6087, 
        n70_adj_6088, n73_adj_6089, n76_adj_6090, cout_adj_6091, cout_adj_6092, 
        n78_adj_6093, n81_adj_6094, n84_adj_6095, n87_adj_6096, n90_adj_6097, 
        n93_adj_6098, n96_adj_6099, n99_adj_6100, n102_adj_6101, n105_adj_6102, 
        n108_adj_6103, n111_adj_6104, n114_adj_6105, n117_adj_6106, 
        n120_adj_6107, n123_adj_6108, n126_adj_6109, n129_adj_6110, 
        n132_adj_6111, n135_adj_6112, n138_adj_6113, n141_adj_6114, 
        n144_adj_6115, n147_adj_6116, n150_adj_6117, n153_adj_6118, 
        n156_adj_6119, n159_adj_6120, n162_adj_6121, n165_adj_6122, 
        n168_adj_6123, n171_adj_6124, n174_adj_6125, n177_adj_6126, 
        n180_adj_6127, n183_adj_6128, cout_adj_6129, n19809, n19732, 
        n19731, n36_adj_6130, n28_adj_6131, n31_adj_6132, n34_adj_6133, 
        n37_adj_6134, n40_adj_6135, n43_adj_6136, n46_adj_6137, n49_adj_6138, 
        n52_adj_6139, n55_adj_6140, n58_adj_6141, n61_adj_6142, n34_adj_6143, 
        n40_adj_6144, n43_adj_6145, n46_adj_6146, n49_adj_6147, n52_adj_6148, 
        n55_adj_6149, n58_adj_6150, n61_adj_6151, n64_adj_6152, n67_adj_6153, 
        n70_adj_6154, n73_adj_6155, n76_adj_6156, n19425, n19723, 
        n34_adj_6157, n40_adj_6158, n43_adj_6159, n46_adj_6160, n49_adj_6161, 
        n52_adj_6162, n55_adj_6163, n58_adj_6164, n61_adj_6165, n64_adj_6166, 
        n67_adj_6167, n70_adj_6168, n73_adj_6169, n76_adj_6170, n34_adj_6171, 
        n40_adj_6172, n43_adj_6173, n46_adj_6174, n49_adj_6175, n52_adj_6176, 
        n55_adj_6177, n58_adj_6178, n61_adj_6179, n64_adj_6180, n67_adj_6181, 
        n70_adj_6182, n73_adj_6183, n76_adj_6184, n19722, n19424, 
        n19423, n19422, n19720, n19719, n17899, n19520, n17202, 
        n17501, n34_adj_6185, n40_adj_6186, n43_adj_6187, n46_adj_6188, 
        n49_adj_6189, n52_adj_6190, n55_adj_6191, n58_adj_6192, n61_adj_6193, 
        n64_adj_6194, n67_adj_6195, n70_adj_6196, n73_adj_6197, n76_adj_6198, 
        n17201, n46_adj_6199, n19519, n19717, n19518, n19629, n19716, 
        n19715, n19517, n19516, n19515, n19514, n19421, n34_adj_6200, 
        n78_adj_6201, n81_adj_6202, n84_adj_6203, n87_adj_6204, n90_adj_6205, 
        n93_adj_6206, n96_adj_6207, n99_adj_6208, n102_adj_6209, n105_adj_6210, 
        n108_adj_6211, n111_adj_6212, n114_adj_6213, n117_adj_6214, 
        n120_adj_6215, n123_adj_6216, n126_adj_6217, n129_adj_6218, 
        n132_adj_6219, n135_adj_6220, n138_adj_6221, n141_adj_6222, 
        n144_adj_6223, n147_adj_6224, n150_adj_6225, n153_adj_6226, 
        n156_adj_6227, n159_adj_6228, n162_adj_6229, n165_adj_6230, 
        n168_adj_6231, n171_adj_6232, n174_adj_6233, n177_adj_6234, 
        n180_adj_6235, n183_adj_6236, n24_adj_6237, n27_adj_6238, n30_adj_6239, 
        n33_adj_6240, n36_adj_6241, n39, n42_adj_6242, n45_adj_6243, 
        n48_adj_6244, n78_adj_6245, n81_adj_6246, n84_adj_6247, n87_adj_6248, 
        n90_adj_6249, n93_adj_6250, n96_adj_6251, n99_adj_6252, n102_adj_6253, 
        n105_adj_6254, n108_adj_6255, n111_adj_6256, n114_adj_6257, 
        n117_adj_6258, n120_adj_6259, n123_adj_6260, n126_adj_6261, 
        n129_adj_6262, n132_adj_6263, n135_adj_6264, n138_adj_6265, 
        n141_adj_6266, n144_adj_6267, n147_adj_6268, n150_adj_6269, 
        n153_adj_6270, n156_adj_6271, n159_adj_6272, n162_adj_6273, 
        n165_adj_6274, n168_adj_6275, n171_adj_6276, n174_adj_6277, 
        n177_adj_6278, n180_adj_6279, n183_adj_6280, n17200, n17199, 
        n17198, n17197, n17196, n17195, n17194, n17193, n17192, 
        n17191, n17190, n19420, n17185, n17184, n17183, n17182, 
        n17181, n17180, n17179, n17177, n17176, n17175, n17174, 
        n17173, n17172, n17171, n17169, n17168, n17167, n17166, 
        n17165, n17164, cout_adj_6281, n17898, n30_adj_6282, n33_adj_6283, 
        n36_adj_6284, n39_adj_6285, n42_adj_6286, n45_adj_6287, n48_adj_6288, 
        cout_adj_6289, n78_adj_6290, n81_adj_6291, n84_adj_6292, n87_adj_6293, 
        n90_adj_6294, n93_adj_6295, n96_adj_6296, n99_adj_6297, n102_adj_6298, 
        n105_adj_6299, n108_adj_6300, n111_adj_6301, n114_adj_6302, 
        n117_adj_6303, n120_adj_6304, n123_adj_6305, n126_adj_6306, 
        n129_adj_6307, n132_adj_6308, n135_adj_6309, n138_adj_6310, 
        n141_adj_6311, n144_adj_6312, n147_adj_6313, n150_adj_6314, 
        n153_adj_6315, n156_adj_6316, n159_adj_6317, n162_adj_6318, 
        n165_adj_6319, n168_adj_6320, n171_adj_6321, n174_adj_6322, 
        n177_adj_6323, n180_adj_6324, n183_adj_6325, n28_adj_6326, n31_adj_6327, 
        n34_adj_6328, n37_adj_6329, n40_adj_6330, n43_adj_6331, n46_adj_6332, 
        n49_adj_6333, n52_adj_6334, n55_adj_6335, n58_adj_6336, n61_adj_6337, 
        n28_adj_6338, n31_adj_6339, n34_adj_6340, n37_adj_6341, n40_adj_6342, 
        n43_adj_6343, n46_adj_6344, n49_adj_6345, n52_adj_6346, n55_adj_6347, 
        n58_adj_6348, n61_adj_6349, n28_adj_6350, n31_adj_6351, n34_adj_6352, 
        n37_adj_6353, n40_adj_6354, n43_adj_6355, n46_adj_6356, n49_adj_6357, 
        n52_adj_6358, n55_adj_6359, n58_adj_6360, n61_adj_6361, n28_adj_6362, 
        n31_adj_6363, n34_adj_6364, n37_adj_6365, n40_adj_6366, n43_adj_6367, 
        n46_adj_6368, n49_adj_6369, n52_adj_6370, n55_adj_6371, n58_adj_6372, 
        n61_adj_6373, n36_adj_6374, n42_adj_6375, n45_adj_6376, n48_adj_6377, 
        n51_adj_6378, n54_adj_6379, n57_adj_6380, n60_adj_6381, n63_adj_6382, 
        n66_adj_6383, n69_adj_6384, n72_adj_6385, n75_adj_6386, n78_adj_6387, 
        n78_adj_6388, n81_adj_6389, n84_adj_6390, n87_adj_6391, n90_adj_6392, 
        n93_adj_6393, n96_adj_6394, n99_adj_6395, n102_adj_6396, n105_adj_6397, 
        n108_adj_6398, n111_adj_6399, n114_adj_6400, n117_adj_6401, 
        n120_adj_6402, n123_adj_6403, n126_adj_6404, n129_adj_6405, 
        n132_adj_6406, n135_adj_6407, n138_adj_6408, n141_adj_6409, 
        n144_adj_6410, n147_adj_6411, n150_adj_6412, n153_adj_6413, 
        n156_adj_6414, n159_adj_6415, n162_adj_6416, n19702, n165_adj_6417, 
        n168_adj_6418, n171_adj_6419, n19701, n174_adj_6420, n177_adj_6421, 
        n180_adj_6422, n183_adj_6423, n19819, n19688, n19509, n78_adj_6424, 
        n81_adj_6425, n84_adj_6426, n87_adj_6427, n90_adj_6428, n93_adj_6429, 
        n96_adj_6430, n99_adj_6431, n102_adj_6432, n105_adj_6433, n108_adj_6434, 
        n111_adj_6435, n114_adj_6436, n117_adj_6437, n120_adj_6438, 
        n123_adj_6439, n126_adj_6440, n129_adj_6441, n132_adj_6442, 
        n135_adj_6443, n138_adj_6444, n19508, n141_adj_6445, n19580, 
        n144_adj_6446, n147_adj_6447, n150_adj_6448, n153_adj_6449, 
        n156_adj_6450, n159_adj_6451, n162_adj_6452, n19418, n165_adj_6453, 
        n168_adj_6454, n171_adj_6455, n174_adj_6456, n177_adj_6457, 
        n19507, n180_adj_6458, n183_adj_6459, n19574, n19416, n19687, 
        n19686, n36_adj_6460, n19417, n42_adj_6461, n18834, n45_adj_6462, 
        n48_adj_6463, n51_adj_6464, n54_adj_6465, n57_adj_6466, n60_adj_6467, 
        n63_adj_6468, n17918, n66_adj_6469, n17917, n69_adj_6470, 
        n17916, n72_adj_6471, n17915, n75_adj_6472, n17914, n78_adj_6473, 
        n17913, n17912, n17897, n17896, n17449, n17895, n17500, 
        n17894, n17499, n17498, n17497, n17374, n17890, n17496, 
        n17889, n17495, n17482, n17888, n17887, n17494, n17481, 
        n17886, clk_80mhz_enable_238, n17885, n17884, n17480, n17479, 
        n17882, n17373, n17881, n17478, n17880, n17477, n17879, 
        n17372, n17878, n17476, n17877, n17493, n17475, n17876, 
        n17371, n17875, n17474, n17464, n17874, n17463, n78_adj_6474, 
        n17453, n81_adj_6475, n17873, n84_adj_6476, n17492, n87_adj_6477, 
        n17473, n90_adj_6478, n17872, n93_adj_6479, n17491, n96_adj_6480, 
        n99_adj_6481, n17871, n102_adj_6482, n105_adj_6483, n108_adj_6484, 
        n17870, n111_adj_6485, n17462, n114_adj_6486, n17452, n117_adj_6487, 
        n17869, n120_adj_6488, n123_adj_6489, n126_adj_6490, n17868, 
        n129_adj_6491, n17490, n132_adj_6492, n17471, n135_adj_6493, 
        n17867, n138_adj_6494, n141_adj_6495, n17163, n144_adj_6496, 
        n17866, n147_adj_6497, n17489, n150_adj_6498, n17865, n153_adj_6499, 
        n17488, n156_adj_6500, n159_adj_6501, n17370, n162_adj_6502, 
        n165_adj_6503, n168_adj_6504, n171_adj_6505, n174_adj_6506, 
        n177_adj_6507, n17860, n180_adj_6508, n183_adj_6509, n17859, 
        n17858, n17857, n17856, n17855, n17854, n17853, n17852, 
        n17851, n17369, n17850, n17368, n17849, n17848, n17367, 
        n17847, n17366, n17846, n17845, n17844, n17487, n17470, 
        n17843, n17842, n17841, n17840, n17839, n17361, n17838, 
        n17837, n17836, n17360, n17835, n17359, n17834, n4_adj_6510, 
        n17833, n17832, n17358, n17831, n17357, n17830, n17486, 
        n17469, n17828, n17356, n17827, n17355, n17826, n17825, 
        n17824, n17354, n17161, n17823, n17160, n17353, n17159, 
        n13890, n17158, n17157, n17156, n17155, n17154, n17153, 
        n13878, n17152, n13876, n17151, n17822, n17150, n19685, 
        n17149, n19684, n17148, n17484, n17147, n17468, n17146, 
        n17820, n17145, n17352, n17144, n17819, n17143, n17351, 
        n17142, n17818, n17141, n17140, n17817, n17139, n17138, 
        n17816, n17137, n17136, n17815, n17135, n17350, n17134, 
        n17814, n17133, n17349, n17132, n17813, n17131, n17130, 
        n17812, n17129, n17348, n17811, n17347, n17810, cout_adj_6511, 
        n17809, n17461, n17808, n17346, n17807, n17460, n17806, 
        n17345, n17805, n17804, n17459, n17803, n17344, n17467, 
        n17458, n17798, n17451, n17797, n13821, n17796, n17340, 
        n13815, n17795, n17794, n17339, n17793, n17450, n17792, 
        n17338, n17790, n17789, n17788, n17787, n17786, n17785, 
        n17466, n17784, n17337, n17336, n17782, n17335, n17781, 
        n17334, n17780, n17333, n17779, n17332, n17331, n17777, 
        n17330, n17776, n17457, n17775, n17774, n17773, n17772, 
        n17329, n19412, n19683, n19411, n17128, n17127, n17126, 
        n17125, n17124, n17123, n17122, n17121, n17120, n17119, 
        n17117, n17116, n17115, n17114, n17113, n19681, n19410, 
        n17771, n17536, n17535, n17534, n17770, n17769, n17328, 
        n17768, n17533, n17767, n17532, n17531, n17766, n17765, 
        n17764, n17530, n17763, n17529, n17528, n17527, n17762, 
        n17526, n17525, n17761, n17760, n19680, n17456, n19678, 
        n17524, n17756, n17112, n19493, n17755, clk_80mhz_enable_235, 
        n17523, n17754, n17753, n17522, n17521, n17752, n17751, 
        n19677, n16231, n17750, n16230, n17520, n16229, n16228, 
        n19492, n17749, n17519, n17518, n17748, n17747, n17746, 
        n17517, n19294, n16227, n17745, n17744, n19676, n19491, 
        n17743, n17516, n17742, n17515, n17741, n17111, n17740, 
        n17739, n17737, n17736, n17514, n17513, n17735, n17512, 
        n17734, n17511, n17733, n17732, n17731, n17455, n17730, 
        n17729, n17728, n17110, n17727, n17510, n17726, n17725, 
        n17509, n17724, n17723, n17722, n17721, n17720, n17719, 
        n17454, n17508, n17507, n17718, n17717, cout_adj_6512, n17716, 
        n17715, n17506, n17714, n17109, n17108, n17713, n17483, 
        n17505, n17504, n17712, n17711, n17710, n17709, n17708, 
        n17707, n17706, n16226, n17705, n17704, n16225, n17703, 
        n16224, n17702, n16223, n16222, n17701, n17700, n17699, 
        n17698, n17697, n17696, n17695, n17694, n17693, n17692, 
        n17691, n17690, n17503, n17502, n17689, n17688, n17465, 
        n17687, n17686, n17685, n17107, n17106, n17105, n17104, 
        n17103, n17102, n17101, n19668, n17100, n17095, n17094, 
        n17093, n17092, n17091, n17090, n19667, n17089, n17088, 
        n17087, n17086, n17085, n17084, n17083, n19666, n17082, 
        n17081, n17080, n17079, n17078, n17077, n17076, n17075, 
        n17074, n17073, n17072, n17071, n17070, n17069, n17068, 
        n17067, n17066, n17065, n17056, n17055, n17054, n17053, 
        n17052, n17051, n17050, n17049, n17048, n17047, n17046, 
        n17045, n17044, n17043, n17042, n17041, n17040, n17039, 
        n17038, n17037, n17036, n17035, n17034, n17033, n17032, 
        n17031, n17030, n17029, n17028, n17027, n17026, n17025, 
        n17024, n17023, n17022, n17021, n17020, n17019, n17018, 
        n17017, n17016, n17015, n17014, n17013, n17012, n17011, 
        n17010, n17009, n17008, n17007, n17006, n17005, n17004, 
        n17003, n17002, n17001, n17000, n16999, n16998, n16997, 
        n16996, n16995, n16994, n16993, n16992, n16991, n19665, 
        n16990, n16989, n16988, n16987, n16986, n16985, n16984, 
        n16983, n16982, n16981, n16980, n16979, n16978, n16977, 
        n16976, n16975, n16974, n16973, n16972, n16971, n16970, 
        n16969, n16968, n16967, n16966, n16965, n16964, n16963, 
        n16962, n16961, n16960, n16959, n16958, n16957, n16956, 
        n16955, n16954, n16953, n16952, n16951, n16950, n16949, 
        n16948, n16947, n16946, n16945, n16944, n16943, n16942, 
        n16941, n16940, n16939, n16938, n16937, n16936, n16935, 
        n16934, n16932, n16931, n16930, n16929, n16928, n16927, 
        n16926, n16925, n16924, n16923, n16922, n16921, n16920, 
        n16919, n16918, n16917, n16916, n36_adj_6513, n16915, n16914, 
        n16913, n42_adj_6514, n16912, n45_adj_6515, n16911, n48_adj_6516, 
        n16910, n51_adj_6517, n16909, n54_adj_6518, n16908, n57_adj_6519, 
        n60_adj_6520, n16906, n63_adj_6521, n16905, n66_adj_6522, 
        n16904, n69_adj_6523, n16903, n72_adj_6524, n16902, n75_adj_6525, 
        n16901, n78_adj_6526, n16900, n16899, n16898, n16897, n16896, 
        n16895, n16894, n16893, n16892, n16891, n16890, n16889, 
        n16888, n16887, n16886, n16885, n16884, n16883, n16882, 
        n16881, n16880, n16879, n16878, n16877, n16876, n16875, 
        n16874, n16873, n16872, n16871, n16870, n16869, n16868, 
        n16867, n16866, n16865, n16864, n16862, n16861, n16860, 
        n16859, n16858, n16857, n16856, n16854, n16853, n16852, 
        n16851, n16850, n16849, n16848, n16847, n16846, n16845, 
        n16844, n76_adj_6527, n16843, n79_adj_6528, n16842, n82_adj_6529, 
        n16841, n85_adj_6530, n16840, n88_adj_6531, n16839, n91_adj_6532, 
        n16838, n94_adj_6533, n16837, n97_adj_6534, n16836, n100_adj_6535, 
        n16835, n103_adj_6536, n16834, n106_adj_6537, n16833, n109_adj_6538, 
        n16832, n112_adj_6539, n16831, n115_adj_6540, n16830, n118_adj_6541, 
        n16829, n19628, n16828, n16827, n16826, n16825, n16824, 
        n16823, n16822, n16821, n16820, n16819, n16818, n16817, 
        n16816, n16815, n16814, n16813, n16812, n16810, n16809, 
        n16808, n16807, n16806, n16805, n16804, n16803, n16802, 
        n16801, n16800, n16799, n16798, n16797, n16796, n16795, 
        n16794, n16793, n16792, n16791, n16790, n16789, n16788, 
        n16787, n16786, n16785, n16784, n16783, n16782, n16781, 
        n16780, n16779, n16778, n16777, n16776, n16775, n16774, 
        n16773, n16772, n16771, n16770, n16769, n16768, n16766, 
        n16765, n16764, n16763, n16762, n16761, n16760, n16759, 
        n16758, n16757, n16756, n16755, n16754, n16753, n16752, 
        n16751, n16750, n16749, n16748, n16747, n16746, n16745, 
        n16744, n16743, n16742, n16741, n16740, n16739, n16738, 
        n16737, n16736, n16734, n16733, n16732, n16731, n16730, 
        n16729, n16728, n16727, n16726, n16725, n16724, n16723, 
        n16722, n16721, n16720, n16719, n16718, n16717, n16715, 
        n16714, n16713, n16712, n16711, n16710, n16709, n16707, 
        n16706, n16705, n16704, n16703, n16702, n16701, n16700, 
        n16699, n16698, n16697, n16696, n16695, n16694, n16693, 
        n16692, n16691, n16690, n16686, n16685, n16684, n19664, 
        n16683, n16682, n16681, n16680, n16679, n16678, n16677, 
        n16676, n16675, n16674, n16673, n16672, n16671, n16670, 
        n16669, n19663, n16667, n16666, n16665, n16664, n16663, 
        n16662, n16661, n16660, n16659, n16658, n16657, n16656, 
        n16655, n16654, n16653, n16652, n16651, n16650, n16649, 
        n16648, n16647, n16646, n16645, n16644, n16643, n16642, 
        n16641, n16640, n16639, n16638, n16637, n16636, n16635, 
        n16634, n16633, n16632, n16631, n16630, n16629, n16628, 
        n16627, n16625, n16624, n16623, n16622, n16621, n16620, 
        n16619, n16618, n16617, n16616, n16615, n16614, n16613, 
        n16612, n16611, n16610, n16609, n16608, n16607, n16606, 
        n16605, n16604, n16603, n16602, n16601, n16600, n16599, 
        n16598, n16597, n16596, n16595, n16594, n16593, n16592, 
        n16591, n16590, n16588, n16587, n16586, n16585, n16584, 
        n16583, n16582, n16581, n16580, n16579, n16578, n16577, 
        n16576, n16575, n16574, n16573, n16572, n16571, n16570, 
        n16569, n16568, n16567, n16566, n16565, n16564, n16562, 
        n16561, n16560, n16559, n16558, n16557, n16556, n16554, 
        n16553, n16552, n16551, n16550, n16549, n16548, n16547, 
        n16546, n16545, n16544, n16543, n16542, n16541, n16540, 
        n16539, n16538, n16537, n16536, n16535, n16534, n16533, 
        n16532, n16531, n16530, n16528, n16527, n16526, n16525, 
        n16524, n16523, n16522, n16520, n16519, n16518, n16517, 
        n16516, n16515, n16514, n16512, n16511, n16510, n16509, 
        n16508, n16507, n16506, n16504, n16503, n16502, n16501, 
        n16500, n16499, n16498, n16497, n16496, n16495, n16494, 
        n16493, n16492, n16491, n16490, n16489, n16488, n16487, 
        n16486, n16485, n16484, n16483, n16482, n16481, n16480, 
        n16478, n16477, n16476, n16475, n16474, n16473, n16472, 
        n16471, n19480, n16470, n16469, n16468, n16467, n16466, 
        n16465, n16464, n16463, n16462, n16461, n16459, n16458, 
        n16457, n16456, n16455, n16454, n16453, n16452, n16451, 
        n16450, n16449, n16448, n16447, n16446, n16445, n16444, 
        n16443, n16442, n16440, n16439, n16438, n16437, n16436, 
        n16435, n16434, n16433, n16432, n16431, n16430, n16429, 
        n16428, n16427, n16426, n16425, n16424, n16423, n16421, 
        n16420, n16419, n16418, n16417, n16416, n16415, n16414, 
        n16413, n16412, n16411, n16410, n16409, n16408, n16407, 
        n16406, n16405, n16404, n16403, n16402, n16401, n16400, 
        n16399, n16398, n16397, n16396, n16395, n16394, n16393, 
        n16392, n16391, n16390, n16389, n16388, n16387, n16386, 
        n16384, n16383, n16382, n34_adj_6542, n16381, n16380, n16379, 
        n16378, n16377, n16376, n16375, n16374, n16373, n16372, 
        n16371, n16370, n16369, n16368, n16367, n16365, n16364, 
        n16363, n16362, n16361, n16360, n16359, n16358, n16357, 
        n16356, n16355, n16354, n16353, n16352, n16351, n16350, 
        n16349, n16348, n16345, n16344, n16343, n16342, n16341, 
        n16340, n16339, n16338, n16337, n16336, n16335, n16334, 
        n16333, n16332, n16331, n16330, n16329, n16328, n16324, 
        n16323, n16322, n16321, n16320, n16319, n16318, n16317, 
        n16316, n16315, n16314, n16313, n16312, n16311, n16310, 
        n16309, n16308, n16307, n16305, n16304, n16303, n16302, 
        n16301, n16300, n16299, n16298, n16297, n16296, n16295, 
        n16294, n16293, n16292, n16291, n16290, n16289, n16288, 
        n16283, n16282, n16281, n16280, n16279, n16278, n16277, 
        n16276, n16275, n16274, n16273, n16272, n16271, n16270, 
        n16269, n16268, n16267, n16266, n19479, n16261, n16260, 
        n16259, n16258, n16257, n16256, n16255, n16254, n16253, 
        n16252, n16251, n16250, n16249, n19816, n19815, n19134, 
        n19814, n19474, n19473, n19630, n19472, n19298, cout_adj_6543, 
        n19813, n19812, cout_adj_6544, clk_80mhz_enable_223, n19810, 
        n19808, n19798, n19640, n19797, n19831, n19796, n19795, 
        n19641, n19794, n19811, n19793, n19642, n19791, n19449, 
        n19790, n19789, n19788, n18704, n19787, n19786, n19785, 
        n18700, n19448, n19446, n19445, n19297, n19444, n19647, 
        n19296, n19648, n19443, n19442, n19441, n18600, n18533, 
        n19649, n19806;
    
    VHI i2 (.Z(VCC_net));
    MUX21 i8412 (.D0(n3794), .D1(n3791), .SD(n19822), .Z(n3797));
    CCU2C _add_1_3699_add_4_10 (.A0(amdemod_out_d_11__N_2370[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2370[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16851), .COUT(n16852), 
          .S0(n57_adj_5817), .S1(n54_adj_5816));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3699_add_4_10.INIT0 = 16'h555f;
    defparam _add_1_3699_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_3699_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3699_add_4_10.INJECT1_1 = "NO";
    FD1S3AX rx_byte_i0 (.D(rx_byte1[0]), .CK(clk_80mhz), .Q(rx_byte[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam rx_byte_i0.GSR = "ENABLED";
    CCU2C _add_1_3699_add_4_8 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2370[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2370[4]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16850), .COUT(n16851), 
          .S0(n63_adj_5819), .S1(n60_adj_5818));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3699_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3699_add_4_8.INIT1 = 16'h555f;
    defparam _add_1_3699_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3699_add_4_8.INJECT1_1 = "NO";
    FD1S3AX phase_increment_0__i117 (.D(\phase_increment[0] [52]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [52]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i117.GSR = "ENABLED";
    CCU2C _add_1_3699_add_4_6 (.A0(amdemod_out_d_11__N_2370[1]), .B0(square_sum[25]), 
          .C0(n30_adj_6282), .D0(n13890), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2370[2]), .D1(VCC_net), .CIN(n16849), 
          .COUT(n16850), .S0(n69_adj_5821), .S1(n66_adj_5820));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3699_add_4_6.INIT0 = 16'h596a;
    defparam _add_1_3699_add_4_6.INIT1 = 16'he1e1;
    defparam _add_1_3699_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3699_add_4_6.INJECT1_1 = "NO";
    OB pwm_out_p_pad_3 (.I(pwm_out_p_c), .O(pwm_out_p[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(43[22:31])
    CCU2C _add_1_3699_add_4_4 (.A0(n19816), .B0(square_sum[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_out_d_11__N_2370[0]), .B1(amdemod_out_d_11__N_2370[11]), 
          .C1(amdemod_out_d_11__N_2363), .D1(amdemod_out_d_11__N_2369[11]), 
          .CIN(n16848), .COUT(n16849), .S0(n75_adj_5823), .S1(n72_adj_5822));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3699_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3699_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_3699_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3699_add_4_4.INJECT1_1 = "NO";
    FD1S3AX phase_increment_0__i116 (.D(\phase_increment[0] [51]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i116.GSR = "ENABLED";
    PFUMX mux_1673_i1 (.BLUT(n2989), .ALUT(n2995), .C0(n19299), .Z(n2998));
    quarterwave_generator nco_inst (.clk_80mhz(clk_80mhz), .\phase_accumulator[63] (phase_accumulator_adj_6545[63]), 
            .\lo_sinewave[0] (lo_sinewave[0]), .\lo_cosinewave[0] (lo_cosinewave[0]), 
            .\lo_cosinewave[9] (lo_cosinewave[9]), .\lo_cosinewave[10] (lo_cosinewave[10]), 
            .\lo_sinewave[5] (lo_sinewave[5]), .\lo_cosinewave[6] (lo_cosinewave[6]), 
            .\lo_cosinewave[7] (lo_cosinewave[7]), .\lo_cosinewave[4] (lo_cosinewave[4]), 
            .\lo_cosinewave[5] (lo_cosinewave[5]), .\lo_sinewave[6] (lo_sinewave[6]), 
            .\lo_sinewave[9] (lo_sinewave[9]), .\lo_sinewave[10] (lo_sinewave[10]), 
            .\lo_sinewave[12] (lo_sinewave[12]), .\lo_sinewave[8] (lo_sinewave[8]), 
            .\lo_sinewave[7] (lo_sinewave[7]), .\lo_sinewave[2] (lo_sinewave[2]), 
            .\lo_sinewave[3] (lo_sinewave[3]), .\lo_sinewave[4] (lo_sinewave[4]), 
            .\lo_sinewave[1] (lo_sinewave[1]), .sine_table_value({sine_table_value}), 
            .n67({n28_adj_6326, n31_adj_6327, n34_adj_6328, n37_adj_6329, 
            n40_adj_6330, n43_adj_6331, n46_adj_6332, n49_adj_6333, 
            n52_adj_6334, n55_adj_6335, n58_adj_6336, n61_adj_6337}), 
            .\phase_accumulator[62] (phase_accumulator_adj_6545[62]), .cosine_table_value({cosine_table_value}), 
            .n67_adj_464({n28_adj_6338, n31_adj_6339, n34_adj_6340, n37_adj_6341, 
            n40_adj_6342, n43_adj_6343, n46_adj_6344, n49_adj_6345, 
            n52_adj_6346, n55_adj_6347, n58_adj_6348, n61_adj_6349}), 
            .\phase_accumulator[56] (phase_accumulator_adj_6545[56]), .\phase_accumulator[57] (phase_accumulator_adj_6545[57]), 
            .\phase_accumulator[58] (phase_accumulator_adj_6545[58]), .\phase_accumulator[59] (phase_accumulator_adj_6545[59]), 
            .\phase_accumulator[60] (phase_accumulator_adj_6545[60]), .\phase_accumulator[61] (phase_accumulator_adj_6545[61]), 
            .\lo_cosinewave[12] (lo_cosinewave[12]), .\lo_cosinewave[8] (lo_cosinewave[8]), 
            .\lo_cosinewave[3] (lo_cosinewave[3]), .\lo_cosinewave[2] (lo_cosinewave[2]), 
            .\lo_cosinewave[1] (lo_cosinewave[1]), .GND_net(GND_net), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(158[7] 165[5])
    FD1S3AX phase_accumulator_e3_i0_i41 (.D(n198), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i41.GSR = "ENABLED";
    CCU2C _add_1_3699_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[16]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16848), .S1(n78_adj_5824));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3699_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3699_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3699_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3699_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_38 (.A0(comb_d9[71]), .B0(comb9[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16847), .S0(n78_adj_5825));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3702_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_36 (.A0(comb_d9[69]), .B0(comb9[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[70]), .B1(comb9[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16846), .COUT(n16847), .S0(n84_adj_5827), 
          .S1(n81_adj_5826));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_34 (.A0(comb_d9[67]), .B0(comb9[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[68]), .B1(comb9[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16845), .COUT(n16846), .S0(n90_adj_5829), 
          .S1(n87_adj_5828));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_32 (.A0(comb_d9[65]), .B0(comb9[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[66]), .B1(comb9[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16844), .COUT(n16845), .S0(n96_adj_5831), 
          .S1(n93_adj_5830));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_30 (.A0(comb_d9[63]), .B0(comb9[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[64]), .B1(comb9[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16843), .COUT(n16844), .S0(n102_adj_5833), 
          .S1(n99_adj_5832));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_28 (.A0(comb_d9[61]), .B0(comb9[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[62]), .B1(comb9[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16842), .COUT(n16843), .S0(n108_adj_5835), 
          .S1(n105_adj_5834));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_26 (.A0(comb_d9[59]), .B0(comb9[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[60]), .B1(comb9[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16841), .COUT(n16842), .S0(n114_adj_5837), 
          .S1(n111_adj_5836));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_24 (.A0(comb_d9[57]), .B0(comb9[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[58]), .B1(comb9[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16840), .COUT(n16841), .S0(n120_adj_5839), 
          .S1(n117_adj_5838));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_22 (.A0(comb_d9[55]), .B0(comb9[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[56]), .B1(comb9[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16839), .COUT(n16840));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_20 (.A0(comb_d9[53]), .B0(comb9[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[54]), .B1(comb9[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16838), .COUT(n16839));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_18 (.A0(comb_d9[51]), .B0(comb9[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[52]), .B1(comb9[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16837), .COUT(n16838));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_16 (.A0(comb_d9[49]), .B0(comb9[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[50]), .B1(comb9[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16836), .COUT(n16837));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_14 (.A0(comb_d9[47]), .B0(comb9[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[48]), .B1(comb9[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16835), .COUT(n16836));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_12 (.A0(comb_d9[45]), .B0(comb9[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[46]), .B1(comb9[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16834), .COUT(n16835));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_10 (.A0(comb_d9[43]), .B0(comb9[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[44]), .B1(comb9[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16833), .COUT(n16834));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_8 (.A0(comb_d9[41]), .B0(comb9[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[42]), .B1(comb9[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16832), .COUT(n16833));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3702_add_4_6 (.A0(comb_d9[39]), .B0(comb9[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[40]), .B1(comb9[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16831), .COUT(n16832));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_6.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i40 (.D(n201), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[40]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i40.GSR = "ENABLED";
    CCU2C _add_1_3702_add_4_4 (.A0(comb_d9[37]), .B0(comb9[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[38]), .B1(comb9[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16830), .COUT(n16831));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3702_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_4.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i63 (.D(n132_adj_5305), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i63.GSR = "ENABLED";
    CCU2C _add_1_3702_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[36]), .B1(comb9[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16830));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3702_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3702_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3702_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3702_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_38 (.A0(comb_d7_adj_6566[35]), .B0(comb7_adj_6565[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16829), .S0(comb8_71__N_2137_adj_6591[35]), 
          .S1(cout_adj_5840));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3705_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_36 (.A0(comb_d7_adj_6566[33]), .B0(comb7_adj_6565[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[34]), .B1(comb7_adj_6565[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16828), .COUT(n16829), .S0(comb8_71__N_2137_adj_6591[33]), 
          .S1(comb8_71__N_2137_adj_6591[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_34 (.A0(comb_d7_adj_6566[31]), .B0(comb7_adj_6565[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[32]), .B1(comb7_adj_6565[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16827), .COUT(n16828), .S0(comb8_71__N_2137_adj_6591[31]), 
          .S1(comb8_71__N_2137_adj_6591[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_32 (.A0(comb_d7_adj_6566[29]), .B0(comb7_adj_6565[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[30]), .B1(comb7_adj_6565[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16826), .COUT(n16827), .S0(comb8_71__N_2137_adj_6591[29]), 
          .S1(comb8_71__N_2137_adj_6591[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_30 (.A0(comb_d7_adj_6566[27]), .B0(comb7_adj_6565[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[28]), .B1(comb7_adj_6565[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16825), .COUT(n16826), .S0(comb8_71__N_2137_adj_6591[27]), 
          .S1(comb8_71__N_2137_adj_6591[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_28 (.A0(comb_d7_adj_6566[25]), .B0(comb7_adj_6565[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[26]), .B1(comb7_adj_6565[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16824), .COUT(n16825), .S0(comb8_71__N_2137_adj_6591[25]), 
          .S1(comb8_71__N_2137_adj_6591[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_26 (.A0(comb_d7_adj_6566[23]), .B0(comb7_adj_6565[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[24]), .B1(comb7_adj_6565[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16823), .COUT(n16824), .S0(comb8_71__N_2137_adj_6591[23]), 
          .S1(comb8_71__N_2137_adj_6591[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_24 (.A0(comb_d7_adj_6566[21]), .B0(comb7_adj_6565[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[22]), .B1(comb7_adj_6565[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16822), .COUT(n16823), .S0(comb8_71__N_2137_adj_6591[21]), 
          .S1(comb8_71__N_2137_adj_6591[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_22 (.A0(comb_d7_adj_6566[19]), .B0(comb7_adj_6565[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[20]), .B1(comb7_adj_6565[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16821), .COUT(n16822), .S0(comb8_71__N_2137_adj_6591[19]), 
          .S1(comb8_71__N_2137_adj_6591[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_20 (.A0(comb_d7_adj_6566[17]), .B0(comb7_adj_6565[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[18]), .B1(comb7_adj_6565[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16820), .COUT(n16821), .S0(comb8_71__N_2137_adj_6591[17]), 
          .S1(comb8_71__N_2137_adj_6591[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_18 (.A0(comb_d7_adj_6566[15]), .B0(comb7_adj_6565[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[16]), .B1(comb7_adj_6565[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16819), .COUT(n16820), .S0(comb8_71__N_2137_adj_6591[15]), 
          .S1(comb8_71__N_2137_adj_6591[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_16 (.A0(comb_d7_adj_6566[13]), .B0(comb7_adj_6565[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[14]), .B1(comb7_adj_6565[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16818), .COUT(n16819), .S0(comb8_71__N_2137_adj_6591[13]), 
          .S1(comb8_71__N_2137_adj_6591[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_14 (.A0(comb_d7_adj_6566[11]), .B0(comb7_adj_6565[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[12]), .B1(comb7_adj_6565[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16817), .COUT(n16818), .S0(comb8_71__N_2137_adj_6591[11]), 
          .S1(comb8_71__N_2137_adj_6591[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3639_add_4_16 (.A0(amdemod_out_d_11__N_2390[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2390[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17277), .S1(n36_adj_6513));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3639_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_3639_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3639_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3639_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_24 (.A0(integrator2[57]), .B0(integrator1[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[58]), .B1(integrator1[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17840), .COUT(n17841), .S0(n120_adj_5315), 
          .S1(n117_adj_5316));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_22 (.A0(integrator2[55]), .B0(integrator1[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[56]), .B1(integrator1[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17839), .COUT(n17840), .S0(n126_adj_5338), 
          .S1(n123_adj_5342));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_12 (.A0(comb_d7_adj_6566[9]), .B0(comb7_adj_6565[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[10]), .B1(comb7_adj_6565[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16816), .COUT(n16817), .S0(comb8_71__N_2137_adj_6591[9]), 
          .S1(comb8_71__N_2137_adj_6591[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_10 (.A0(comb_d7_adj_6566[7]), .B0(comb7_adj_6565[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[8]), .B1(comb7_adj_6565[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16815), .COUT(n16816), .S0(comb8_71__N_2137_adj_6591[7]), 
          .S1(comb8_71__N_2137_adj_6591[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_20 (.A0(integrator2[53]), .B0(integrator1[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[54]), .B1(integrator1[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17838), .COUT(n17839), .S0(n132_adj_5311), 
          .S1(n129_adj_5312));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_18 (.A0(integrator2[51]), .B0(integrator1[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[52]), .B1(integrator1[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17837), .COUT(n17838), .S0(n138_adj_5345), 
          .S1(n135_adj_5343));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_16 (.A0(integrator2[49]), .B0(integrator1[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[50]), .B1(integrator1[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17836), .COUT(n17837), .S0(n144_adj_5348), 
          .S1(n141));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_14 (.A0(integrator2[47]), .B0(integrator1[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[48]), .B1(integrator1[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17835), .COUT(n17836), .S0(n150_adj_5346), 
          .S1(n147_adj_5344));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_12 (.A0(integrator2[45]), .B0(integrator1[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[46]), .B1(integrator1[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17834), .COUT(n17835), .S0(n156_adj_5352), 
          .S1(n153_adj_5349));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_10 (.A0(integrator2[43]), .B0(integrator1[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[44]), .B1(integrator1[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17833), .COUT(n17834), .S0(n162_adj_5309), 
          .S1(n159_adj_5307));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_8 (.A0(integrator2[41]), .B0(integrator1[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[42]), .B1(integrator1[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17832), .COUT(n17833), .S0(n168_adj_5350), 
          .S1(n165_adj_5347));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_6 (.A0(integrator2[39]), .B0(integrator1[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[40]), .B1(integrator1[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17831), .COUT(n17832), .S0(n174_adj_5303), 
          .S1(n171_adj_5306));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_4 (.A0(integrator2[37]), .B0(integrator1[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[38]), .B1(integrator1[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17830), .COUT(n17831), .S0(n180_adj_5325), 
          .S1(n177_adj_5351));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3639_add_4_14 (.A0(amdemod_out_d_11__N_2390[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2390[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17276), .COUT(n17277), 
          .S0(n45_adj_6515), .S1(n42_adj_6514));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3639_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_3639_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_3639_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3639_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator2[36]), .B1(integrator1[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17830), .S1(n183_adj_5324));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3525_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3762_add_4_15 (.A0(amdemod_out_d_11__N_2370[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2370[11]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17828), .S1(n34_adj_6171));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3762_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3762_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3762_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3762_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3639_add_4_12 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2390[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2390[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17275), .COUT(n17276), 
          .S0(n51_adj_6517), .S1(n48_adj_6516));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3639_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3639_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_3639_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3639_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3639_add_4_10 (.A0(amdemod_out_d_11__N_2390[5]), .B0(square_sum[25]), 
          .C0(n30_adj_6282), .D0(n13890), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2390[6]), .D1(VCC_net), .CIN(n17274), 
          .COUT(n17275), .S0(n57_adj_6519), .S1(n54_adj_6518));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3639_add_4_10.INIT0 = 16'h596a;
    defparam _add_1_3639_add_4_10.INIT1 = 16'he1e1;
    defparam _add_1_3639_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3639_add_4_10.INJECT1_1 = "NO";
    LUT4 i8271_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19449), 
         .D(n1616), .Z(n1632)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8271_3_lut_4_lut.init = 16'hf780;
    CCU2C _add_1_3639_add_4_8 (.A0(n19815), .B0(amdemod_out_d_11__N_2390[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2390[4]), 
          .B1(amdemod_out_d_11__N_2370[11]), .C1(amdemod_out_d_11__N_2363), 
          .D1(amdemod_out_d_11__N_2369[11]), .CIN(n17273), .COUT(n17274), 
          .S0(n63_adj_6521), .S1(n60_adj_6520));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3639_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3639_add_4_8.INIT1 = 16'h656a;
    defparam _add_1_3639_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3639_add_4_8.INJECT1_1 = "NO";
    LUT4 i8166_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19474), 
         .D(n2744), .Z(n2760)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8166_3_lut_4_lut.init = 16'hf780;
    PFUMX i8576 (.BLUT(n19602), .ALUT(n19601), .C0(rx_byte[2]), .Z(n19603));
    CCU2C _add_1_3762_add_4_13 (.A0(amdemod_out_d_11__N_2370[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2370[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17827), .COUT(n17828), 
          .S0(n43_adj_6173), .S1(n40_adj_6172));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3762_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3762_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3762_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3762_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3639_add_4_6 (.A0(n19813), .B0(amdemod_out_d_11__N_2390[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2390[2]), 
          .B1(amdemod_out_d_11__N_2380[14]), .C1(n19815), .D1(amdemod_out_d_11__N_2379[14]), 
          .CIN(n17272), .COUT(n17273), .S0(n69_adj_6523), .S1(n66_adj_6522));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3639_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3639_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_3639_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3639_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3762_add_4_11 (.A0(amdemod_out_d_11__N_2370[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2370[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17826), .COUT(n17827), 
          .S0(n49_adj_6175), .S1(n46_adj_6174));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3762_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3762_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3762_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3762_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_33 (.A0(\phase_increment[0] [32]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [33]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17614), .COUT(n17615), .S0(phase_increment_1__63__N_20[32]), 
          .S1(phase_increment_1__63__N_20[33]));
    defparam _add_1_3813_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3762_add_4_9 (.A0(amdemod_out_d_11__N_2370[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2370[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17825), .COUT(n17826), 
          .S0(n55_adj_6177), .S1(n52_adj_6176));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3762_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_3762_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_3762_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3762_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3639_add_4_4 (.A0(n19812), .B0(square_sum[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_out_d_11__N_2390[0]), .B1(amdemod_out_d_11__N_2390[14]), 
          .C1(n19813), .D1(amdemod_out_d_11__N_2389[14]), .CIN(n17271), 
          .COUT(n17272), .S0(n75_adj_6525), .S1(n72_adj_6524));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3639_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3639_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_3639_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3639_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3639_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17271), .S1(n78_adj_6526));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3639_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3639_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3639_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3639_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3762_add_4_7 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2370[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2370[4]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17824), .COUT(n17825), 
          .S0(n61_adj_6179), .S1(n58_adj_6178));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3762_add_4_7.INIT0 = 16'h666a;
    defparam _add_1_3762_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_3762_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3762_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3762_add_4_5 (.A0(amdemod_out_d_11__N_2363), .B0(amdemod_out_d_11__N_2370[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2370[2]), .D1(VCC_net), .CIN(n17823), 
          .COUT(n17824), .S0(n67_adj_6181), .S1(n64_adj_6180));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3762_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3762_add_4_5.INIT1 = 16'h1e1e;
    defparam _add_1_3762_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3762_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3762_add_4_3 (.A0(square_sum[17]), .B0(amdemod_out_d_11__N_2370[11]), 
          .C0(amdemod_out_d_11__N_2363), .D0(amdemod_out_d_11__N_2369[11]), 
          .A1(n19816), .B1(amdemod_out_d_11__N_2370[0]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17822), .COUT(n17823), .S0(n73_adj_6183), 
          .S1(n70_adj_6182));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3762_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_3762_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3762_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3762_add_4_3.INJECT1_1 = "NO";
    LUT4 i1_4_lut_then_4_lut (.A(rx_byte[4]), .B(rx_byte[0]), .C(rx_byte[3]), 
         .D(rx_byte[2]), .Z(n19863)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0400;
    CCU2C _add_1_3762_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[16]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17822), .S1(n76_adj_6184));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3762_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3762_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3762_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3762_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_else_4_lut (.A(rx_byte[4]), .B(rx_byte[0]), .C(rx_byte[3]), 
         .D(rx_byte[2]), .Z(n19862)) /* synthesis lut_function=(!(A+!(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h4014;
    FD1S3AX phase_accumulator_e3_i0_i62 (.D(n135_adj_5287), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[62]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i62.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i61 (.D(n138_adj_5292), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i61.GSR = "ENABLED";
    FD1S3AX rx_data_valid_255 (.D(rx_data_valid1), .CK(clk_80mhz), .Q(rx_data_valid));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam rx_data_valid_255.GSR = "ENABLED";
    CCU2C _add_1_3765_add_4_37 (.A0(integrator4[70]), .B0(cout_adj_5293), 
          .C0(n81_adj_6001), .D0(integrator5[70]), .A1(integrator4[71]), 
          .B1(cout_adj_5293), .C1(n78_adj_6000), .D1(integrator5[71]), 
          .CIN(n17820), .S0(integrator5_71__N_1248[70]), .S1(integrator5_71__N_1248[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_35 (.A0(integrator4[68]), .B0(cout_adj_5293), 
          .C0(n87_adj_6003), .D0(integrator5[68]), .A1(integrator4[69]), 
          .B1(cout_adj_5293), .C1(n84_adj_6002), .D1(integrator5[69]), 
          .CIN(n17819), .COUT(n17820), .S0(integrator5_71__N_1248[68]), 
          .S1(integrator5_71__N_1248[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_33 (.A0(integrator4[66]), .B0(cout_adj_5293), 
          .C0(n93_adj_6005), .D0(integrator5[66]), .A1(integrator4[67]), 
          .B1(cout_adj_5293), .C1(n90_adj_6004), .D1(integrator5[67]), 
          .CIN(n17818), .COUT(n17819), .S0(integrator5_71__N_1248[66]), 
          .S1(integrator5_71__N_1248[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_31 (.A0(integrator4[64]), .B0(cout_adj_5293), 
          .C0(n99_adj_6007), .D0(integrator5[64]), .A1(integrator4[65]), 
          .B1(cout_adj_5293), .C1(n96_adj_6006), .D1(integrator5[65]), 
          .CIN(n17817), .COUT(n17818), .S0(integrator5_71__N_1248[64]), 
          .S1(integrator5_71__N_1248[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_29 (.A0(integrator4[62]), .B0(cout_adj_5293), 
          .C0(n105_adj_6009), .D0(integrator5[62]), .A1(integrator4[63]), 
          .B1(cout_adj_5293), .C1(n102_adj_6008), .D1(integrator5[63]), 
          .CIN(n17816), .COUT(n17817), .S0(integrator5_71__N_1248[62]), 
          .S1(integrator5_71__N_1248[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_27 (.A0(integrator4[60]), .B0(cout_adj_5293), 
          .C0(n111_adj_6011), .D0(integrator5[60]), .A1(integrator4[61]), 
          .B1(cout_adj_5293), .C1(n108_adj_6010), .D1(integrator5[61]), 
          .CIN(n17815), .COUT(n17816), .S0(integrator5_71__N_1248[60]), 
          .S1(integrator5_71__N_1248[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_25 (.A0(integrator4[58]), .B0(cout_adj_5293), 
          .C0(n117_adj_6013), .D0(integrator5[58]), .A1(integrator4[59]), 
          .B1(cout_adj_5293), .C1(n114_adj_6012), .D1(integrator5[59]), 
          .CIN(n17814), .COUT(n17815), .S0(integrator5_71__N_1248[58]), 
          .S1(integrator5_71__N_1248[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_23 (.A0(integrator4[56]), .B0(cout_adj_5293), 
          .C0(n123_adj_6015), .D0(integrator5[56]), .A1(integrator4[57]), 
          .B1(cout_adj_5293), .C1(n120_adj_6014), .D1(integrator5[57]), 
          .CIN(n17813), .COUT(n17814), .S0(integrator5_71__N_1248[56]), 
          .S1(integrator5_71__N_1248[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_21 (.A0(integrator4[54]), .B0(cout_adj_5293), 
          .C0(n129_adj_6017), .D0(integrator5[54]), .A1(integrator4[55]), 
          .B1(cout_adj_5293), .C1(n126_adj_6016), .D1(integrator5[55]), 
          .CIN(n17812), .COUT(n17813), .S0(integrator5_71__N_1248[54]), 
          .S1(integrator5_71__N_1248[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_19 (.A0(integrator4[52]), .B0(cout_adj_5293), 
          .C0(n135_adj_6019), .D0(integrator5[52]), .A1(integrator4[53]), 
          .B1(cout_adj_5293), .C1(n132_adj_6018), .D1(integrator5[53]), 
          .CIN(n17811), .COUT(n17812), .S0(integrator5_71__N_1248[52]), 
          .S1(integrator5_71__N_1248[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_17 (.A0(integrator4[50]), .B0(cout_adj_5293), 
          .C0(n141_adj_6021), .D0(integrator5[50]), .A1(integrator4[51]), 
          .B1(cout_adj_5293), .C1(n138_adj_6020), .D1(integrator5[51]), 
          .CIN(n17810), .COUT(n17811), .S0(integrator5_71__N_1248[50]), 
          .S1(integrator5_71__N_1248[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_15 (.A0(integrator4[48]), .B0(cout_adj_5293), 
          .C0(n147_adj_6023), .D0(integrator5[48]), .A1(integrator4[49]), 
          .B1(cout_adj_5293), .C1(n144_adj_6022), .D1(integrator5[49]), 
          .CIN(n17809), .COUT(n17810), .S0(integrator5_71__N_1248[48]), 
          .S1(integrator5_71__N_1248[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_13 (.A0(integrator4[46]), .B0(cout_adj_5293), 
          .C0(n153_adj_6025), .D0(integrator5[46]), .A1(integrator4[47]), 
          .B1(cout_adj_5293), .C1(n150_adj_6024), .D1(integrator5[47]), 
          .CIN(n17808), .COUT(n17809), .S0(integrator5_71__N_1248[46]), 
          .S1(integrator5_71__N_1248[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_11 (.A0(integrator4[44]), .B0(cout_adj_5293), 
          .C0(n159_adj_6027), .D0(integrator5[44]), .A1(integrator4[45]), 
          .B1(cout_adj_5293), .C1(n156_adj_6026), .D1(integrator5[45]), 
          .CIN(n17807), .COUT(n17808), .S0(integrator5_71__N_1248[44]), 
          .S1(integrator5_71__N_1248[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_9 (.A0(integrator4[42]), .B0(cout_adj_5293), 
          .C0(n165_adj_6029), .D0(integrator5[42]), .A1(integrator4[43]), 
          .B1(cout_adj_5293), .C1(n162_adj_6028), .D1(integrator5[43]), 
          .CIN(n17806), .COUT(n17807), .S0(integrator5_71__N_1248[42]), 
          .S1(integrator5_71__N_1248[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_7 (.A0(integrator4[40]), .B0(cout_adj_5293), 
          .C0(n171_adj_6031), .D0(integrator5[40]), .A1(integrator4[41]), 
          .B1(cout_adj_5293), .C1(n168_adj_6030), .D1(integrator5[41]), 
          .CIN(n17805), .COUT(n17806), .S0(integrator5_71__N_1248[40]), 
          .S1(integrator5_71__N_1248[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_5 (.A0(integrator4[38]), .B0(cout_adj_5293), 
          .C0(n177_adj_6033), .D0(integrator5[38]), .A1(integrator4[39]), 
          .B1(cout_adj_5293), .C1(n174_adj_6032), .D1(integrator5[39]), 
          .CIN(n17804), .COUT(n17805), .S0(integrator5_71__N_1248[38]), 
          .S1(integrator5_71__N_1248[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_3 (.A0(integrator4[36]), .B0(cout_adj_5293), 
          .C0(n183_adj_6035), .D0(integrator5[36]), .A1(integrator4[37]), 
          .B1(cout_adj_5293), .C1(n180_adj_6034), .D1(integrator5[37]), 
          .CIN(n17803), .COUT(n17804), .S0(integrator5_71__N_1248[36]), 
          .S1(integrator5_71__N_1248[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3765_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3765_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5293), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17803));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3765_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3765_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3765_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3768_add_4_16 (.A0(amdemod_out_d_11__N_2801), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2798), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17798), .S1(amdemod_out_d_11__N_2409[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3768_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_3768_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3768_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3768_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3768_add_4_14 (.A0(square_sum[25]), .B0(n19824), .C0(amdemod_out_d_11__N_2807), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(amdemod_out_d_11__N_2804), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17797), .COUT(n17798), .S0(amdemod_out_d_11__N_2409[11]), 
          .S1(amdemod_out_d_11__N_2409[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3768_add_4_14.INIT0 = 16'he1e1;
    defparam _add_1_3768_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3768_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3768_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3768_add_4_12 (.A0(amdemod_out_d_11__N_2813), .B0(amdemod_out_d_11__N_2370[11]), 
          .C0(amdemod_out_d_11__N_2363), .D0(amdemod_out_d_11__N_2369[11]), 
          .A1(amdemod_out_d_11__N_2810), .B1(square_sum[25]), .C1(n30_adj_6282), 
          .D1(n13890), .CIN(n17796), .COUT(n17797), .S0(amdemod_out_d_11__N_2409[9]), 
          .S1(amdemod_out_d_11__N_2409[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3768_add_4_12.INIT0 = 16'h656a;
    defparam _add_1_3768_add_4_12.INIT1 = 16'h596a;
    defparam _add_1_3768_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3768_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3768_add_4_10 (.A0(amdemod_out_d_11__N_2819), .B0(amdemod_out_d_11__N_2380[14]), 
          .C0(n19815), .D0(amdemod_out_d_11__N_2379[14]), .A1(n19815), 
          .B1(amdemod_out_d_11__N_2816), .C1(GND_net), .D1(VCC_net), .CIN(n17795), 
          .COUT(n17796), .S0(amdemod_out_d_11__N_2409[7]), .S1(amdemod_out_d_11__N_2409[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3768_add_4_10.INIT0 = 16'h656a;
    defparam _add_1_3768_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3768_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3768_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3768_add_4_8 (.A0(amdemod_out_d_11__N_2825), .B0(amdemod_out_d_11__N_2390[14]), 
          .C0(n19813), .D0(amdemod_out_d_11__N_2389[14]), .A1(n19813), 
          .B1(amdemod_out_d_11__N_2822), .C1(GND_net), .D1(VCC_net), .CIN(n17794), 
          .COUT(n17795), .S0(amdemod_out_d_11__N_2409[5]), .S1(amdemod_out_d_11__N_2409[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3768_add_4_8.INIT0 = 16'h656a;
    defparam _add_1_3768_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3768_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3768_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3768_add_4_6 (.A0(amdemod_out_d_11__N_2831), .B0(amdemod_out_d_11__N_2400[14]), 
          .C0(n19811), .D0(amdemod_out_d_11__N_2399[14]), .A1(n19811), 
          .B1(amdemod_out_d_11__N_2828), .C1(GND_net), .D1(VCC_net), .CIN(n17793), 
          .COUT(n17794), .S0(amdemod_out_d_11__N_2409[3]), .S1(amdemod_out_d_11__N_2409[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3768_add_4_6.INIT0 = 16'h656a;
    defparam _add_1_3768_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3768_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3768_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3768_add_4_4 (.A0(n19809), .B0(square_sum[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19809), .B1(amdemod_out_d_11__N_2834), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17792), .COUT(n17793), .S0(amdemod_out_d_11__N_2409[1]), 
          .S1(amdemod_out_d_11__N_2409[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3768_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3768_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3768_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3768_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3768_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17792), .S1(amdemod_out_d_11__N_2409[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3768_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3768_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3768_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3768_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3774_add_4_15 (.A0(amdemod_out_d_11__N_2369[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2369[11]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17790), .S1(n34_adj_6185));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3774_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3774_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3774_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3774_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3774_add_4_13 (.A0(amdemod_out_d_11__N_2369[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2369[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17789), .COUT(n17790), 
          .S0(n43_adj_6187), .S1(n40_adj_6186));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3774_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3774_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3774_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3774_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3774_add_4_11 (.A0(amdemod_out_d_11__N_2369[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2369[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17788), .COUT(n17789), 
          .S0(n49_adj_6189), .S1(n46_adj_6188));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3774_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3774_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3774_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3774_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3774_add_4_9 (.A0(amdemod_out_d_11__N_2369[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2369[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17787), .COUT(n17788), 
          .S0(n55_adj_6191), .S1(n52_adj_6190));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3774_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_3774_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_3774_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3774_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3774_add_4_7 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2369[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2369[4]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17786), .COUT(n17787), 
          .S0(n61_adj_6193), .S1(n58_adj_6192));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3774_add_4_7.INIT0 = 16'h666a;
    defparam _add_1_3774_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_3774_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3774_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3774_add_4_5 (.A0(amdemod_out_d_11__N_2363), .B0(amdemod_out_d_11__N_2369[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2369[2]), .D1(VCC_net), .CIN(n17785), 
          .COUT(n17786), .S0(n67_adj_6195), .S1(n64_adj_6194));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3774_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3774_add_4_5.INIT1 = 16'h1e1e;
    defparam _add_1_3774_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3774_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3774_add_4_3 (.A0(square_sum[17]), .B0(amdemod_out_d_11__N_2370[11]), 
          .C0(amdemod_out_d_11__N_2363), .D0(amdemod_out_d_11__N_2369[11]), 
          .A1(n19816), .B1(amdemod_out_d_11__N_2369[0]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17784), .COUT(n17785), .S0(n73_adj_6197), 
          .S1(n70_adj_6196));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3774_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_3774_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3774_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3774_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3774_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[16]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17784), .S1(n76_adj_6198));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3774_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3774_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3774_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3774_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3777_add_4_9 (.A0(square_sum[25]), .B0(n19824), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17782), .S0(amdemod_out_d_11__N_2365[7]), 
          .S1(amdemod_out_d_11__N_2365[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3777_add_4_9.INIT0 = 16'h1111;
    defparam _add_1_3777_add_4_9.INIT1 = 16'h1111;
    defparam _add_1_3777_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3777_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3777_add_4_7 (.A0(n19828), .B0(n19827), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17781), .COUT(n17782), .S0(amdemod_out_d_11__N_2365[5]), 
          .S1(amdemod_out_d_11__N_2365[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3777_add_4_7.INIT0 = 16'h1111;
    defparam _add_1_3777_add_4_7.INIT1 = 16'h9999;
    defparam _add_1_3777_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3777_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3777_add_4_5 (.A0(square_sum[25]), .B0(n4_adj_6510), .C0(GND_net), 
          .D0(VCC_net), .A1(n19828), .B1(n19827), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17780), .COUT(n17781), .S0(amdemod_out_d_11__N_2365[3]), 
          .S1(amdemod_out_d_11__N_2365[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3777_add_4_5.INIT0 = 16'h3339;
    defparam _add_1_3777_add_4_5.INIT1 = 16'h1111;
    defparam _add_1_3777_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3777_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3777_add_4_3 (.A0(square_sum[25]), .B0(n19824), .C0(square_sum[21]), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), .C1(square_sum[22]), 
          .D1(VCC_net), .CIN(n17779), .COUT(n17780), .S0(amdemod_out_d_11__N_2365[1]), 
          .S1(amdemod_out_d_11__N_2365[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3777_add_4_3.INIT0 = 16'he1e1;
    defparam _add_1_3777_add_4_3.INIT1 = 16'he1ee;
    defparam _add_1_3777_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3777_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3777_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[20]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17779), .S1(n46_adj_6199));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3777_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3777_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3777_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3777_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_37 (.A0(integrator1_adj_6558[70]), .B0(cout_adj_5328), 
          .C0(n81_adj_5267), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[71]), 
          .B1(cout_adj_5328), .C1(n78_adj_5268), .D1(mix_cosinewave[11]), 
          .CIN(n17777), .S0(integrator1_71__N_960_adj_6573[70]), .S1(integrator1_71__N_960_adj_6573[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_35 (.A0(integrator1_adj_6558[68]), .B0(cout_adj_5328), 
          .C0(n87_adj_5265), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[69]), 
          .B1(cout_adj_5328), .C1(n84_adj_5266), .D1(mix_cosinewave[11]), 
          .CIN(n17776), .COUT(n17777), .S0(integrator1_71__N_960_adj_6573[68]), 
          .S1(integrator1_71__N_960_adj_6573[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_33 (.A0(integrator1_adj_6558[66]), .B0(cout_adj_5328), 
          .C0(n93), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[67]), 
          .B1(cout_adj_5328), .C1(n90_adj_5264), .D1(mix_cosinewave[11]), 
          .CIN(n17775), .COUT(n17776), .S0(integrator1_71__N_960_adj_6573[66]), 
          .S1(integrator1_71__N_960_adj_6573[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_31 (.A0(integrator1_adj_6558[64]), .B0(cout_adj_5328), 
          .C0(n99), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[65]), 
          .B1(cout_adj_5328), .C1(n96), .D1(mix_cosinewave[11]), .CIN(n17774), 
          .COUT(n17775), .S0(integrator1_71__N_960_adj_6573[64]), .S1(integrator1_71__N_960_adj_6573[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_29 (.A0(integrator1_adj_6558[62]), .B0(cout_adj_5328), 
          .C0(n105), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[63]), 
          .B1(cout_adj_5328), .C1(n102), .D1(mix_cosinewave[11]), .CIN(n17773), 
          .COUT(n17774), .S0(integrator1_71__N_960_adj_6573[62]), .S1(integrator1_71__N_960_adj_6573[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_27 (.A0(integrator1_adj_6558[60]), .B0(cout_adj_5328), 
          .C0(n111), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[61]), 
          .B1(cout_adj_5328), .C1(n108), .D1(mix_cosinewave[11]), .CIN(n17772), 
          .COUT(n17773), .S0(integrator1_71__N_960_adj_6573[60]), .S1(integrator1_71__N_960_adj_6573[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_25 (.A0(integrator1_adj_6558[58]), .B0(cout_adj_5328), 
          .C0(n117), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[59]), 
          .B1(cout_adj_5328), .C1(n114), .D1(mix_cosinewave[11]), .CIN(n17771), 
          .COUT(n17772), .S0(integrator1_71__N_960_adj_6573[58]), .S1(integrator1_71__N_960_adj_6573[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_23 (.A0(integrator1_adj_6558[56]), .B0(cout_adj_5328), 
          .C0(n123), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[57]), 
          .B1(cout_adj_5328), .C1(n120), .D1(mix_cosinewave[11]), .CIN(n17770), 
          .COUT(n17771), .S0(integrator1_71__N_960_adj_6573[56]), .S1(integrator1_71__N_960_adj_6573[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_21 (.A0(integrator1_adj_6558[54]), .B0(cout_adj_5328), 
          .C0(n129), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[55]), 
          .B1(cout_adj_5328), .C1(n126), .D1(mix_cosinewave[11]), .CIN(n17769), 
          .COUT(n17770), .S0(integrator1_71__N_960_adj_6573[54]), .S1(integrator1_71__N_960_adj_6573[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_19 (.A0(integrator1_adj_6558[52]), .B0(cout_adj_5328), 
          .C0(n135), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[53]), 
          .B1(cout_adj_5328), .C1(n132), .D1(mix_cosinewave[11]), .CIN(n17768), 
          .COUT(n17769), .S0(integrator1_71__N_960_adj_6573[52]), .S1(integrator1_71__N_960_adj_6573[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_17 (.A0(integrator1_adj_6558[50]), .B0(cout_adj_5328), 
          .C0(n141_adj_4975), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[51]), 
          .B1(cout_adj_5328), .C1(n138), .D1(mix_cosinewave[11]), .CIN(n17767), 
          .COUT(n17768), .S0(integrator1_71__N_960_adj_6573[50]), .S1(integrator1_71__N_960_adj_6573[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_15 (.A0(integrator1_adj_6558[48]), .B0(cout_adj_5328), 
          .C0(n147), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[49]), 
          .B1(cout_adj_5328), .C1(n144), .D1(mix_cosinewave[11]), .CIN(n17766), 
          .COUT(n17767), .S0(integrator1_71__N_960_adj_6573[48]), .S1(integrator1_71__N_960_adj_6573[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_13 (.A0(integrator1_adj_6558[46]), .B0(cout_adj_5328), 
          .C0(n153), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[47]), 
          .B1(cout_adj_5328), .C1(n150), .D1(mix_cosinewave[11]), .CIN(n17765), 
          .COUT(n17766), .S0(integrator1_71__N_960_adj_6573[46]), .S1(integrator1_71__N_960_adj_6573[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_11 (.A0(integrator1_adj_6558[44]), .B0(cout_adj_5328), 
          .C0(n159), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[45]), 
          .B1(cout_adj_5328), .C1(n156), .D1(mix_cosinewave[11]), .CIN(n17764), 
          .COUT(n17765), .S0(integrator1_71__N_960_adj_6573[44]), .S1(integrator1_71__N_960_adj_6573[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_9 (.A0(integrator1_adj_6558[42]), .B0(cout_adj_5328), 
          .C0(n165), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[43]), 
          .B1(cout_adj_5328), .C1(n162), .D1(mix_cosinewave[11]), .CIN(n17763), 
          .COUT(n17764), .S0(integrator1_71__N_960_adj_6573[42]), .S1(integrator1_71__N_960_adj_6573[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_7 (.A0(integrator1_adj_6558[40]), .B0(cout_adj_5328), 
          .C0(n171), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[41]), 
          .B1(cout_adj_5328), .C1(n168), .D1(mix_cosinewave[11]), .CIN(n17762), 
          .COUT(n17763), .S0(integrator1_71__N_960_adj_6573[40]), .S1(integrator1_71__N_960_adj_6573[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_5 (.A0(integrator1_adj_6558[38]), .B0(cout_adj_5328), 
          .C0(n177), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[39]), 
          .B1(cout_adj_5328), .C1(n174), .D1(mix_cosinewave[11]), .CIN(n17761), 
          .COUT(n17762), .S0(integrator1_71__N_960_adj_6573[38]), .S1(integrator1_71__N_960_adj_6573[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_3 (.A0(integrator1_adj_6558[36]), .B0(cout_adj_5328), 
          .C0(n183), .D0(mix_cosinewave[11]), .A1(integrator1_adj_6558[37]), 
          .B1(cout_adj_5328), .C1(n180), .D1(mix_cosinewave[11]), .CIN(n17760), 
          .COUT(n17761), .S0(integrator1_71__N_960_adj_6573[36]), .S1(integrator1_71__N_960_adj_6573[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3780_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3780_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3780_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5328), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17760));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3780_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3780_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3780_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3780_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_38 (.A0(mix_sinewave[11]), .B0(integrator1[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17756), .S0(n78_adj_6201));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3792_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_36 (.A0(mix_sinewave[11]), .B0(integrator1[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17755), .COUT(n17756), .S0(n84_adj_6203), 
          .S1(n81_adj_6202));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_8 (.A0(comb_d7_adj_6566[5]), .B0(comb7_adj_6565[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[6]), .B1(comb7_adj_6565[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16814), .COUT(n16815), .S0(comb8_71__N_2137_adj_6591[5]), 
          .S1(comb8_71__N_2137_adj_6591[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_8.INJECT1_1 = "NO";
    LUT4 i4985_2_lut_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[19]), 
         .Z(n3501)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i4985_2_lut_2_lut.init = 16'h4444;
    CCU2C _add_1_3705_add_4_6 (.A0(comb_d7_adj_6566[3]), .B0(comb7_adj_6565[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[4]), .B1(comb7_adj_6565[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16813), .COUT(n16814), .S0(comb8_71__N_2137_adj_6591[3]), 
          .S1(comb8_71__N_2137_adj_6591[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_4 (.A0(comb_d7_adj_6566[1]), .B0(comb7_adj_6565[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[2]), .B1(comb7_adj_6565[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16812), .COUT(n16813), .S0(comb8_71__N_2137_adj_6591[1]), 
          .S1(comb8_71__N_2137_adj_6591[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3705_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_4.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_59__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[59]), .Z(n19448)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_59__bdd_2_lut_2_lut.init = 16'h4444;
    CCU2C _add_1_3642_add_4_37 (.A0(comb_d9[71]), .B0(comb9[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17270), .S0(n76_adj_6527));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_37.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_37.INIT1 = 16'h0000;
    defparam _add_1_3642_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_37.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_4__bdd_4_lut_4_lut (.A(rx_byte[0]), .B(rx_byte[2]), 
         .C(n19799), .D(phase_increment_1__63__N_21[4]), .Z(n19807)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_4__bdd_4_lut_4_lut.init = 16'hd1c0;
    CCU2C _add_1_3642_add_4_35 (.A0(comb_d9[69]), .B0(comb9[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[70]), .B1(comb9[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17269), .COUT(n17270), .S0(n82_adj_6529), 
          .S1(n79_adj_6528));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_35.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_35.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3705_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7_adj_6566[0]), .B1(comb7_adj_6565[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16812), .S1(comb8_71__N_2137_adj_6591[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3705_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3705_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3705_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3705_add_4_2.INJECT1_1 = "NO";
    LUT4 mux_1122_i1_3_lut (.A(phase_increment_1__63__N_16[45]), .B(phase_increment_1__63__N_18[45]), 
         .C(rx_byte[0]), .Z(n2259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1122_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3708_add_4_16 (.A0(amdemod_out_d_11__N_2369[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2369[11]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16810), .S1(n36_adj_5841));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3708_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_3708_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3708_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3708_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3708_add_4_14 (.A0(amdemod_out_d_11__N_2369[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2369[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16809), .COUT(n16810), 
          .S0(n45_adj_5843), .S1(n42_adj_5842));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3708_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_3708_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_3708_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3708_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3708_add_4_12 (.A0(amdemod_out_d_11__N_2369[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2369[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16808), .COUT(n16809), 
          .S0(n51_adj_5845), .S1(n48_adj_5844));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3708_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_3708_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_3708_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3708_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3708_add_4_10 (.A0(amdemod_out_d_11__N_2369[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2369[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16807), .COUT(n16808), 
          .S0(n57_adj_5847), .S1(n54_adj_5846));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3708_add_4_10.INIT0 = 16'h555f;
    defparam _add_1_3708_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_3708_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3708_add_4_10.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_25__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[25]), .Z(n19479)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_25__bdd_2_lut_2_lut.init = 16'h4444;
    CCU2C _add_1_3708_add_4_8 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2369[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2369[4]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16806), .COUT(n16807), 
          .S0(n63_adj_5849), .S1(n60_adj_5848));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3708_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3708_add_4_8.INIT1 = 16'h555f;
    defparam _add_1_3708_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3708_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3708_add_4_6 (.A0(amdemod_out_d_11__N_2369[1]), .B0(square_sum[25]), 
          .C0(n30_adj_6282), .D0(n13890), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2369[2]), .D1(VCC_net), .CIN(n16805), 
          .COUT(n16806), .S0(n69_adj_5851), .S1(n66_adj_5850));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3708_add_4_6.INIT0 = 16'h596a;
    defparam _add_1_3708_add_4_6.INIT1 = 16'he1e1;
    defparam _add_1_3708_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3708_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3708_add_4_4 (.A0(n19816), .B0(square_sum[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_out_d_11__N_2369[0]), .B1(amdemod_out_d_11__N_2370[11]), 
          .C1(amdemod_out_d_11__N_2363), .D1(amdemod_out_d_11__N_2369[11]), 
          .CIN(n16804), .COUT(n16805), .S0(n75_adj_5853), .S1(n72_adj_5852));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3708_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3708_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_3708_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3708_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3708_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[16]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16804), .S1(n78_adj_5854));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3708_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3708_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3708_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3708_add_4_2.INJECT1_1 = "NO";
    Mixer mixer_inst (.mix_sinewave({mix_sinewave}), .clk_80mhz(clk_80mhz), 
          .mix_cosinewave({mix_cosinewave}), .diff_out_c(diff_out_c), .rf_in_c(rf_in_c), 
          .\lo_sinewave[0] (lo_sinewave[0]), .n67({n28_adj_6350, n31_adj_6351, 
          n34_adj_6352, n37_adj_6353, n40_adj_6354, n43_adj_6355, n46_adj_6356, 
          n49_adj_6357, n52_adj_6358, n55_adj_6359, n58_adj_6360, n61_adj_6361}), 
          .\lo_sinewave[8] (lo_sinewave[8]), .\lo_cosinewave[0] (lo_cosinewave[0]), 
          .n67_adj_451({n28_adj_6362, n31_adj_6363, n34_adj_6364, n37_adj_6365, 
          n40_adj_6366, n43_adj_6367, n46_adj_6368, n49_adj_6369, n52_adj_6370, 
          n55_adj_6371, n58_adj_6372, n61_adj_6373}), .\lo_sinewave[9] (lo_sinewave[9]), 
          .\lo_sinewave[12] (lo_sinewave[12]), .\lo_sinewave[10] (lo_sinewave[10]), 
          .\lo_sinewave[6] (lo_sinewave[6]), .\lo_sinewave[3] (lo_sinewave[3]), 
          .\lo_cosinewave[12] (lo_cosinewave[12]), .\lo_cosinewave[10] (lo_cosinewave[10]), 
          .\lo_cosinewave[9] (lo_cosinewave[9]), .\lo_cosinewave[8] (lo_cosinewave[8]), 
          .\lo_cosinewave[7] (lo_cosinewave[7]), .\lo_cosinewave[6] (lo_cosinewave[6]), 
          .\lo_cosinewave[5] (lo_cosinewave[5]), .\lo_cosinewave[4] (lo_cosinewave[4]), 
          .\lo_cosinewave[3] (lo_cosinewave[3]), .\lo_cosinewave[2] (lo_cosinewave[2]), 
          .\lo_cosinewave[1] (lo_cosinewave[1]), .\lo_sinewave[1] (lo_sinewave[1]), 
          .\lo_sinewave[2] (lo_sinewave[2]), .\lo_sinewave[4] (lo_sinewave[4]), 
          .\lo_sinewave[5] (lo_sinewave[5]), .\lo_sinewave[7] (lo_sinewave[7])) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(172[6] 180[5])
    CCU2C _add_1_3642_add_4_33 (.A0(comb_d9[67]), .B0(comb9[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[68]), .B1(comb9[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17268), .COUT(n17269), .S0(n88_adj_6531), 
          .S1(n85_adj_6530));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_33.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_33.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_33.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i1 (.D(n19579), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(phase_increment_1__63__N_21[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i1.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i115 (.D(\phase_increment[0] [50]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [50]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i115.GSR = "ENABLED";
    LUT4 phase_increment_1__63__N_21_53__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[53]), .Z(n19492)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_53__bdd_2_lut_2_lut.init = 16'h4444;
    CCU2C _add_1_3711_add_4_38 (.A0(comb_d8[71]), .B0(comb8[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16803), .S0(n78_adj_5855));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3711_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_38.INJECT1_1 = "NO";
    FD1S3AX phase_increment_0__i114 (.D(\phase_increment[0] [49]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i114.GSR = "ENABLED";
    LUT4 phase_increment_1__63__N_21_51__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[51]), .Z(n19508)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_51__bdd_2_lut_2_lut.init = 16'h4444;
    CCU2C _add_1_3711_add_4_36 (.A0(comb_d8[69]), .B0(comb8[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[70]), .B1(comb8[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16802), .COUT(n16803), .S0(n84_adj_5857), 
          .S1(n81_adj_5856));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_36.INJECT1_1 = "NO";
    FD1S3AX phase_increment_0__i113 (.D(\phase_increment[0] [48]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [48]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i113.GSR = "ENABLED";
    CCU2C _add_1_3642_add_4_31 (.A0(comb_d9[65]), .B0(comb9[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[66]), .B1(comb9[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17267), .COUT(n17268), .S0(n94_adj_6533), 
          .S1(n91_adj_6532));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_31.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_31.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_31.INJECT1_1 = "NO";
    FD1S3AX phase_increment_0__i112 (.D(\phase_increment[0] [47]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i112.GSR = "ENABLED";
    CCU2C _add_1_3711_add_4_34 (.A0(comb_d8[67]), .B0(comb8[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[68]), .B1(comb8[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16801), .COUT(n16802), .S0(n90_adj_5859), 
          .S1(n87_adj_5858));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_34.INJECT1_1 = "NO";
    FD1S3AX phase_increment_0__i111 (.D(\phase_increment[0] [46]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [46]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i111.GSR = "ENABLED";
    LUT4 mux_2067_i1_3_lut (.A(phase_increment_1__63__N_16[18]), .B(phase_increment_1__63__N_18[18]), 
         .C(rx_byte[0]), .Z(n3528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2067_i1_3_lut.init = 16'hcaca;
    FD1S3AX phase_increment_0__i110 (.D(\phase_increment[0] [45]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i110.GSR = "ENABLED";
    CCU2C _add_1_3711_add_4_32 (.A0(comb_d8[65]), .B0(comb8[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[66]), .B1(comb8[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16800), .COUT(n16801), .S0(n96_adj_5861), 
          .S1(n93_adj_5860));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_30 (.A0(comb_d8[63]), .B0(comb8[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[64]), .B1(comb8[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16799), .COUT(n16800), .S0(n102_adj_5863), 
          .S1(n99_adj_5862));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_28 (.A0(comb_d8[61]), .B0(comb8[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[62]), .B1(comb8[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16798), .COUT(n16799), .S0(n108_adj_5865), 
          .S1(n105_adj_5864));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_28.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i39 (.D(n204), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i39.GSR = "ENABLED";
    CCU2C _add_1_3711_add_4_26 (.A0(comb_d8[59]), .B0(comb8[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[60]), .B1(comb8[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16797), .COUT(n16798), .S0(n114_adj_5867), 
          .S1(n111_adj_5866));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_24 (.A0(comb_d8[57]), .B0(comb8[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[58]), .B1(comb8[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16796), .COUT(n16797), .S0(n120_adj_5869), 
          .S1(n117_adj_5868));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_22 (.A0(comb_d8[55]), .B0(comb8[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[56]), .B1(comb8[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16795), .COUT(n16796), .S0(n126_adj_5871), 
          .S1(n123_adj_5870));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_20 (.A0(comb_d8[53]), .B0(comb8[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[54]), .B1(comb8[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16794), .COUT(n16795), .S0(n132_adj_5873), 
          .S1(n129_adj_5872));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_18 (.A0(comb_d8[51]), .B0(comb8[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[52]), .B1(comb8[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16793), .COUT(n16794), .S0(n138_adj_5875), 
          .S1(n135_adj_5874));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_16 (.A0(comb_d8[49]), .B0(comb8[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[50]), .B1(comb8[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16792), .COUT(n16793), .S0(n144_adj_5877), 
          .S1(n141_adj_5876));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_14 (.A0(comb_d8[47]), .B0(comb8[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[48]), .B1(comb8[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16791), .COUT(n16792), .S0(n150_adj_5879), 
          .S1(n147_adj_5878));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_12 (.A0(comb_d8[45]), .B0(comb8[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[46]), .B1(comb8[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16790), .COUT(n16791), .S0(n156_adj_5881), 
          .S1(n153_adj_5880));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_10 (.A0(comb_d8[43]), .B0(comb8[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[44]), .B1(comb8[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16789), .COUT(n16790), .S0(n162_adj_5883), 
          .S1(n159_adj_5882));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_8 (.A0(comb_d8[41]), .B0(comb8[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[42]), .B1(comb8[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16788), .COUT(n16789), .S0(n168_adj_5885), 
          .S1(n165_adj_5884));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_6 (.A0(comb_d8[39]), .B0(comb8[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[40]), .B1(comb8[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16787), .COUT(n16788), .S0(n174_adj_5887), 
          .S1(n171_adj_5886));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_4 (.A0(comb_d8[37]), .B0(comb8[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[38]), .B1(comb8[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16786), .COUT(n16787), .S0(n180_adj_5889), 
          .S1(n177_adj_5888));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3711_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3711_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[36]), .B1(comb8[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16786), .S1(n183_adj_5890));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3711_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3711_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3711_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3711_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_38 (.A0(comb_d8_adj_6568[35]), .B0(comb8_adj_6567[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16785), .S0(comb9_71__N_2209_adj_6592[35]), 
          .S1(cout_adj_5891));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3714_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_36 (.A0(comb_d8_adj_6568[33]), .B0(comb8_adj_6567[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[34]), .B1(comb8_adj_6567[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16784), .COUT(n16785), .S0(comb9_71__N_2209_adj_6592[33]), 
          .S1(comb9_71__N_2209_adj_6592[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_34 (.A0(comb_d8_adj_6568[31]), .B0(comb8_adj_6567[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[32]), .B1(comb8_adj_6567[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16783), .COUT(n16784), .S0(comb9_71__N_2209_adj_6592[31]), 
          .S1(comb9_71__N_2209_adj_6592[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_32 (.A0(comb_d8_adj_6568[29]), .B0(comb8_adj_6567[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[30]), .B1(comb8_adj_6567[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16782), .COUT(n16783), .S0(comb9_71__N_2209_adj_6592[29]), 
          .S1(comb9_71__N_2209_adj_6592[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_30 (.A0(comb_d8_adj_6568[27]), .B0(comb8_adj_6567[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[28]), .B1(comb8_adj_6567[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16781), .COUT(n16782), .S0(comb9_71__N_2209_adj_6592[27]), 
          .S1(comb9_71__N_2209_adj_6592[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_28 (.A0(comb_d8_adj_6568[25]), .B0(comb8_adj_6567[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[26]), .B1(comb8_adj_6567[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16780), .COUT(n16781), .S0(comb9_71__N_2209_adj_6592[25]), 
          .S1(comb9_71__N_2209_adj_6592[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_26 (.A0(comb_d8_adj_6568[23]), .B0(comb8_adj_6567[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[24]), .B1(comb8_adj_6567[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16779), .COUT(n16780), .S0(comb9_71__N_2209_adj_6592[23]), 
          .S1(comb9_71__N_2209_adj_6592[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_24 (.A0(comb_d8_adj_6568[21]), .B0(comb8_adj_6567[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[22]), .B1(comb8_adj_6567[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16778), .COUT(n16779), .S0(comb9_71__N_2209_adj_6592[21]), 
          .S1(comb9_71__N_2209_adj_6592[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_24.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i38 (.D(n207), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[38]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i38.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i109 (.D(\phase_increment[0] [44]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [44]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i109.GSR = "ENABLED";
    CCU2C _add_1_3714_add_4_22 (.A0(comb_d8_adj_6568[19]), .B0(comb8_adj_6567[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[20]), .B1(comb8_adj_6567[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16777), .COUT(n16778), .S0(comb9_71__N_2209_adj_6592[19]), 
          .S1(comb9_71__N_2209_adj_6592[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_20 (.A0(comb_d8_adj_6568[17]), .B0(comb8_adj_6567[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[18]), .B1(comb8_adj_6567[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16776), .COUT(n16777), .S0(comb9_71__N_2209_adj_6592[17]), 
          .S1(comb9_71__N_2209_adj_6592[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_20.INJECT1_1 = "NO";
    LUT4 mux_1799_i1_3_lut (.A(phase_increment_1__63__N_19[26]), .B(phase_increment_1__63__N_20[26]), 
         .C(rx_byte[0]), .Z(n3167)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1799_i1_3_lut.init = 16'hcaca;
    FD1S3AX phase_increment_0__i108 (.D(\phase_increment[0] [43]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i108.GSR = "ENABLED";
    CCU2C _add_1_3792_add_4_34 (.A0(mix_sinewave[11]), .B0(integrator1[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17754), .COUT(n17755), .S0(n90_adj_6205), 
          .S1(n87_adj_6204));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_34.INJECT1_1 = "NO";
    FD1S3AX phase_increment_0__i107 (.D(\phase_increment[0] [42]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [42]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i107.GSR = "ENABLED";
    CCU2C _add_1_3714_add_4_18 (.A0(comb_d8_adj_6568[15]), .B0(comb8_adj_6567[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[16]), .B1(comb8_adj_6567[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16775), .COUT(n16776), .S0(comb9_71__N_2209_adj_6592[15]), 
          .S1(comb9_71__N_2209_adj_6592[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3642_add_4_29 (.A0(comb_d9[63]), .B0(comb9[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[64]), .B1(comb9[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17266), .COUT(n17267), .S0(n100_adj_6535), 
          .S1(n97_adj_6534));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_29.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_29.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_16 (.A0(comb_d8_adj_6568[13]), .B0(comb8_adj_6567[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[14]), .B1(comb8_adj_6567[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16774), .COUT(n16775), .S0(comb9_71__N_2209_adj_6592[13]), 
          .S1(comb9_71__N_2209_adj_6592[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_14 (.A0(comb_d8_adj_6568[11]), .B0(comb8_adj_6567[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[12]), .B1(comb8_adj_6567[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16773), .COUT(n16774), .S0(comb9_71__N_2209_adj_6592[11]), 
          .S1(comb9_71__N_2209_adj_6592[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_12 (.A0(comb_d8_adj_6568[9]), .B0(comb8_adj_6567[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[10]), .B1(comb8_adj_6567[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16772), .COUT(n16773), .S0(comb9_71__N_2209_adj_6592[9]), 
          .S1(comb9_71__N_2209_adj_6592[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_10 (.A0(comb_d8_adj_6568[7]), .B0(comb8_adj_6567[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[8]), .B1(comb8_adj_6567[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16771), .COUT(n16772), .S0(comb9_71__N_2209_adj_6592[7]), 
          .S1(comb9_71__N_2209_adj_6592[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_8 (.A0(comb_d8_adj_6568[5]), .B0(comb8_adj_6567[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[6]), .B1(comb8_adj_6567[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16770), .COUT(n16771), .S0(comb9_71__N_2209_adj_6592[5]), 
          .S1(comb9_71__N_2209_adj_6592[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_6 (.A0(comb_d8_adj_6568[3]), .B0(comb8_adj_6567[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[4]), .B1(comb8_adj_6567[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16769), .COUT(n16770), .S0(comb9_71__N_2209_adj_6592[3]), 
          .S1(comb9_71__N_2209_adj_6592[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3714_add_4_4 (.A0(comb_d8_adj_6568[1]), .B0(comb8_adj_6567[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[2]), .B1(comb8_adj_6567[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16768), .COUT(n16769), .S0(comb9_71__N_2209_adj_6592[1]), 
          .S1(comb9_71__N_2209_adj_6592[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3714_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3642_add_4_27 (.A0(comb_d9[61]), .B0(comb9[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[62]), .B1(comb9[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17265), .COUT(n17266), .S0(n106_adj_6537), 
          .S1(n103_adj_6536));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_27.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_27.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_27.INJECT1_1 = "NO";
    LUT4 mux_1717_i1_3_lut (.A(phase_increment_1__63__N_16[28]), .B(phase_increment_1__63__N_18[28]), 
         .C(rx_byte[0]), .Z(n3058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1717_i1_3_lut.init = 16'hcaca;
    FD1S3AX phase_accumulator_e3_i0_i37 (.D(n210), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i37.GSR = "ENABLED";
    CCU2C _add_1_3714_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8_adj_6568[0]), .B1(comb8_adj_6567[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16768), .S1(comb9_71__N_2209_adj_6592[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3714_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3714_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3714_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3714_add_4_2.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i36 (.D(n213), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[36]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i36.GSR = "ENABLED";
    CCU2C phase_accumulator_add_4_64 (.A0(\phase_increment[1] [62]), .B0(phase_accumulator_adj_6545[62]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [63]), .B1(phase_accumulator_adj_6545[63]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16766), .S0(n135_adj_5287), 
          .S1(n132_adj_5305));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_64.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_64.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_64.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_64.INJECT1_1 = "NO";
    PFUMX mux_1638_i1 (.BLUT(n2942), .ALUT(n2948), .C0(n19297), .Z(n2951));
    PFUMX mux_726_i1 (.BLUT(n1710), .ALUT(n1720), .C0(led_0_6), .Z(n1726));
    CCU2C phase_accumulator_add_4_62 (.A0(\phase_increment[1] [60]), .B0(phase_accumulator_adj_6545[60]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [61]), .B1(phase_accumulator_adj_6545[61]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16765), .COUT(n16766), .S0(n141_adj_3522), 
          .S1(n138_adj_5292));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_62.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_62.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_62.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_62.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_10__bdd_2_lut_8995 (.A(phase_increment_1__63__N_21[10]), 
         .B(rx_byte[0]), .Z(n19542)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_10__bdd_2_lut_8995.init = 16'heeee;
    CCU2C phase_accumulator_add_4_60 (.A0(\phase_increment[1] [58]), .B0(phase_accumulator_adj_6545[58]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [59]), .B1(phase_accumulator_adj_6545[59]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16764), .COUT(n16765), .S0(n147_adj_5320), 
          .S1(n144_adj_5332));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_60.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_60.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_60.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_60.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i35 (.D(n216), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i35.GSR = "ENABLED";
    CCU2C _add_1_3792_add_4_32 (.A0(mix_sinewave[11]), .B0(integrator1[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17753), .COUT(n17754), .S0(n96_adj_6207), 
          .S1(n93_adj_6206));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3642_add_4_25 (.A0(comb_d9[59]), .B0(comb9[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[60]), .B1(comb9[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17264), .COUT(n17265), .S0(n112_adj_6539), 
          .S1(n109_adj_6538));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_25.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_25.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3642_add_4_23 (.A0(comb_d9[57]), .B0(comb9[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[58]), .B1(comb9[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17263), .COUT(n17264), .S0(n118_adj_6541), 
          .S1(n115_adj_6540));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_23.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_23.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_23.INJECT1_1 = "NO";
    CCU2C phase_accumulator_add_4_58 (.A0(\phase_increment[1] [56]), .B0(phase_accumulator_adj_6545[56]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [57]), .B1(phase_accumulator_adj_6545[57]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16763), .COUT(n16764), .S0(n153_adj_5302), 
          .S1(n150_adj_5329));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_58.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_58.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_58.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_58.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i34 (.D(n219), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i34.GSR = "ENABLED";
    CCU2C phase_accumulator_add_4_56 (.A0(\phase_increment[1] [54]), .B0(phase_accumulator_adj_6545[54]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [55]), .B1(phase_accumulator_adj_6545[55]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16762), .COUT(n16763), .S0(n159_adj_5321), 
          .S1(n156_adj_5297));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_56.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_56.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_56.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_56.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_18__bdd_2_lut_8650_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[18]), .Z(n19515)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_18__bdd_2_lut_8650_2_lut.init = 16'h4444;
    CCU2C phase_accumulator_add_4_54 (.A0(\phase_increment[1] [52]), .B0(phase_accumulator_adj_6545[52]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [53]), .B1(phase_accumulator_adj_6545[53]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16761), .COUT(n16762), .S0(n165_adj_5308), 
          .S1(n162_adj_5317));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_54.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_54.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_54.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_54.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i33 (.D(n222), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i33.GSR = "ENABLED";
    CCU2C phase_accumulator_add_4_52 (.A0(\phase_increment[1] [50]), .B0(phase_accumulator_adj_6545[50]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [51]), .B1(phase_accumulator_adj_6545[51]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16760), .COUT(n16761), .S0(n171_adj_5291), 
          .S1(n168_adj_5353));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_52.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_52.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_52.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_52.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_31 (.A0(\phase_increment[0] [30]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [31]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17613), .COUT(n17614), .S0(phase_increment_1__63__N_20[30]), 
          .S1(phase_increment_1__63__N_20[31]));
    defparam _add_1_3813_add_4_31.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_30 (.A0(mix_sinewave[11]), .B0(integrator1[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17752), .COUT(n17753), .S0(n102_adj_6209), 
          .S1(n99_adj_6208));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_28 (.A0(mix_sinewave[11]), .B0(integrator1[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17751), .COUT(n17752), .S0(n108_adj_6211), 
          .S1(n105_adj_6210));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3642_add_4_21 (.A0(comb_d9[55]), .B0(comb9[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[56]), .B1(comb9[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17262), .COUT(n17263));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_21.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_21.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_26 (.A0(mix_sinewave[11]), .B0(integrator1[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17750), .COUT(n17751), .S0(n114_adj_6213), 
          .S1(n111_adj_6212));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_24 (.A0(mix_sinewave[11]), .B0(integrator1[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17749), .COUT(n17750), .S0(n120_adj_6215), 
          .S1(n117_adj_6214));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_22 (.A0(mix_sinewave[11]), .B0(integrator1[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17748), .COUT(n17749), .S0(n126_adj_6217), 
          .S1(n123_adj_6216));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_22.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_48__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[48]), .Z(n19525)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_48__bdd_2_lut_2_lut.init = 16'h4444;
    CCU2C _add_1_3813_add_4_29 (.A0(\phase_increment[0] [28]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [29]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17612), .COUT(n17613), .S0(phase_increment_1__63__N_20[28]), 
          .S1(phase_increment_1__63__N_20[29]));
    defparam _add_1_3813_add_4_29.INIT0 = 16'haaa0;
    defparam _add_1_3813_add_4_29.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_29.INJECT1_1 = "NO";
    CCU2C phase_accumulator_add_4_50 (.A0(\phase_increment[1] [48]), .B0(phase_accumulator_adj_6545[48]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [49]), .B1(phase_accumulator_adj_6545[49]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16759), .COUT(n16760), .S0(n177_adj_5326), 
          .S1(n174_adj_5285));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_50.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_50.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_50.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_50.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i32 (.D(n225), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i32.GSR = "ENABLED";
    CCU2C phase_accumulator_add_4_48 (.A0(\phase_increment[1] [46]), .B0(phase_accumulator_adj_6545[46]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [47]), .B1(phase_accumulator_adj_6545[47]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16758), .COUT(n16759), .S0(n183_adj_5295), 
          .S1(n180_adj_5341));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_48.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_48.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_48.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_48.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_46__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[46]), .Z(n19551)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_46__bdd_2_lut_2_lut.init = 16'h4444;
    LUT4 i8043_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19762), 
         .D(n3966), .Z(n3982)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8043_3_lut_4_lut.init = 16'hf780;
    LUT4 phase_increment_1__63__N_21_33__bdd_2_lut_8654 (.A(phase_increment_1__63__N_17[33]), 
         .B(led_0_6), .Z(n19700)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_33__bdd_2_lut_8654.init = 16'heeee;
    LUT4 i8224_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19555), 
         .D(n2180), .Z(n2196)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8224_3_lut_4_lut.init = 16'hf780;
    CCU2C phase_accumulator_add_4_46 (.A0(\phase_increment[1] [44]), .B0(phase_accumulator_adj_6545[44]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [45]), .B1(phase_accumulator_adj_6545[45]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16757), .COUT(n16758), .S0(n189), 
          .S1(n186));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_46.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_46.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_46.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_46.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i31 (.D(n228), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i31.GSR = "ENABLED";
    CCU2C phase_accumulator_add_4_44 (.A0(\phase_increment[1] [42]), .B0(phase_accumulator_adj_6545[42]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [43]), .B1(phase_accumulator_adj_6545[43]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16756), .COUT(n16757), .S0(n195), 
          .S1(n192));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_44.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_44.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_44.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_44.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_20 (.A0(mix_sinewave[11]), .B0(integrator1[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17747), .COUT(n17748), .S0(n132_adj_6219), 
          .S1(n129_adj_6218));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_18 (.A0(mix_sinewave[11]), .B0(integrator1[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17746), .COUT(n17747), .S0(n138_adj_6221), 
          .S1(n135_adj_6220));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3642_add_4_19 (.A0(comb_d9[53]), .B0(comb9[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[54]), .B1(comb9[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17261), .COUT(n17262));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_19.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_19.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3642_add_4_17 (.A0(comb_d9[51]), .B0(comb9[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[52]), .B1(comb9[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17260), .COUT(n17261));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_17.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_17.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_16 (.A0(mix_sinewave[11]), .B0(integrator1[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17745), .COUT(n17746), .S0(n144_adj_6223), 
          .S1(n141_adj_6222));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_14 (.A0(mix_sinewave[11]), .B0(integrator1[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17744), .COUT(n17745), .S0(n150_adj_6225), 
          .S1(n147_adj_6224));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_27 (.A0(\phase_increment[0] [26]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [27]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17611), .COUT(n17612), .S0(phase_increment_1__63__N_20[26]), 
          .S1(phase_increment_1__63__N_20[27]));
    defparam _add_1_3813_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_25 (.A0(\phase_increment[0] [24]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [25]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17610), .COUT(n17611), .S0(phase_increment_1__63__N_20[24]), 
          .S1(phase_increment_1__63__N_20[25]));
    defparam _add_1_3813_add_4_25.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_25.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_23 (.A0(\phase_increment[0] [22]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [23]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17609), .COUT(n17610), .S0(phase_increment_1__63__N_20[22]), 
          .S1(phase_increment_1__63__N_20[23]));
    defparam _add_1_3813_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_21 (.A0(\phase_increment[0] [20]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [21]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17608), .COUT(n17609), .S0(phase_increment_1__63__N_20[20]), 
          .S1(phase_increment_1__63__N_20[21]));
    defparam _add_1_3813_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_19 (.A0(\phase_increment[0] [18]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [19]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17607), .COUT(n17608), .S0(phase_increment_1__63__N_20[18]), 
          .S1(phase_increment_1__63__N_20[19]));
    defparam _add_1_3813_add_4_19.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_17 (.A0(\phase_increment[0] [16]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [17]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17606), .COUT(n17607), .S0(phase_increment_1__63__N_20[16]), 
          .S1(phase_increment_1__63__N_20[17]));
    defparam _add_1_3813_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_3813_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_17.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_33__bdd_2_lut_8973 (.A(phase_increment_1__63__N_21[33]), 
         .B(rx_byte[0]), .Z(n19701)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_33__bdd_2_lut_8973.init = 16'heeee;
    CCU2C phase_accumulator_add_4_42 (.A0(\phase_increment[1] [40]), .B0(phase_accumulator_adj_6545[40]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [41]), .B1(phase_accumulator_adj_6545[41]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16755), .COUT(n16756), .S0(n201), 
          .S1(n198));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_42.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_42.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_42.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_42.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i30 (.D(n231), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i30.GSR = "ENABLED";
    CCU2C phase_accumulator_add_4_40 (.A0(\phase_increment[1] [38]), .B0(phase_accumulator_adj_6545[38]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [39]), .B1(phase_accumulator_adj_6545[39]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16754), .COUT(n16755), .S0(n207), 
          .S1(n204));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_40.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_40.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_40.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_40.INJECT1_1 = "NO";
    PFUMX mux_584_i1 (.BLUT(n1527), .ALUT(n1512), .C0(rx_byte[2]), .Z(n1535));
    LUT4 mux_1227_i1_3_lut (.A(phase_increment_1__63__N_16[42]), .B(phase_increment_1__63__N_18[42]), 
         .C(rx_byte[0]), .Z(n2400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1227_i1_3_lut.init = 16'hcaca;
    LUT4 phase_increment_1__63__N_21_0__bdd_4_lut_3_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_19[0]), 
         .C(phase_increment_1__63__N_21[0]), .Z(n19577)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_0__bdd_4_lut_3_lut.init = 16'he4e4;
    CCU2C phase_accumulator_add_4_38 (.A0(\phase_increment[1] [36]), .B0(phase_accumulator_adj_6545[36]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [37]), .B1(phase_accumulator_adj_6545[37]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16753), .COUT(n16754), .S0(n213), 
          .S1(n210));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_38.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_38.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_38.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_38.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i29 (.D(n234), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i29.GSR = "ENABLED";
    CCU2C phase_accumulator_add_4_36 (.A0(\phase_increment[1] [34]), .B0(phase_accumulator_adj_6545[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [35]), .B1(phase_accumulator_adj_6545[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16752), .COUT(n16753), .S0(n219), 
          .S1(n216));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_36.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_36.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_36.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_15 (.A0(\phase_increment[0] [14]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [15]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17605), .COUT(n17606), .S0(phase_increment_1__63__N_20[14]), 
          .S1(phase_increment_1__63__N_20[15]));
    defparam _add_1_3813_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_13 (.A0(\phase_increment[0] [12]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [13]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17604), .COUT(n17605), .S0(phase_increment_1__63__N_20[12]), 
          .S1(phase_increment_1__63__N_20[13]));
    defparam _add_1_3813_add_4_13.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_11 (.A0(\phase_increment[0] [10]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [11]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17603), .COUT(n17604), .S0(phase_increment_1__63__N_20[10]), 
          .S1(phase_increment_1__63__N_20[11]));
    defparam _add_1_3813_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3813_add_4_11.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_12 (.A0(mix_sinewave[11]), .B0(integrator1[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17743), .COUT(n17744), .S0(n156_adj_6227), 
          .S1(n153_adj_6226));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_10 (.A0(mix_sinewave[11]), .B0(integrator1[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17742), .COUT(n17743), .S0(n162_adj_6229), 
          .S1(n159_adj_6228));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_8 (.A0(mix_sinewave[11]), .B0(integrator1[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17741), .COUT(n17742), .S0(n168_adj_6231), 
          .S1(n165_adj_6230));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_6 (.A0(mix_sinewave[11]), .B0(integrator1[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17740), .COUT(n17741), .S0(n174_adj_6233), 
          .S1(n171_adj_6232));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_4 (.A0(mix_sinewave[11]), .B0(integrator1[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17739), .COUT(n17740), .S0(n180_adj_6235), 
          .S1(n177_adj_6234));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3792_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3792_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17739), .S1(n183_adj_6236));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3792_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3792_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3792_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3792_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3795_add_4_10 (.A0(square_sum[25]), .B0(n19824), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17737), .S0(n27_adj_6238), .S1(n24_adj_6237));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3795_add_4_10.INIT0 = 16'heee1;
    defparam _add_1_3795_add_4_10.INIT1 = 16'heee1;
    defparam _add_1_3795_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3795_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3642_add_4_15 (.A0(comb_d9[49]), .B0(comb9[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[50]), .B1(comb9[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17259), .COUT(n17260));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_15.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_15.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_15.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_42__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[42]), .Z(n19602)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_42__bdd_2_lut_2_lut.init = 16'h4444;
    CCU2C phase_accumulator_add_4_34 (.A0(\phase_increment[1] [32]), .B0(phase_accumulator_adj_6545[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [33]), .B1(phase_accumulator_adj_6545[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16751), .COUT(n16752), .S0(n225), 
          .S1(n222));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_34.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_34.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_34.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_34.INJECT1_1 = "NO";
    CCU2C phase_accumulator_add_4_32 (.A0(\phase_increment[1] [30]), .B0(phase_accumulator_adj_6545[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [31]), .B1(phase_accumulator_adj_6545[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16750), .COUT(n16751), .S0(n231), 
          .S1(n228));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_32.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_32.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_32.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_9 (.A0(\phase_increment[0] [8]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [9]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17602), .COUT(n17603), .S0(phase_increment_1__63__N_20[8]), 
          .S1(phase_increment_1__63__N_20[9]));
    defparam _add_1_3813_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_3813_add_4_9.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3642_add_4_13 (.A0(comb_d9[47]), .B0(comb9[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[48]), .B1(comb9[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17258), .COUT(n17259));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_13.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_13.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_13.INJECT1_1 = "NO";
    CCU2C phase_accumulator_add_4_30 (.A0(\phase_increment[1] [28]), .B0(phase_accumulator_adj_6545[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [29]), .B1(phase_accumulator_adj_6545[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16749), .COUT(n16750), .S0(n237), 
          .S1(n234));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_30.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_30.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_30.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_30.INJECT1_1 = "NO";
    CCU2C phase_accumulator_add_4_28 (.A0(\phase_increment[1] [26]), .B0(phase_accumulator_adj_6545[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [27]), .B1(phase_accumulator_adj_6545[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16748), .COUT(n16749), .S0(n243), 
          .S1(n240));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_28.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_28.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_28.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_28.INJECT1_1 = "NO";
    FD1S3AX phase_increment_0__i106 (.D(\phase_increment[0] [41]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i106.GSR = "ENABLED";
    CCU2C phase_accumulator_add_4_26 (.A0(\phase_increment[1] [24]), .B0(phase_accumulator_adj_6545[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [25]), .B1(phase_accumulator_adj_6545[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16747), .COUT(n16748), .S0(n249), 
          .S1(n246));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_26.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_26.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_26.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_26.INJECT1_1 = "NO";
    LUT4 i8111_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19480), 
         .D(n3214), .Z(n3230)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8111_3_lut_4_lut.init = 16'hf780;
    CCU2C phase_accumulator_add_4_24 (.A0(\phase_increment[1] [22]), .B0(phase_accumulator_adj_6545[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [23]), .B1(phase_accumulator_adj_6545[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16746), .COUT(n16747), .S0(n255), 
          .S1(n252));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_24.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_24.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_24.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_24.INJECT1_1 = "NO";
    LUT4 mux_1842_i1_3_lut (.A(rx_byte[2]), .B(n3199), .C(rx_byte[3]), 
         .Z(n3224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1842_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3813_add_4_7 (.A0(\phase_increment[0] [6]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [7]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17601), .COUT(n17602), .S0(phase_increment_1__63__N_20[6]), 
          .S1(phase_increment_1__63__N_20[7]));
    defparam _add_1_3813_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_3813_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_5 (.A0(\phase_increment[0] [4]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [5]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17600), .COUT(n17601), .S0(phase_increment_1__63__N_20[4]), 
          .S1(phase_increment_1__63__N_20[5]));
    defparam _add_1_3813_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_3813_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_3 (.A0(phase_increment_1__63__N_17[2]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_increment_1__63__N_17[3]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17599), .COUT(n17600), 
          .S0(phase_increment_1__63__N_20[2]), .S1(phase_increment_1__63__N_20[3]));
    defparam _add_1_3813_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_3813_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_increment_1__63__N_17[1]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .COUT(n17599), .S1(phase_increment_1__63__N_20[1]));
    defparam _add_1_3813_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3813_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17598), .S0(cout_adj_6289));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_36 (.A0(mix_sinewave[11]), .B0(integrator1[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17597), .COUT(n17598), .S0(integrator1_71__N_960[34]), 
          .S1(integrator1_71__N_960[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_34 (.A0(mix_sinewave[11]), .B0(integrator1[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17596), .COUT(n17597), .S0(integrator1_71__N_960[32]), 
          .S1(integrator1_71__N_960[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_32 (.A0(mix_sinewave[11]), .B0(integrator1[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17595), .COUT(n17596), .S0(integrator1_71__N_960[30]), 
          .S1(integrator1_71__N_960[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_add_4_32.INJECT1_1 = "NO";
    CCU2C phase_accumulator_add_4_22 (.A0(\phase_increment[1] [20]), .B0(phase_accumulator_adj_6545[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [21]), .B1(phase_accumulator_adj_6545[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16745), .COUT(n16746), .S0(n261), 
          .S1(n258));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_22.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_22.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_22.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3795_add_4_8 (.A0(n19828), .B0(n19827), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17736), .COUT(n17737), .S0(n33_adj_6240), 
          .S1(n30_adj_6239));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3795_add_4_8.INIT0 = 16'heee1;
    defparam _add_1_3795_add_4_8.INIT1 = 16'h6669;
    defparam _add_1_3795_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3795_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3795_add_4_6 (.A0(square_sum[25]), .B0(n4_adj_6510), .C0(amdemod_out_d_11__N_2358[5]), 
          .D0(VCC_net), .A1(n19828), .B1(n19827), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17735), .COUT(n17736), .S0(n39), .S1(n36_adj_6241));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3795_add_4_6.INIT0 = 16'h6969;
    defparam _add_1_3795_add_4_6.INIT1 = 16'heee1;
    defparam _add_1_3795_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3795_add_4_6.INJECT1_1 = "NO";
    LUT4 mux_1192_i1_3_lut (.A(phase_increment_1__63__N_16[43]), .B(phase_increment_1__63__N_18[43]), 
         .C(rx_byte[0]), .Z(n2353)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1192_i1_3_lut.init = 16'hcaca;
    CCU2C phase_accumulator_add_4_20 (.A0(\phase_increment[1] [18]), .B0(phase_accumulator_adj_6545[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [19]), .B1(phase_accumulator_adj_6545[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16744), .COUT(n16745), .S0(n267), 
          .S1(n264));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_20.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_20.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_20.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_30 (.A0(mix_sinewave[11]), .B0(integrator1[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17594), .COUT(n17595), .S0(integrator1_71__N_960[28]), 
          .S1(integrator1_71__N_960[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_add_4_30.INJECT1_1 = "NO";
    CCU2C phase_accumulator_add_4_18 (.A0(\phase_increment[1] [16]), .B0(phase_accumulator_adj_6545[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [17]), .B1(phase_accumulator_adj_6545[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16743), .COUT(n16744), .S0(n273), 
          .S1(n270));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_18.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_18.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_18.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_18.INJECT1_1 = "NO";
    CCU2C phase_accumulator_add_4_16 (.A0(\phase_increment[1] [14]), .B0(phase_accumulator_adj_6545[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [15]), .B1(phase_accumulator_adj_6545[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16742), .COUT(n16743), .S0(n279), 
          .S1(n276));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_16.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_16.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_16.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_16.INJECT1_1 = "NO";
    CCU2C phase_accumulator_add_4_14 (.A0(\phase_increment[1] [12]), .B0(phase_accumulator_adj_6545[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [13]), .B1(phase_accumulator_adj_6545[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16741), .COUT(n16742), .S0(n285), 
          .S1(n282));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_14.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_14.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_14.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_28 (.A0(mix_sinewave[11]), .B0(integrator1[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17593), .COUT(n17594), .S0(integrator1_71__N_960[26]), 
          .S1(integrator1_71__N_960[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_add_4_28.INJECT1_1 = "NO";
    CCU2C phase_accumulator_add_4_12 (.A0(\phase_increment[1] [10]), .B0(phase_accumulator_adj_6545[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [11]), .B1(phase_accumulator_adj_6545[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16740), .COUT(n16741), .S0(n291), 
          .S1(n288));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_12.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_12.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_12.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3795_add_4_4 (.A0(square_sum[25]), .B0(n19824), .C0(square_sum[21]), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), .C1(square_sum[22]), 
          .D1(VCC_net), .CIN(n17734), .COUT(n17735), .S0(n45_adj_6243), 
          .S1(n42_adj_6242));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3795_add_4_4.INIT0 = 16'h1e1e;
    defparam _add_1_3795_add_4_4.INIT1 = 16'h1e11;
    defparam _add_1_3795_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3795_add_4_4.INJECT1_1 = "NO";
    OB pwm_out_pad (.I(pwm_out_c), .O(pwm_out));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(42[22:29])
    CCU2C phase_accumulator_add_4_10 (.A0(\phase_increment[1] [8]), .B0(phase_accumulator_adj_6545[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [9]), .B1(phase_accumulator_adj_6545[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16739), .COUT(n16740), .S0(n297), 
          .S1(n294));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_10.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_10.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_10.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_26 (.A0(mix_sinewave[11]), .B0(integrator1[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17592), .COUT(n17593), .S0(integrator1_71__N_960[24]), 
          .S1(integrator1_71__N_960[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_add_4_26.INJECT1_1 = "NO";
    CCU2C phase_accumulator_add_4_8 (.A0(\phase_increment[1] [6]), .B0(phase_accumulator_adj_6545[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [7]), .B1(phase_accumulator_adj_6545[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16738), .COUT(n16739), .S0(n303), 
          .S1(n300));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_8.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_8.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_8.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_8.INJECT1_1 = "NO";
    L6MUX21 i8445 (.D0(n19424), .D1(n19421), .SD(n19822), .Z(n19425));
    CCU2C phase_accumulator_add_4_6 (.A0(\phase_increment[1] [4]), .B0(phase_accumulator_adj_6545[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [5]), .B1(phase_accumulator_adj_6545[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16737), .COUT(n16738), .S0(n309), 
          .S1(n306));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_6.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_6.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_6.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_6.INJECT1_1 = "NO";
    CCU2C phase_accumulator_add_4_4 (.A0(\phase_increment[1] [2]), .B0(phase_accumulator_adj_6545[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [3]), .B1(phase_accumulator_adj_6545[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16736), .COUT(n16737), .S0(n315), 
          .S1(n312));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_4.INIT0 = 16'h666a;
    defparam phase_accumulator_add_4_4.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_4.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_4.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i60 (.D(n141_adj_3522), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[60]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i60.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i59 (.D(n144_adj_5332), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i59.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i58 (.D(n147_adj_5320), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[58]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i58.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i57 (.D(n150_adj_5329), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i57.GSR = "ENABLED";
    CCU2C _add_1_3621_add_4_20 (.A0(comb_d9[17]), .B0(comb9[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[18]), .B1(comb9[18]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17393), .COUT(n17394));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3621_add_4_22 (.A0(comb_d9[19]), .B0(comb9[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[20]), .B1(comb9[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17394), .COUT(n17395));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_22.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i56 (.D(n153_adj_5302), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[56]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i56.GSR = "ENABLED";
    CCU2C _add_1_add_4_24 (.A0(mix_sinewave[11]), .B0(integrator1[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17591), .COUT(n17592), .S0(integrator1_71__N_960[22]), 
          .S1(integrator1_71__N_960[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_add_4_24.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i55 (.D(n156_adj_5297), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i55.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i54 (.D(n159_adj_5321), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[54]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i54.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i53 (.D(n162_adj_5317), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i53.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i52 (.D(n165_adj_5308), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[52]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i52.GSR = "ENABLED";
    CCU2C _add_1_3642_add_4_11 (.A0(comb_d9[45]), .B0(comb9[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[46]), .B1(comb9[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17257), .COUT(n17258));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3642_add_4_9 (.A0(comb_d9[43]), .B0(comb9[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[44]), .B1(comb9[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17256), .COUT(n17257));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_9.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i51 (.D(n168_adj_5353), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i51.GSR = "ENABLED";
    LUT4 i8234_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19526), 
         .D(n2133), .Z(n2149)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8234_3_lut_4_lut.init = 16'hf780;
    CCU2C _add_1_3621_add_4_18 (.A0(comb_d9[15]), .B0(comb9[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[16]), .B1(comb9[16]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17392), .COUT(n17393));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3795_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[20]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17734), .S1(n48_adj_6244));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3795_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3795_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3795_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3795_add_4_2.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_43__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[43]), .Z(n19605)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_43__bdd_2_lut_2_lut.init = 16'h4444;
    CCU2C _add_1_3621_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[0]), .B1(comb9[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17385));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3621_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_2.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i50 (.D(n171_adj_5291), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[50]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i50.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i49 (.D(n174_adj_5285), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i49.GSR = "ENABLED";
    CCU2C phase_accumulator_add_4_2 (.A0(\phase_increment[1] [0]), .B0(phase_accumulator_adj_6545[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[1] [1]), .B1(phase_accumulator_adj_6545[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16736), .S1(n318));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_add_4_2.INIT0 = 16'h0008;
    defparam phase_accumulator_add_4_2.INIT1 = 16'h666a;
    defparam phase_accumulator_add_4_2.INJECT1_0 = "NO";
    defparam phase_accumulator_add_4_2.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i48 (.D(n177_adj_5326), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[48]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i48.GSR = "ENABLED";
    LUT4 phase_increment_1__63__N_21_35__bdd_2_lut_8941 (.A(phase_increment_1__63__N_21[35]), 
         .B(rx_byte[0]), .Z(n19473)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_35__bdd_2_lut_8941.init = 16'heeee;
    LUT4 mux_2289_i1_3_lut (.A(phase_increment_1__63__N_19[12]), .B(phase_increment_1__63__N_20[12]), 
         .C(rx_byte[0]), .Z(n3825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2289_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3624_add_4_33 (.A0(integrator_tmp[66]), .B0(cout_adj_5271), 
          .C0(n93_adj_5969), .D0(n7), .A1(integrator_tmp[67]), .B1(cout_adj_5271), 
          .C1(n90_adj_5968), .D1(n6), .CIN(n17381), .COUT(n17382), .S0(comb6_71__N_1993[66]), 
          .S1(comb6_71__N_1993[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_27 (.A0(integrator_tmp[60]), .B0(cout_adj_5271), 
          .C0(n111_adj_5975), .D0(n13), .A1(integrator_tmp[61]), .B1(cout_adj_5271), 
          .C1(n108_adj_5974), .D1(n12), .CIN(n17378), .COUT(n17379), 
          .S0(comb6_71__N_1993[60]), .S1(comb6_71__N_1993[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_19 (.A0(integrator_tmp[52]), .B0(cout_adj_5271), 
          .C0(n135_adj_5983), .D0(n21), .A1(integrator_tmp[53]), .B1(cout_adj_5271), 
          .C1(n132_adj_5982), .D1(n20), .CIN(n17374), .COUT(n17375), 
          .S0(comb6_71__N_1993[52]), .S1(comb6_71__N_1993[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_25 (.A0(integrator_tmp[58]), .B0(cout_adj_5271), 
          .C0(n117_adj_5977), .D0(n15), .A1(integrator_tmp[59]), .B1(cout_adj_5271), 
          .C1(n114_adj_5976), .D1(n14), .CIN(n17377), .COUT(n17378), 
          .S0(comb6_71__N_1993[58]), .S1(comb6_71__N_1993[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_17 (.A0(integrator_tmp[50]), .B0(cout_adj_5271), 
          .C0(n141_adj_5985), .D0(n23), .A1(integrator_tmp[51]), .B1(cout_adj_5271), 
          .C1(n138_adj_5984), .D1(n22), .CIN(n17373), .COUT(n17374), 
          .S0(comb6_71__N_1993[50]), .S1(comb6_71__N_1993[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_31 (.A0(integrator_tmp[64]), .B0(cout_adj_5271), 
          .C0(n99_adj_5971), .D0(n9), .A1(integrator_tmp[65]), .B1(cout_adj_5271), 
          .C1(n96_adj_5970), .D1(n8), .CIN(n17380), .COUT(n17381), .S0(comb6_71__N_1993[64]), 
          .S1(comb6_71__N_1993[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_23 (.A0(integrator_tmp[56]), .B0(cout_adj_5271), 
          .C0(n123_adj_5979), .D0(n17), .A1(integrator_tmp[57]), .B1(cout_adj_5271), 
          .C1(n120_adj_5978), .D1(n16), .CIN(n17376), .COUT(n17377), 
          .S0(comb6_71__N_1993[56]), .S1(comb6_71__N_1993[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_15 (.A0(integrator_tmp[48]), .B0(cout_adj_5271), 
          .C0(n147_adj_5987), .D0(n25), .A1(integrator_tmp[49]), .B1(cout_adj_5271), 
          .C1(n144_adj_5986), .D1(n24), .CIN(n17372), .COUT(n17373), 
          .S0(comb6_71__N_1993[48]), .S1(comb6_71__N_1993[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_29 (.A0(integrator_tmp[62]), .B0(cout_adj_5271), 
          .C0(n105_adj_5973), .D0(n11), .A1(integrator_tmp[63]), .B1(cout_adj_5271), 
          .C1(n102_adj_5972), .D1(n10), .CIN(n17379), .COUT(n17380), 
          .S0(comb6_71__N_1993[62]), .S1(comb6_71__N_1993[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_21 (.A0(integrator_tmp[54]), .B0(cout_adj_5271), 
          .C0(n129_adj_5981), .D0(n19), .A1(integrator_tmp[55]), .B1(cout_adj_5271), 
          .C1(n126_adj_5980), .D1(n18), .CIN(n17375), .COUT(n17376), 
          .S0(comb6_71__N_1993[54]), .S1(comb6_71__N_1993[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_21.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_38__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[38]), .Z(n19641)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_38__bdd_2_lut_2_lut.init = 16'h4444;
    LUT4 i5009_4_lut (.A(phase_increment_1__63__N_16[11]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[11]), .D(rx_byte[0]), .Z(n3882)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i5009_4_lut.init = 16'hc088;
    LUT4 mux_2324_i1_3_lut (.A(phase_increment_1__63__N_19[11]), .B(phase_increment_1__63__N_20[11]), 
         .C(rx_byte[0]), .Z(n3872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2324_i1_3_lut.init = 16'hcaca;
    FD1S3AX phase_accumulator_e3_i0_i0 (.D(n321), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i0.GSR = "ENABLED";
    CCU2C _add_1_3624_add_4_13 (.A0(integrator_tmp[46]), .B0(cout_adj_5271), 
          .C0(n153_adj_5989), .D0(n27), .A1(integrator_tmp[47]), .B1(cout_adj_5271), 
          .C1(n150_adj_5988), .D1(n26), .CIN(n17371), .COUT(n17372), 
          .S0(comb6_71__N_1993[46]), .S1(comb6_71__N_1993[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_7 (.A0(integrator_tmp[40]), .B0(cout_adj_5271), 
          .C0(n171_adj_5995), .D0(n33), .A1(integrator_tmp[41]), .B1(cout_adj_5271), 
          .C1(n168_adj_5994), .D1(n32), .CIN(n17368), .COUT(n17369), 
          .S0(comb6_71__N_1993[40]), .S1(comb6_71__N_1993[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_5 (.A0(integrator_tmp[38]), .B0(cout_adj_5271), 
          .C0(n177_adj_5997), .D0(n35), .A1(integrator_tmp[39]), .B1(cout_adj_5271), 
          .C1(n174_adj_5996), .D1(n34_adj_5272), .CIN(n17367), .COUT(n17368), 
          .S0(comb6_71__N_1993[38]), .S1(comb6_71__N_1993[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_11 (.A0(integrator_tmp[44]), .B0(cout_adj_5271), 
          .C0(n159_adj_5991), .D0(n29), .A1(integrator_tmp[45]), .B1(cout_adj_5271), 
          .C1(n156_adj_5990), .D1(n28_adj_5274), .CIN(n17370), .COUT(n17371), 
          .S0(comb6_71__N_1993[44]), .S1(comb6_71__N_1993[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_3 (.A0(integrator_tmp[36]), .B0(cout_adj_5271), 
          .C0(n183_adj_5999), .D0(n37), .A1(integrator_tmp[37]), .B1(cout_adj_5271), 
          .C1(n180_adj_5998), .D1(n36), .CIN(n17366), .COUT(n17367), 
          .S0(comb6_71__N_1993[36]), .S1(comb6_71__N_1993[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_37 (.A0(comb6[70]), .B0(cout_adj_6129), .C0(n81_adj_5929), 
          .D0(n3_adj_5304), .A1(comb6[71]), .B1(cout_adj_6129), .C1(n78_adj_5928), 
          .D1(n2_adj_5354), .CIN(n17361), .S0(comb7_71__N_2065[70]), .S1(comb7_71__N_2065[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_9 (.A0(integrator_tmp[42]), .B0(cout_adj_5271), 
          .C0(n165_adj_5993), .D0(n31_adj_5273), .A1(integrator_tmp[43]), 
          .B1(cout_adj_5271), .C1(n162_adj_5992), .D1(n30), .CIN(n17369), 
          .COUT(n17370), .S0(comb6_71__N_1993[42]), .S1(comb6_71__N_1993[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5271), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17366));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3624_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3624_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_1.INJECT1_1 = "NO";
    PFUMX mux_761_i1 (.BLUT(n1757), .ALUT(n1767), .C0(led_0_6), .Z(n1773));
    LUT4 i8189_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19642), 
         .D(n2603), .Z(n2619)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8189_3_lut_4_lut.init = 16'hf780;
    CCU2C _add_1_3798_add_4_38 (.A0(integrator3[71]), .B0(integrator2[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17733), .S0(n78_adj_6245));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3798_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_38.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_32__bdd_2_lut_8646_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[32]), .Z(n19663)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_32__bdd_2_lut_8646_2_lut.init = 16'h4444;
    LUT4 phase_increment_1__63__N_21_37__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[37]), .Z(n19680)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_37__bdd_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_3_lut_3_lut_3_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[3]), 
         .C(rx_byte[2]), .Z(n18645)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i1_3_lut_3_lut_3_lut.init = 16'h0404;
    LUT4 phase_increment_1__63__N_21_30__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[30]), .Z(n19716)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_30__bdd_2_lut_2_lut.init = 16'h4444;
    LUT4 phase_increment_1__63__N_21_28__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[28]), .Z(n19764)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_28__bdd_2_lut_2_lut.init = 16'h4444;
    LUT4 phase_increment_1__63__N_21_60__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[60]), .Z(n19786)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_60__bdd_2_lut_2_lut.init = 16'h4444;
    LUT4 phase_increment_1__63__N_21_58__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[58]), .Z(n19793)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_58__bdd_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_rep_284_2_lut (.A(rx_byte[0]), .B(led_0_6), .Z(n19823)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i1_2_lut_rep_284_2_lut.init = 16'h4444;
    LUT4 phase_increment_1__63__N_21_31__bdd_2_lut_8781 (.A(phase_increment_1__63__N_21[31]), 
         .B(rx_byte[0]), .Z(n19719)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_31__bdd_2_lut_8781.init = 16'heeee;
    LUT4 phase_increment_1__63__N_21_24__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[24]), .Z(n19732)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_24__bdd_2_lut_2_lut.init = 16'h4444;
    LUT4 i8394_4_lut (.A(n18834), .B(rx_byte[0]), .C(rx_byte[5]), .D(rx_byte[2]), 
         .Z(cic_gain_7__N_544[0])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i8394_4_lut.init = 16'h0040;
    LUT4 i8053_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19543), 
         .D(n3919), .Z(n3935)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8053_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut (.A(rx_byte[4]), .B(rx_byte[3]), .C(rx_byte[6]), .D(rx_byte[7]), 
         .Z(n18834)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut.init = 16'hfffd;
    LUT4 i8246_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19493), 
         .D(n1898), .Z(n1914)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8246_3_lut_4_lut.init = 16'hf780;
    LUT4 phase_increment_1__63__N_21_34__bdd_2_lut_8592_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[34]), .Z(n19624)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_34__bdd_2_lut_8592_2_lut.init = 16'h4444;
    LUT4 phase_increment_1__63__N_21_47__bdd_2_lut_8545 (.A(phase_increment_1__63__N_17[47]), 
         .B(led_0_6), .Z(n19553)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_47__bdd_2_lut_8545.init = 16'heeee;
    OB led_pad_6 (.I(led_0_6), .O(led[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(45[22:25])
    OB led_pad_5 (.I(led_0_5), .O(led[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(45[22:25])
    PFUMX mux_1986_i1 (.BLUT(n3402), .ALUT(n3412), .C0(led_0_6), .Z(n3418));
    CCU2C _add_1_3627_add_4_35 (.A0(comb6[68]), .B0(cout_adj_6129), .C0(n87_adj_5931), 
          .D0(n5_adj_5300), .A1(comb6[69]), .B1(cout_adj_6129), .C1(n84_adj_5930), 
          .D1(n4_adj_5301), .CIN(n17360), .COUT(n17361), .S0(comb7_71__N_2065[68]), 
          .S1(comb7_71__N_2065[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_29 (.A0(comb6[62]), .B0(cout_adj_6129), .C0(n105_adj_5937), 
          .D0(n11_adj_5357), .A1(comb6[63]), .B1(cout_adj_6129), .C1(n102_adj_5936), 
          .D1(n10_adj_5356), .CIN(n17357), .COUT(n17358), .S0(comb7_71__N_2065[62]), 
          .S1(comb7_71__N_2065[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_23 (.A0(comb6[56]), .B0(cout_adj_6129), .C0(n123_adj_5943), 
          .D0(n17_adj_5363), .A1(comb6[57]), .B1(cout_adj_6129), .C1(n120_adj_5942), 
          .D1(n16_adj_5362), .CIN(n17354), .COUT(n17355), .S0(comb7_71__N_2065[56]), 
          .S1(comb7_71__N_2065[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_23.INJECT1_1 = "NO";
    LUT4 mux_2382_i1_3_lut (.A(phase_increment_1__63__N_16[9]), .B(phase_increment_1__63__N_18[9]), 
         .C(rx_byte[0]), .Z(n3951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2382_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3627_add_4_27 (.A0(comb6[60]), .B0(cout_adj_6129), .C0(n111_adj_5939), 
          .D0(n13_adj_5359), .A1(comb6[61]), .B1(cout_adj_6129), .C1(n108_adj_5938), 
          .D1(n12_adj_5358), .CIN(n17356), .COUT(n17357), .S0(comb7_71__N_2065[60]), 
          .S1(comb7_71__N_2065[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_33 (.A0(comb6[66]), .B0(cout_adj_6129), .C0(n93_adj_5933), 
          .D0(n7_adj_5294), .A1(comb6[67]), .B1(cout_adj_6129), .C1(n90_adj_5932), 
          .D1(n6_adj_5298), .CIN(n17359), .COUT(n17360), .S0(comb7_71__N_2065[66]), 
          .S1(comb7_71__N_2065[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_25 (.A0(comb6[58]), .B0(cout_adj_6129), .C0(n117_adj_5941), 
          .D0(n15_adj_5361), .A1(comb6[59]), .B1(cout_adj_6129), .C1(n114_adj_5940), 
          .D1(n14_adj_5360), .CIN(n17355), .COUT(n17356), .S0(comb7_71__N_2065[58]), 
          .S1(comb7_71__N_2065[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_21 (.A0(comb6[54]), .B0(cout_adj_6129), .C0(n129_adj_5945), 
          .D0(n19_adj_5365), .A1(comb6[55]), .B1(cout_adj_6129), .C1(n126_adj_5944), 
          .D1(n18_adj_5364), .CIN(n17353), .COUT(n17354), .S0(comb7_71__N_2065[54]), 
          .S1(comb7_71__N_2065[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_31 (.A0(comb6[64]), .B0(cout_adj_6129), .C0(n99_adj_5935), 
          .D0(n9_adj_5355), .A1(comb6[65]), .B1(cout_adj_6129), .C1(n96_adj_5934), 
          .D1(n8_adj_5286), .CIN(n17358), .COUT(n17359), .S0(comb7_71__N_2065[64]), 
          .S1(comb7_71__N_2065[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_31.INJECT1_1 = "NO";
    LUT4 i8029_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n18645), 
         .D(n4258), .Z(n4264)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8029_3_lut_4_lut.init = 16'hf780;
    LUT4 phase_increment_1__63__N_21_16__bdd_2_lut_8886 (.A(phase_increment_1__63__N_21[16]), 
         .B(rx_byte[0]), .Z(n19722)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_16__bdd_2_lut_8886.init = 16'heeee;
    CCU2C _add_1_3798_add_4_36 (.A0(integrator3[69]), .B0(integrator2[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[70]), .B1(integrator2[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17732), .COUT(n17733), .S0(n84_adj_6247), 
          .S1(n81_adj_6246));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3621_add_4_16 (.A0(comb_d9[13]), .B0(comb9[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[14]), .B1(comb9[14]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17391), .COUT(n17392));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_16.INJECT1_1 = "NO";
    OB led_pad_4 (.I(led_0_4), .O(led[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(45[22:25])
    LUT4 i4989_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[17]), 
         .Z(n3580)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4989_2_lut_2_lut.init = 16'h4444;
    PFUMX mux_796_i1 (.BLUT(n1804), .ALUT(n1814), .C0(led_0_6), .Z(n1820));
    LUT4 phase_increment_1__63__N_21_5__bdd_2_lut_8447_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[5]), .Z(n19426)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_5__bdd_2_lut_8447_2_lut.init = 16'h4444;
    OB led_pad_3 (.I(led_0_3), .O(led[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(45[22:25])
    FD1S3AX phase_increment_0__i126 (.D(\phase_increment[0] [61]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i126.GSR = "ENABLED";
    PFUMX i8565 (.BLUT(n19586), .ALUT(n19585), .C0(rx_byte[2]), .Z(n19587));
    LUT4 phase_increment_1__63__N_21_45__bdd_2_lut_8564_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[45]), .Z(n19585)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_45__bdd_2_lut_8564_2_lut.init = 16'h4444;
    LUT4 i8025_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19806), 
         .D(n4154), .Z(n4170)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8025_3_lut_4_lut.init = 16'hf780;
    LUT4 i5001_4_lut (.A(phase_increment_1__63__N_16[13]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[13]), .D(rx_byte[0]), .Z(n3788)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i5001_4_lut.init = 16'hc088;
    LUT4 i8386_4_lut (.A(n18700), .B(n18704), .C(n19819), .D(n19822), 
         .Z(clk_80mhz_enable_238)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(265[5] 289[6])
    defparam i8386_4_lut.init = 16'h5010;
    LUT4 i8180_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19678), 
         .D(n2697), .Z(n2713)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8180_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_912_i1_3_lut (.A(phase_increment_1__63__N_16[51]), .B(phase_increment_1__63__N_18[51]), 
         .C(rx_byte[0]), .Z(n1977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_912_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3642_add_4_7 (.A0(comb_d9[41]), .B0(comb9[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[42]), .B1(comb9[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17255), .COUT(n17256));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_7.INJECT1_1 = "NO";
    FD1S3AX phase_increment_0__i127 (.D(\phase_increment[0] [62]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [62]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i127.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i128 (.D(\phase_increment[0] [63]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i128.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i120 (.D(\phase_increment[0] [55]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i120.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i121 (.D(\phase_increment[0] [56]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [56]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i121.GSR = "ENABLED";
    LUT4 i6755_2_lut (.A(integrator2[0]), .B(integrator1[0]), .Z(integrator2_71__N_1032[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i6755_2_lut.init = 16'h6666;
    FD1S3AX phase_increment_0__i125 (.D(\phase_increment[0] [60]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [60]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i125.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i124 (.D(\phase_increment[0] [59]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i124.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i122 (.D(\phase_increment[0] [57]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i122.GSR = "ENABLED";
    LUT4 phase_increment_1__63__N_21_28__bdd_2_lut_8706_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[28]), .Z(n19763)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_28__bdd_2_lut_8706_2_lut.init = 16'h4444;
    LUT4 mux_2254_i1_3_lut (.A(phase_increment_1__63__N_19[13]), .B(phase_increment_1__63__N_20[13]), 
         .C(rx_byte[0]), .Z(n3778)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2254_i1_3_lut.init = 16'hcaca;
    LUT4 i4984_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[19]), 
         .Z(n3486)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4984_2_lut_2_lut.init = 16'h4444;
    LUT4 i4912_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[50]), 
         .Z(n2029)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4912_2_lut_2_lut.init = 16'h4444;
    LUT4 i8217_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19587), 
         .D(n2274), .Z(n2290)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8217_3_lut_4_lut.init = 16'hf780;
    FD1S3AX phase_increment_0__i123 (.D(\phase_increment[0] [58]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [58]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i123.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i118 (.D(\phase_increment[0] [53]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i118.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i119 (.D(\phase_increment[0] [54]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [54]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i119.GSR = "ENABLED";
    OB led_pad_2 (.I(led_0_2), .O(led[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(45[22:25])
    OB led_pad_1 (.I(led_0_1), .O(led[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(45[22:25])
    CCU2C _add_1_3657_add_4_37 (.A0(comb_d9_adj_6570[71]), .B0(comb9_adj_6569[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16734), .S0(n76));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_37.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_37.INIT1 = 16'h0000;
    defparam _add_1_3657_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_37.INJECT1_1 = "NO";
    IB rx_serial_pad (.I(rx_serial), .O(rx_serial_c));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(39[22:31])
    PFUMX i8562 (.BLUT(n19581), .ALUT(n19580), .C0(rx_byte[2]), .Z(n19582));
    FD1S3AX phase_increment_0__i105 (.D(\phase_increment[0] [40]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [40]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i105.GSR = "ENABLED";
    IB rf_in_pad (.I(rf_in), .O(rf_in_c));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(40[22:27])
    FD1S3AX phase_increment_0__i104 (.D(\phase_increment[0] [39]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i104.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i103 (.D(\phase_increment[0] [38]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [38]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i103.GSR = "ENABLED";
    IB clk_25mhz_pad (.I(clk_25mhz), .O(clk_25mhz_c));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(38[22:31])
    OB led_pad_0 (.I(led_0_0), .O(led[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(45[22:25])
    CCU2C _add_1_3642_add_4_5 (.A0(comb_d9[39]), .B0(comb9[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[40]), .B1(comb9[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17254), .COUT(n17255));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_5.INJECT1_1 = "NO";
    FD1S3AX phase_increment_0__i102 (.D(\phase_increment[0] [37]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i102.GSR = "ENABLED";
    CCU2C _add_1_3798_add_4_34 (.A0(integrator3[67]), .B0(integrator2[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[68]), .B1(integrator2[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17731), .COUT(n17732), .S0(n90_adj_6249), 
          .S1(n87_adj_6248));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_34.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_42__bdd_2_lut_8575_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[42]), .Z(n19601)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_42__bdd_2_lut_8575_2_lut.init = 16'h4444;
    CCU2C _add_1_add_4_22 (.A0(mix_sinewave[11]), .B0(integrator1[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17590), .COUT(n17591), .S0(integrator1_71__N_960[20]), 
          .S1(integrator1_71__N_960[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_add_4_22.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i47 (.D(n180_adj_5341), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i47.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i46 (.D(n183_adj_5295), .CK(clk_80mhz), 
            .Q(phase_accumulator_adj_6545[46]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i46.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i45 (.D(n186), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i45.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i101 (.D(\phase_increment[0] [36]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [36]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i101.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i100 (.D(\phase_increment[0] [35]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i100.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i99 (.D(\phase_increment[0] [34]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i99.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i98 (.D(\phase_increment[0] [33]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i98.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i97 (.D(\phase_increment[0] [32]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i97.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i96 (.D(\phase_increment[0] [31]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i96.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i95 (.D(\phase_increment[0] [30]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i95.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i94 (.D(\phase_increment[0] [29]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i94.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i44 (.D(n189), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[44]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i44.GSR = "ENABLED";
    CCU2C _add_1_3642_add_4_3 (.A0(comb_d9[37]), .B0(comb9[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[38]), .B1(comb9[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17253), .COUT(n17254));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_3642_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_3.INJECT1_1 = "NO";
    FD1S3AX phase_increment_0__i93 (.D(\phase_increment[0] [28]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i93.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i92 (.D(\phase_increment[0] [27]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i92.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i91 (.D(\phase_increment[0] [26]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i91.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i90 (.D(\phase_increment[0] [25]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i90.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i89 (.D(\phase_increment[0] [24]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i89.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i88 (.D(\phase_increment[0] [23]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i88.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i87 (.D(\phase_increment[0] [22]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i87.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i86 (.D(\phase_increment[0] [21]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i86.GSR = "ENABLED";
    LUT4 phase_increment_1__63__N_21_24__bdd_2_lut_8677 (.A(led_0_6), .B(phase_increment_1__63__N_17[24]), 
         .Z(n19731)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_24__bdd_2_lut_8677.init = 16'heeee;
    FD1S3AX phase_increment_0__i85 (.D(\phase_increment[0] [20]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i85.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i84 (.D(\phase_increment[0] [19]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i84.GSR = "ENABLED";
    CCU2C _add_1_add_4_20 (.A0(mix_sinewave[11]), .B0(integrator1[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17589), .COUT(n17590), .S0(integrator1_71__N_960[18]), 
          .S1(integrator1_71__N_960[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_add_4_20.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i43 (.D(n192), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i43.GSR = "ENABLED";
    CCU2C _add_1_add_4_18 (.A0(mix_sinewave[11]), .B0(integrator1[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17588), .COUT(n17589), .S0(integrator1_71__N_960[16]), 
          .S1(integrator1_71__N_960[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_add_4_18.INJECT1_1 = "NO";
    FD1S3AX phase_increment_0__i83 (.D(\phase_increment[0] [18]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i83.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i82 (.D(\phase_increment[0] [17]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i82.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i81 (.D(\phase_increment[0] [16]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i81.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i80 (.D(\phase_increment[0] [15]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i80.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i79 (.D(\phase_increment[0] [14]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i79.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i78 (.D(\phase_increment[0] [13]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i78.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i77 (.D(\phase_increment[0] [12]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i77.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i28 (.D(n237), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i28.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i27 (.D(n240), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i27.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i26 (.D(n243), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i26.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i25 (.D(n246), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i25.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i76 (.D(\phase_increment[0] [11]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i76.GSR = "ENABLED";
    CCU2C _add_1_add_4_16 (.A0(mix_sinewave[11]), .B0(integrator1[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17587), .COUT(n17588), .S0(integrator1_71__N_960[14]), 
          .S1(integrator1_71__N_960[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_add_4_16.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_8__bdd_2_lut_8461_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[8]), .Z(n19440)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_8__bdd_2_lut_8461_2_lut.init = 16'h4444;
    FD1S3AX phase_increment_0__i75 (.D(\phase_increment[0] [10]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i75.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i74 (.D(\phase_increment[0] [9]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i74.GSR = "ENABLED";
    LUT4 mux_1729_i1_3_lut (.A(phase_increment_1__63__N_19[28]), .B(phase_increment_1__63__N_20[28]), 
         .C(rx_byte[0]), .Z(n3073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1729_i1_3_lut.init = 16'hcaca;
    FD1S3AX phase_increment_0__i73 (.D(\phase_increment[0] [8]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i73.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i72 (.D(\phase_increment[0] [7]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i72.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i71 (.D(\phase_increment[0] [6]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i71.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i70 (.D(\phase_increment[0] [5]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i70.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i69 (.D(\phase_increment[0] [4]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i69.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i68 (.D(phase_increment_1__63__N_17[3]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i68.GSR = "ENABLED";
    FD1S3AX phase_increment_0__i67 (.D(phase_increment_1__63__N_17[2]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i67.GSR = "ENABLED";
    LUT4 i8143_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19717), 
         .D(n2979), .Z(n2995)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8143_3_lut_4_lut.init = 16'hf780;
    FD1S3AX phase_increment_0__i66 (.D(phase_increment_1__63__N_17[1]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i66.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i24 (.D(n249), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i24.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i23 (.D(n252), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i23.GSR = "ENABLED";
    CCU2C _add_1_3657_add_4_35 (.A0(comb_d9_adj_6570[69]), .B0(comb9_adj_6569[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[70]), .B1(comb9_adj_6569[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16733), .COUT(n16734), .S0(n82), 
          .S1(n79));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_35.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_35.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_35.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i22 (.D(n255), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i22.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i21 (.D(n258), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i21.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i20 (.D(n261), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i20.GSR = "ENABLED";
    LUT4 i4909_4_lut (.A(phase_increment_1__63__N_16[52]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[52]), .D(rx_byte[0]), .Z(n1955)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4909_4_lut.init = 16'hc088;
    FD1S3AX phase_increment_0__i65 (.D(phase_increment_1__63__N_21[0]), .CK(clk_80mhz), 
            .Q(\phase_increment[1] [0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i65.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i64 (.D(n1447), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i64.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i63 (.D(n1494), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [62]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i63.GSR = "ENABLED";
    CCU2C _add_1_3798_add_4_32 (.A0(integrator3[65]), .B0(integrator2[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[66]), .B1(integrator2[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17730), .COUT(n17731), .S0(n96_adj_6251), 
          .S1(n93_adj_6250));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3798_add_4_30 (.A0(integrator3[63]), .B0(integrator2[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[64]), .B1(integrator2[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17729), .COUT(n17730), .S0(n102_adj_6253), 
          .S1(n99_adj_6252));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3642_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[36]), .B1(comb9[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17253));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3642_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3642_add_4_1.INIT1 = 16'h9995;
    defparam _add_1_3642_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3642_add_4_1.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i62 (.D(n1541), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i62.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i61 (.D(n19791), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [60]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i61.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i60 (.D(n1635), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i60.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i59 (.D(n19798), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [58]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i59.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i58 (.D(n1729), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i58.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i57 (.D(n1776), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [56]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i57.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i56 (.D(n1823), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i56.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i55 (.D(n19425), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [54]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i55.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i54 (.D(n1917), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i54.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i53 (.D(n1964), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [52]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i53.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i52 (.D(n2011), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i52.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i19 (.D(n264), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i19.GSR = "ENABLED";
    CCU2C _add_1_add_4_14 (.A0(mix_sinewave[11]), .B0(integrator1[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17586), .COUT(n17587), .S0(integrator1_71__N_960[12]), 
          .S1(integrator1_71__N_960[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_add_4_14.INJECT1_1 = "NO";
    PFUMX i8559 (.BLUT(n19577), .ALUT(n19576), .C0(led_0_6), .Z(n19578));
    LUT4 i8187_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19649), 
         .D(n2556), .Z(n2572)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8187_3_lut_4_lut.init = 16'hf780;
    FD1S3AX phase_accumulator_e3_i0_i18 (.D(n267), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i18.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i17 (.D(n270), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i17.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i16 (.D(n273), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i16.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i42 (.D(n195), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[42]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i42.GSR = "ENABLED";
    CCU2C _add_1_3798_add_4_28 (.A0(integrator3[61]), .B0(integrator2[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[62]), .B1(integrator2[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17728), .COUT(n17729), .S0(n108_adj_6255), 
          .S1(n105_adj_6254));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_28.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i51 (.D(n2058), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [50]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i51.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i50 (.D(n2105), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i50.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i49 (.D(n2152), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [48]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i49.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i48 (.D(n2199), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i48.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i47 (.D(n2246), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [46]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i47.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i46 (.D(n2293), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i46.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i45 (.D(n2340), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [44]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i45.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i44 (.D(n2387), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i44.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i43 (.D(n2434), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [42]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i43.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i42 (.D(n2481), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i42.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i41 (.D(n2528), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [40]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i41.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i15 (.D(n276), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i15.GSR = "ENABLED";
    CCU2C _add_1_add_4_12 (.A0(mix_sinewave[10]), .B0(integrator1[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_sinewave[11]), .B1(integrator1[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17585), .COUT(n17586), .S0(integrator1_71__N_960[10]), 
          .S1(integrator1_71__N_960[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_add_4_12.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i14 (.D(n279), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i14.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i13 (.D(n282), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i13.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i12 (.D(n285), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i12.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i11 (.D(n288), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i11.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i10 (.D(n291), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i10.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i40 (.D(n2575), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i40.GSR = "ENABLED";
    CCU2C _add_1_3657_add_4_33 (.A0(comb_d9_adj_6570[67]), .B0(comb9_adj_6569[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[68]), .B1(comb9_adj_6569[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16732), .COUT(n16733), .S0(n88), 
          .S1(n85));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_33.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_33.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_33.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i39 (.D(n2622), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [38]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i39.GSR = "ENABLED";
    CCU2C _add_1_3657_add_4_31 (.A0(comb_d9_adj_6570[65]), .B0(comb9_adj_6569[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[66]), .B1(comb9_adj_6569[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16731), .COUT(n16732), .S0(n94), 
          .S1(n91));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_31.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_31.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_31.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i38 (.D(n2669), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i38.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i37 (.D(n2716), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [36]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i37.GSR = "ENABLED";
    CCU2C _add_1_3657_add_4_29 (.A0(comb_d9_adj_6570[63]), .B0(comb9_adj_6569[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[64]), .B1(comb9_adj_6569[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16730), .COUT(n16731), .S0(n100), 
          .S1(n97));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_29.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_29.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_29.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i36 (.D(n2763), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i36.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i35 (.D(n19630), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i35.GSR = "ENABLED";
    CCU2C _add_1_3657_add_4_27 (.A0(comb_d9_adj_6570[61]), .B0(comb9_adj_6569[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[62]), .B1(comb9_adj_6569[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16729), .COUT(n16730), .S0(n106), 
          .S1(n103));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_27.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_27.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_27.INJECT1_1 = "NO";
    PFUMX mux_759_i1 (.BLUT(n1762), .ALUT(n1747), .C0(rx_byte[2]), .Z(n1770));
    FD1P3AX phase_increment_0__i34 (.D(n2857), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i34.GSR = "ENABLED";
    CCU2C _add_1_3657_add_4_25 (.A0(comb_d9_adj_6570[59]), .B0(comb9_adj_6569[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[60]), .B1(comb9_adj_6569[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16728), .COUT(n16729), .S0(n112), 
          .S1(n109));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_25.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_25.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_25.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i33 (.D(n19668), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i33.GSR = "ENABLED";
    CCU2C _add_1_3657_add_4_23 (.A0(comb_d9_adj_6570[57]), .B0(comb9_adj_6569[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[58]), .B1(comb9_adj_6569[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16727), .COUT(n16728), .S0(n118), 
          .S1(n115));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_23.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_23.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_23.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i32 (.D(n2951), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i32.GSR = "ENABLED";
    CCU2C _add_1_3657_add_4_21 (.A0(comb_d9_adj_6570[55]), .B0(comb9_adj_6569[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[56]), .B1(comb9_adj_6569[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16726), .COUT(n16727));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_21.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_21.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_21.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i31 (.D(n2998), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i31.GSR = "ENABLED";
    PFUMX mux_868_i1 (.BLUT(n1908), .ALUT(n1914), .C0(n19297), .Z(n1917));
    CCU2C _add_1_3657_add_4_19 (.A0(comb_d9_adj_6570[53]), .B0(comb9_adj_6569[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[54]), .B1(comb9_adj_6569[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16725), .COUT(n16726));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_19.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_19.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_19.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i30 (.D(n3045), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i30.GSR = "ENABLED";
    CCU2C _add_1_3657_add_4_17 (.A0(comb_d9_adj_6570[51]), .B0(comb9_adj_6569[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[52]), .B1(comb9_adj_6569[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16724), .COUT(n16725));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_17.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_17.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_17.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i29 (.D(n3092), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i29.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i28 (.D(n3139), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i28.GSR = "ENABLED";
    CCU2C _add_1_3657_add_4_15 (.A0(comb_d9_adj_6570[49]), .B0(comb9_adj_6569[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[50]), .B1(comb9_adj_6569[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16723), .COUT(n16724));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_15.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_15.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_15.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i27 (.D(n3186), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i27.GSR = "ENABLED";
    CCU2C _add_1_3657_add_4_13 (.A0(comb_d9_adj_6570[47]), .B0(comb9_adj_6569[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[48]), .B1(comb9_adj_6569[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16722), .COUT(n16723));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_13.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_13.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_13.INJECT1_1 = "NO";
    PFUMX mux_1951_i1 (.BLUT(n3355), .ALUT(n3365), .C0(led_0_6), .Z(n3371));
    LUT4 mux_889_i1_3_lut (.A(phase_increment_1__63__N_19[52]), .B(phase_increment_1__63__N_20[52]), 
         .C(rx_byte[0]), .Z(n1945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_889_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1807_i1_3_lut (.A(rx_byte[2]), .B(n3152), .C(rx_byte[3]), 
         .Z(n3177)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1807_i1_3_lut.init = 16'hcaca;
    LUT4 i8120_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19418), 
         .D(n3120), .Z(n3136)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8120_3_lut_4_lut.init = 16'hf780;
    LUT4 i8122_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19412), 
         .D(n3167), .Z(n3183)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8122_3_lut_4_lut.init = 16'hf780;
    LUT4 i5005_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[11]), 
         .Z(n3862)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i5005_2_lut_2_lut.init = 16'h4444;
    LUT4 i4933_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[41]), 
         .Z(n2452)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4933_2_lut_2_lut.init = 16'h4444;
    LUT4 phase_increment_1__63__N_21_36__bdd_2_lut_8632_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[36]), .Z(n19676)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_36__bdd_2_lut_8632_2_lut.init = 16'h4444;
    FD1P3AX phase_increment_0__i26 (.D(n3233), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i26.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i25 (.D(n19737), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i25.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i24 (.D(n3327), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i24.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i23 (.D(n3374), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i23.GSR = "ENABLED";
    CCU2C _add_1_3645_add_4_37 (.A0(integrator_tmp_adj_6556[70]), .B0(cout_adj_6512), 
          .C0(n81_adj_5762), .D0(n3_adj_5457), .A1(integrator_tmp_adj_6556[71]), 
          .B1(cout_adj_6512), .C1(n78_adj_5761), .D1(n2_adj_5456), .CIN(n17251), 
          .S0(comb6_71__N_1993_adj_6589[70]), .S1(comb6_71__N_1993_adj_6589[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_37.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i22 (.D(n3421), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i22.GSR = "ENABLED";
    PFUMX mux_724_i1 (.BLUT(n1715), .ALUT(n1700), .C0(rx_byte[2]), .Z(n1723));
    FD1P3AX phase_increment_0__i21 (.D(n19436), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i21.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i20 (.D(n3515), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i20.GSR = "ENABLED";
    PFUMX i8443 (.BLUT(n19423), .ALUT(n19422), .C0(led_0_6), .Z(n19424));
    CCU2C _add_1_3627_add_4_19 (.A0(comb6[52]), .B0(cout_adj_6129), .C0(n135_adj_5947), 
          .D0(n21_adj_5367), .A1(comb6[53]), .B1(cout_adj_6129), .C1(n132_adj_5946), 
          .D1(n20_adj_5366), .CIN(n17352), .COUT(n17353), .S0(comb7_71__N_2065[52]), 
          .S1(comb7_71__N_2065[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_13 (.A0(comb6[46]), .B0(cout_adj_6129), .C0(n153_adj_5953), 
          .D0(n27_adj_5373), .A1(comb6[47]), .B1(cout_adj_6129), .C1(n150_adj_5952), 
          .D1(n26_adj_5372), .CIN(n17349), .COUT(n17350), .S0(comb7_71__N_2065[46]), 
          .S1(comb7_71__N_2065[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_5 (.A0(comb6[38]), .B0(cout_adj_6129), .C0(n177_adj_5961), 
          .D0(n35_adj_5381), .A1(comb6[39]), .B1(cout_adj_6129), .C1(n174_adj_5960), 
          .D1(n34_adj_5380), .CIN(n17345), .COUT(n17346), .S0(comb7_71__N_2065[38]), 
          .S1(comb7_71__N_2065[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_11 (.A0(comb6[44]), .B0(cout_adj_6129), .C0(n159_adj_5955), 
          .D0(n29_adj_5375), .A1(comb6[45]), .B1(cout_adj_6129), .C1(n156_adj_5954), 
          .D1(n28_adj_5374), .CIN(n17348), .COUT(n17349), .S0(comb7_71__N_2065[44]), 
          .S1(comb7_71__N_2065[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_3 (.A0(comb6[36]), .B0(cout_adj_6129), .C0(n183_adj_5963), 
          .D0(n37_adj_5383), .A1(comb6[37]), .B1(cout_adj_6129), .C1(n180_adj_5962), 
          .D1(n36_adj_5382), .CIN(n17344), .COUT(n17345), .S0(comb7_71__N_2065[36]), 
          .S1(comb7_71__N_2065[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_17 (.A0(comb6[50]), .B0(cout_adj_6129), .C0(n141_adj_5949), 
          .D0(n23_adj_5369), .A1(comb6[51]), .B1(cout_adj_6129), .C1(n138_adj_5948), 
          .D1(n22_adj_5368), .CIN(n17351), .COUT(n17352), .S0(comb7_71__N_2065[50]), 
          .S1(comb7_71__N_2065[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_9 (.A0(comb6[42]), .B0(cout_adj_6129), .C0(n165_adj_5957), 
          .D0(n31_adj_5377), .A1(comb6[43]), .B1(cout_adj_6129), .C1(n162_adj_5956), 
          .D1(n30_adj_5376), .CIN(n17347), .COUT(n17348), .S0(comb7_71__N_2065[42]), 
          .S1(comb7_71__N_2065[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_6129), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17344));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3627_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3627_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_15 (.A0(comb6[48]), .B0(cout_adj_6129), .C0(n147_adj_5951), 
          .D0(n25_adj_5371), .A1(comb6[49]), .B1(cout_adj_6129), .C1(n144_adj_5950), 
          .D1(n24_adj_5370), .CIN(n17350), .COUT(n17351), .S0(comb7_71__N_2065[48]), 
          .S1(comb7_71__N_2065[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3627_add_4_7 (.A0(comb6[40]), .B0(cout_adj_6129), .C0(n171_adj_5959), 
          .D0(n33_adj_5379), .A1(comb6[41]), .B1(cout_adj_6129), .C1(n168_adj_5958), 
          .D1(n32_adj_5378), .CIN(n17346), .COUT(n17347), .S0(comb7_71__N_2065[40]), 
          .S1(comb7_71__N_2065[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3627_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3627_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3627_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3627_add_4_7.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i19 (.D(n19520), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i19.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i18 (.D(n3609), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i18.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i17 (.D(n3656), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i17.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i16 (.D(n3703), .SP(clk_80mhz_enable_223), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i16.GSR = "ENABLED";
    PFUMX mux_2408_i1 (.BLUT(n3976), .ALUT(n3982), .C0(n19296), .Z(n3985));
    FD1P3AX phase_increment_0__i15 (.D(n19688), .SP(clk_80mhz_enable_235), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i15.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i14 (.D(n3797), .SP(clk_80mhz_enable_235), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i14.GSR = "ENABLED";
    CCU2C _add_1_3630_add_4_34 (.A0(integrator_d_tmp_adj_6557[31]), .B0(integrator_tmp_adj_6556[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[32]), 
          .B1(integrator_tmp_adj_6556[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17338), .COUT(n17339), .S0(comb6_71__N_1993_adj_6589[31]), 
          .S1(comb6_71__N_1993_adj_6589[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_26 (.A0(integrator_d_tmp_adj_6557[23]), .B0(integrator_tmp_adj_6556[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[24]), 
          .B1(integrator_tmp_adj_6556[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17334), .COUT(n17335), .S0(comb6_71__N_1993_adj_6589[23]), 
          .S1(comb6_71__N_1993_adj_6589[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_26.INJECT1_1 = "NO";
    PFUMX i8546 (.BLUT(n19554), .ALUT(n19553), .C0(rx_byte[2]), .Z(n19555));
    CCU2C _add_1_3630_add_4_32 (.A0(integrator_d_tmp_adj_6557[29]), .B0(integrator_tmp_adj_6556[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[30]), 
          .B1(integrator_tmp_adj_6556[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17337), .COUT(n17338), .S0(comb6_71__N_1993_adj_6589[29]), 
          .S1(comb6_71__N_1993_adj_6589[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_24 (.A0(integrator_d_tmp_adj_6557[21]), .B0(integrator_tmp_adj_6556[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[22]), 
          .B1(integrator_tmp_adj_6556[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17333), .COUT(n17334), .S0(comb6_71__N_1993_adj_6589[21]), 
          .S1(comb6_71__N_1993_adj_6589[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_38 (.A0(integrator_d_tmp_adj_6557[35]), .B0(integrator_tmp_adj_6556[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17340), .S0(comb6_71__N_1993_adj_6589[35]), 
          .S1(cout_adj_6512));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3630_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_30 (.A0(integrator_d_tmp_adj_6557[27]), .B0(integrator_tmp_adj_6556[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[28]), 
          .B1(integrator_tmp_adj_6556[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17336), .COUT(n17337), .S0(comb6_71__N_1993_adj_6589[27]), 
          .S1(comb6_71__N_1993_adj_6589[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_22 (.A0(integrator_d_tmp_adj_6557[19]), .B0(integrator_tmp_adj_6556[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[20]), 
          .B1(integrator_tmp_adj_6556[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17332), .COUT(n17333), .S0(comb6_71__N_1993_adj_6589[19]), 
          .S1(comb6_71__N_1993_adj_6589[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_36 (.A0(integrator_d_tmp_adj_6557[33]), .B0(integrator_tmp_adj_6556[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[34]), 
          .B1(integrator_tmp_adj_6556[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17339), .COUT(n17340), .S0(comb6_71__N_1993_adj_6589[33]), 
          .S1(comb6_71__N_1993_adj_6589[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_28 (.A0(integrator_d_tmp_adj_6557[25]), .B0(integrator_tmp_adj_6556[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[26]), 
          .B1(integrator_tmp_adj_6556[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17335), .COUT(n17336), .S0(comb6_71__N_1993_adj_6589[25]), 
          .S1(comb6_71__N_1993_adj_6589[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_28.INJECT1_1 = "NO";
    LUT4 i8027_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19807), 
         .D(n4201), .Z(n4217)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8027_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_2149_i1_3_lut (.A(phase_increment_1__63__N_19[16]), .B(phase_increment_1__63__N_20[16]), 
         .C(rx_byte[0]), .Z(n3637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2149_i1_3_lut.init = 16'hcaca;
    LUT4 i8141_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19720), 
         .D(n2932), .Z(n2948)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8141_3_lut_4_lut.init = 16'hf780;
    CCU2C _add_1_3798_add_4_26 (.A0(integrator3[59]), .B0(integrator2[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[60]), .B1(integrator2[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17727), .COUT(n17728), .S0(n114_adj_6257), 
          .S1(n111_adj_6256));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_26.INJECT1_1 = "NO";
    FD1P3AX phase_increment_0__i13 (.D(n3844), .SP(clk_80mhz_enable_235), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i13.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i12 (.D(n3891), .SP(clk_80mhz_enable_235), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i12.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i11 (.D(n3938), .SP(clk_80mhz_enable_235), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i11.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i10 (.D(n3985), .SP(clk_80mhz_enable_235), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i10.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i9 (.D(n19446), .SP(clk_80mhz_enable_235), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i9.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i8 (.D(n4079), .SP(clk_80mhz_enable_235), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i8.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i7 (.D(n4126), .SP(clk_80mhz_enable_235), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i7.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i6 (.D(n4173), .SP(clk_80mhz_enable_235), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i6.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i5 (.D(n4220), .SP(clk_80mhz_enable_235), 
            .CK(clk_80mhz), .Q(\phase_increment[0] [4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i5.GSR = "ENABLED";
    FD1P3AX phase_increment_0__i4 (.D(n4267), .SP(clk_80mhz_enable_238), 
            .CK(clk_80mhz), .Q(phase_increment_1__63__N_17[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i4.GSR = "ENABLED";
    LUT4 i4996_4_lut (.A(phase_increment_1__63__N_16[15]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[15]), .D(rx_byte[0]), .Z(n3694)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4996_4_lut.init = 16'hc088;
    LUT4 mux_2184_i1_3_lut (.A(phase_increment_1__63__N_19[15]), .B(phase_increment_1__63__N_20[15]), 
         .C(rx_byte[0]), .Z(n3684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2184_i1_3_lut.init = 16'hcaca;
    FD1P3AX phase_increment_0__i3 (.D(n4314), .SP(clk_80mhz_enable_238), 
            .CK(clk_80mhz), .Q(phase_increment_1__63__N_17[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i3.GSR = "ENABLED";
    LUT4 phase_increment_1__63__N_21_14__bdd_2_lut_8638_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[14]), .Z(n19682)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_14__bdd_2_lut_8638_2_lut.init = 16'h4444;
    FD1P3AX phase_increment_0__i2 (.D(n4361), .SP(clk_80mhz_enable_238), 
            .CK(clk_80mhz), .Q(phase_increment_1__63__N_17[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_0__i2.GSR = "ENABLED";
    LUT4 i4999_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[13]), 
         .Z(n3768)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4999_2_lut_2_lut.init = 16'h4444;
    LUT4 n3246_bdd_3_lut_8680 (.A(n3246), .B(rx_byte[2]), .C(rx_byte[3]), 
         .Z(n19734)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n3246_bdd_3_lut_8680.init = 16'hacac;
    LUT4 i8075_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19723), 
         .D(n3637), .Z(n3653)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8075_3_lut_4_lut.init = 16'hf780;
    LUT4 i4867_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[61]), 
         .Z(n1512)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4867_2_lut_2_lut.init = 16'h4444;
    LUT4 phase_increment_1__63__N_21_48__bdd_2_lut_8528_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[48]), .Z(n19524)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_48__bdd_2_lut_8528_2_lut.init = 16'h4444;
    LUT4 mux_1892_i1_3_lut (.A(phase_increment_1__63__N_16[23]), .B(phase_increment_1__63__N_18[23]), 
         .C(rx_byte[0]), .Z(n3293)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1892_i1_3_lut.init = 16'hcaca;
    LUT4 mux_597_i1_3_lut (.A(phase_increment_1__63__N_16[60]), .B(phase_increment_1__63__N_18[60]), 
         .C(rx_byte[0]), .Z(n1554)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_597_i1_3_lut.init = 16'hcaca;
    LUT4 mux_667_i1_3_lut (.A(phase_increment_1__63__N_16[58]), .B(phase_increment_1__63__N_18[58]), 
         .C(rx_byte[0]), .Z(n1648)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_667_i1_3_lut.init = 16'hcaca;
    LUT4 mux_632_i1_3_lut (.A(phase_increment_1__63__N_16[59]), .B(phase_increment_1__63__N_18[59]), 
         .C(rx_byte[0]), .Z(n1601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_632_i1_3_lut.init = 16'hcaca;
    LUT4 n3246_bdd_3_lut (.A(phase_increment_1__63__N_19[24]), .B(phase_increment_1__63__N_20[24]), 
         .C(rx_byte[0]), .Z(n19735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3246_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_2499_i1_3_lut (.A(phase_increment_1__63__N_19[6]), .B(phase_increment_1__63__N_20[6]), 
         .C(rx_byte[0]), .Z(n4107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2499_i1_3_lut.init = 16'hcaca;
    LUT4 i4888_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[57]), 
         .Z(n1700)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4888_2_lut_2_lut.init = 16'h4444;
    LUT4 phase_increment_1__63__N_21_51__bdd_2_lut_8512_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[51]), .Z(n19507)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_51__bdd_2_lut_8512_2_lut.init = 16'h4444;
    LUT4 i4980_2_lut (.A(phase_increment_1__63__N_21[21]), .B(rx_byte[0]), 
         .Z(n3407)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4980_2_lut.init = 16'heeee;
    LUT4 mux_1624_i1_3_lut (.A(phase_increment_1__63__N_19[31]), .B(phase_increment_1__63__N_20[31]), 
         .C(rx_byte[0]), .Z(n2932)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1624_i1_3_lut.init = 16'hcaca;
    PFUMX mux_938_i1 (.BLUT(n2002), .ALUT(n2008), .C0(n19294), .Z(n2011));
    LUT4 mux_1659_i1_3_lut (.A(phase_increment_1__63__N_19[30]), .B(phase_increment_1__63__N_20[30]), 
         .C(rx_byte[0]), .Z(n2979)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1659_i1_3_lut.init = 16'hcaca;
    LUT4 i8241_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19509), 
         .D(n1992), .Z(n2008)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8241_3_lut_4_lut.init = 16'hf780;
    LUT4 i8101_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19582), 
         .D(n3308), .Z(n3324)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8101_3_lut_4_lut.init = 16'hf780;
    FD1S3AX phase_accumulator_e3_i0_i9 (.D(n294), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i9.GSR = "ENABLED";
    LUT4 phase_increment_1__63__N_21_16__bdd_2_lut_8668_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[16]), .Z(n19721)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_16__bdd_2_lut_8668_2_lut.init = 16'h4444;
    LUT4 i8206_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19606), 
         .D(n2368), .Z(n2384)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8206_3_lut_4_lut.init = 16'hf780;
    LUT4 phase_increment_1__63__N_21_53__bdd_2_lut_8501 (.A(phase_increment_1__63__N_17[53]), 
         .B(led_0_6), .Z(n19491)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_53__bdd_2_lut_8501.init = 16'heeee;
    LUT4 phase_increment_1__63__N_21_26__bdd_2_lut_8430_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[26]), .Z(n19410)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_26__bdd_2_lut_8430_2_lut.init = 16'h4444;
    LUT4 phase_increment_1__63__N_21_38__bdd_2_lut_8602_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[38]), .Z(n19640)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_38__bdd_2_lut_8602_2_lut.init = 16'h4444;
    LUT4 mux_1484_i1_3_lut (.A(phase_increment_1__63__N_19[35]), .B(phase_increment_1__63__N_20[35]), 
         .C(rx_byte[0]), .Z(n2744)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1484_i1_3_lut.init = 16'hcaca;
    FD1S3AX phase_accumulator_e3_i0_i8 (.D(n297), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i8.GSR = "ENABLED";
    CCU2C _add_1_add_4_10 (.A0(mix_sinewave[8]), .B0(integrator1[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(mix_sinewave[9]), .B1(integrator1[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17584), .COUT(n17585), .S0(integrator1_71__N_960[8]), 
          .S1(integrator1_71__N_960[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_add_4_10.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i7 (.D(n300), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i7.GSR = "ENABLED";
    LUT4 phase_increment_1__63__N_21_31__bdd_2_lut_8665_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[31]), .Z(n19718)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_31__bdd_2_lut_8665_2_lut.init = 16'h4444;
    LUT4 i4915_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[49]), 
         .Z(n2076)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4915_2_lut_2_lut.init = 16'h4444;
    FD1S3AX phase_accumulator_e3_i0_i6 (.D(n303), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i6.GSR = "ENABLED";
    LUT4 i4893_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[63]), 
         .Z(n1416)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4893_2_lut_2_lut.init = 16'h4444;
    PFUMX mux_901_i1 (.BLUT(n1945), .ALUT(n1955), .C0(led_0_6), .Z(n1961));
    FD1S3AX phase_accumulator_e3_i0_i5 (.D(n306), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i5.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i4 (.D(n309), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i4.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i3 (.D(n312), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i3.GSR = "ENABLED";
    FD1S3AX phase_accumulator_e3_i0_i2 (.D(n315), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i2.GSR = "ENABLED";
    LUT4 mux_1562_i1_3_lut (.A(rx_byte[2]), .B(n2823), .C(rx_byte[3]), 
         .Z(n2848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1562_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_add_4_8 (.A0(mix_sinewave[6]), .B0(integrator1[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(mix_sinewave[7]), .B1(integrator1[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17583), .COUT(n17584), .S0(integrator1_71__N_960[6]), 
          .S1(integrator1_71__N_960[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_add_4_8.INJECT1_1 = "NO";
    LUT4 i6754_2_lut (.A(integrator3[0]), .B(integrator2[0]), .Z(integrator3_71__N_1104[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i6754_2_lut.init = 16'h6666;
    CCU2C _add_1_3633_add_4_37 (.A0(comb7[70]), .B0(cout_adj_6543), .C0(n81_adj_5893), 
          .D0(n3_adj_5385), .A1(comb7[71]), .B1(cout_adj_6543), .C1(n78_adj_5892), 
          .D1(n2_adj_5384), .CIN(n17321), .S0(comb8_71__N_2137[70]), .S1(comb8_71__N_2137[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_10 (.A0(integrator_d_tmp_adj_6557[7]), .B0(integrator_tmp_adj_6556[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[8]), 
          .B1(integrator_tmp_adj_6556[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17326), .COUT(n17327), .S0(comb6_71__N_1993_adj_6589[7]), 
          .S1(comb6_71__N_1993_adj_6589[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_35 (.A0(comb7[68]), .B0(cout_adj_6543), .C0(n87_adj_5895), 
          .D0(n5_adj_5387), .A1(comb7[69]), .B1(cout_adj_6543), .C1(n84_adj_5894), 
          .D1(n4_adj_5386), .CIN(n17320), .COUT(n17321), .S0(comb8_71__N_2137[68]), 
          .S1(comb8_71__N_2137[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_8 (.A0(integrator_d_tmp_adj_6557[5]), .B0(integrator_tmp_adj_6556[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[6]), 
          .B1(integrator_tmp_adj_6556[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17325), .COUT(n17326), .S0(comb6_71__N_1993_adj_6589[5]), 
          .S1(comb6_71__N_1993_adj_6589[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_18 (.A0(integrator_d_tmp_adj_6557[15]), .B0(integrator_tmp_adj_6556[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[16]), 
          .B1(integrator_tmp_adj_6556[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17330), .COUT(n17331), .S0(comb6_71__N_1993_adj_6589[15]), 
          .S1(comb6_71__N_1993_adj_6589[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_18.INJECT1_1 = "NO";
    FD1S3AX phase_accumulator_e3_i0_i1 (.D(n318), .CK(clk_80mhz), .Q(phase_accumulator_adj_6545[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(38[58:93])
    defparam phase_accumulator_e3_i0_i1.GSR = "ENABLED";
    LUT4 i6753_2_lut (.A(integrator4[0]), .B(integrator3[0]), .Z(integrator4_71__N_1176[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i6753_2_lut.init = 16'h6666;
    CCU2C _add_1_add_4_6 (.A0(mix_sinewave[4]), .B0(integrator1[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(mix_sinewave[5]), .B1(integrator1[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17582), .COUT(n17583), .S0(integrator1_71__N_960[4]), 
          .S1(integrator1_71__N_960[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3657_add_4_11 (.A0(comb_d9_adj_6570[45]), .B0(comb9_adj_6569[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[46]), .B1(comb9_adj_6569[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16721), .COUT(n16722));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3645_add_4_35 (.A0(integrator_tmp_adj_6556[68]), .B0(cout_adj_6512), 
          .C0(n87_adj_5764), .D0(n5_adj_5459), .A1(integrator_tmp_adj_6556[69]), 
          .B1(cout_adj_6512), .C1(n84_adj_5763), .D1(n4_adj_5458), .CIN(n17250), 
          .COUT(n17251), .S0(comb6_71__N_1993_adj_6589[68]), .S1(comb6_71__N_1993_adj_6589[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_35.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_23__bdd_2_lut_8561_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[23]), .Z(n19580)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_23__bdd_2_lut_8561_2_lut.init = 16'h4444;
    PFUMX mux_2299_i1 (.BLUT(n3830), .ALUT(n3815), .C0(rx_byte[2]), .Z(n3838));
    CCU2C _add_1_add_4_4 (.A0(mix_sinewave[2]), .B0(integrator1[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(mix_sinewave[3]), .B1(integrator1[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17581), .COUT(n17582), .S0(integrator1_71__N_960[2]), 
          .S1(integrator1_71__N_960[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_add_4_4.INJECT1_1 = "NO";
    \uart_rx(CLKS_PER_BIT=87)  uart_rx_inst (.rx_byte1({rx_byte1}), .clk_80mhz(clk_80mhz), 
            .rx_serial_c(rx_serial_c), .GND_net(GND_net), .VCC_net(VCC_net), 
            .rx_data_valid1(rx_data_valid1)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(245[7] 250[5])
    PFUMX mux_2264_i1 (.BLUT(n3783), .ALUT(n3768), .C0(rx_byte[2]), .Z(n3791));
    CCU2C _add_1_3630_add_4_20 (.A0(integrator_d_tmp_adj_6557[17]), .B0(integrator_tmp_adj_6556[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[18]), 
          .B1(integrator_tmp_adj_6556[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17331), .COUT(n17332), .S0(comb6_71__N_1993_adj_6589[17]), 
          .S1(comb6_71__N_1993_adj_6589[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_12 (.A0(integrator_d_tmp_adj_6557[9]), .B0(integrator_tmp_adj_6556[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[10]), 
          .B1(integrator_tmp_adj_6556[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17327), .COUT(n17328), .S0(comb6_71__N_1993_adj_6589[9]), 
          .S1(comb6_71__N_1993_adj_6589[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_12.INJECT1_1 = "NO";
    LUT4 i6752_2_lut (.A(integrator5[0]), .B(integrator4[0]), .Z(integrator5_71__N_1248[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i6752_2_lut.init = 16'h6666;
    PFUMX mux_794_i1 (.BLUT(n1809), .ALUT(n1794), .C0(rx_byte[2]), .Z(n1817));
    PFUMX mux_1043_i1 (.BLUT(n2143), .ALUT(n2149), .C0(n19296), .Z(n2152));
    PFUMX mux_1006_i1 (.BLUT(n2086), .ALUT(n2096), .C0(led_0_6), .Z(n2102));
    CCU2C _add_1_add_4_2 (.A0(mix_sinewave[0]), .B0(integrator1[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(mix_sinewave[1]), .B1(integrator1[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17581), .S1(integrator1_71__N_960[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_add_4_2.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_4__bdd_2_lut_8742_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[4]), .Z(n19799)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_4__bdd_2_lut_8742_2_lut.init = 16'h4444;
    PFUMX mux_971_i1 (.BLUT(n2039), .ALUT(n2049), .C0(led_0_6), .Z(n2055));
    CCU2C _add_1_3657_add_4_9 (.A0(comb_d9_adj_6570[43]), .B0(comb9_adj_6569[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[44]), .B1(comb9_adj_6569[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16720), .COUT(n16721));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_9.INJECT1_1 = "NO";
    LUT4 mux_1017_i1_3_lut (.A(phase_increment_1__63__N_16[48]), .B(phase_increment_1__63__N_18[48]), 
         .C(rx_byte[0]), .Z(n2118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1017_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3588_add_4_38 (.A0(integrator2_adj_6559[71]), .B0(integrator1_adj_6558[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17579), .S0(n78_adj_6290));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3588_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_36 (.A0(integrator2_adj_6559[69]), .B0(integrator1_adj_6558[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[70]), .B1(integrator1_adj_6558[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17578), .COUT(n17579), .S0(n84_adj_6292), 
          .S1(n81_adj_6291));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3657_add_4_7 (.A0(comb_d9_adj_6570[41]), .B0(comb9_adj_6569[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[42]), .B1(comb9_adj_6569[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16719), .COUT(n16720));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_34 (.A0(integrator2_adj_6559[67]), .B0(integrator1_adj_6558[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[68]), .B1(integrator1_adj_6558[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17577), .COUT(n17578), .S0(n90_adj_6294), 
          .S1(n87_adj_6293));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_34.INJECT1_1 = "NO";
    LUT4 i4979_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[21]), 
         .Z(n3392)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4979_2_lut_2_lut.init = 16'h4444;
    PFUMX mux_899_i1 (.BLUT(n1950), .ALUT(n1935), .C0(rx_byte[2]), .Z(n1958));
    CCU2C _add_1_3588_add_4_32 (.A0(integrator2_adj_6559[65]), .B0(integrator1_adj_6558[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[66]), .B1(integrator1_adj_6558[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17576), .COUT(n17577), .S0(n96_adj_6296), 
          .S1(n93_adj_6295));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3657_add_4_5 (.A0(comb_d9_adj_6570[39]), .B0(comb9_adj_6569[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[40]), .B1(comb9_adj_6569[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16718), .COUT(n16719));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_30 (.A0(integrator2_adj_6559[63]), .B0(integrator1_adj_6558[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[64]), .B1(integrator1_adj_6558[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17575), .COUT(n17576), .S0(n102_adj_6298), 
          .S1(n99_adj_6297));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3657_add_4_3 (.A0(comb_d9_adj_6570[37]), .B0(comb9_adj_6569[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[38]), .B1(comb9_adj_6569[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16717), .COUT(n16718));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_3657_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_28 (.A0(integrator2_adj_6559[61]), .B0(integrator1_adj_6558[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[62]), .B1(integrator1_adj_6558[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17574), .COUT(n17575), .S0(n108_adj_6300), 
          .S1(n105_adj_6299));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_28.INJECT1_1 = "NO";
    LUT4 i4894_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[52]), 
         .Z(n1935)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4894_2_lut_2_lut.init = 16'h4444;
    CCU2C _add_1_3798_add_4_24 (.A0(integrator3[57]), .B0(integrator2[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[58]), .B1(integrator2[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17726), .COUT(n17727), .S0(n120_adj_6259), 
          .S1(n117_adj_6258));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_26 (.A0(integrator2_adj_6559[59]), .B0(integrator1_adj_6558[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[60]), .B1(integrator1_adj_6558[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17573), .COUT(n17574), .S0(n114_adj_6302), 
          .S1(n111_adj_6301));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_26.INJECT1_1 = "NO";
    LUT4 mux_2542_i1_3_lut (.A(rx_byte[2]), .B(n4139), .C(rx_byte[3]), 
         .Z(n4164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2542_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3657_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9_adj_6570[36]), .B1(comb9_adj_6569[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16717));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3657_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3657_add_4_1.INIT1 = 16'h9995;
    defparam _add_1_3657_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3657_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_24 (.A0(integrator2_adj_6559[57]), .B0(integrator1_adj_6558[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[58]), .B1(integrator1_adj_6558[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17572), .COUT(n17573), .S0(n120_adj_6304), 
          .S1(n117_adj_6303));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_24.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_35__bdd_2_lut_8489_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[35]), .Z(n19472)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_35__bdd_2_lut_8489_2_lut.init = 16'h4444;
    CCU2C _add_1_3588_add_4_22 (.A0(integrator2_adj_6559[55]), .B0(integrator1_adj_6558[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[56]), .B1(integrator1_adj_6558[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17571), .COUT(n17572), .S0(n126_adj_6306), 
          .S1(n123_adj_6305));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_22.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_39__bdd_2_lut_8607_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[39]), .Z(n19647)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_39__bdd_2_lut_8607_2_lut.init = 16'h4444;
    CCU2C _add_1_3588_add_4_20 (.A0(integrator2_adj_6559[53]), .B0(integrator1_adj_6558[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[54]), .B1(integrator1_adj_6558[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17570), .COUT(n17571), .S0(n132_adj_6308), 
          .S1(n129_adj_6307));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_20.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_30__bdd_2_lut_8662_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[30]), .Z(n19715)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_30__bdd_2_lut_8662_2_lut.init = 16'h4444;
    CCU2C _add_1_3504_add_4_16 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2410[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2410[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16715), .S1(n36_adj_5310));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3504_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3504_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3504_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3504_add_4_16.INJECT1_1 = "NO";
    PFUMX i8543 (.BLUT(n19551), .ALUT(n19550), .C0(rx_byte[2]), .Z(n19552));
    CCU2C _add_1_3588_add_4_18 (.A0(integrator2_adj_6559[51]), .B0(integrator1_adj_6558[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[52]), .B1(integrator1_adj_6558[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17569), .COUT(n17570), .S0(n138_adj_6310), 
          .S1(n135_adj_6309));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_18.INJECT1_1 = "NO";
    LUT4 n19578_bdd_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19574), 
         .D(n19578), .Z(n19579)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam n19578_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 i5002_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[12]), 
         .Z(n3815)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i5002_2_lut_2_lut.init = 16'h4444;
    CCU2C _add_1_3588_add_4_16 (.A0(integrator2_adj_6559[49]), .B0(integrator1_adj_6558[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[50]), .B1(integrator1_adj_6558[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17568), .COUT(n17569), .S0(n144_adj_6312), 
          .S1(n141_adj_6311));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_14 (.A0(integrator2_adj_6559[47]), .B0(integrator1_adj_6558[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[48]), .B1(integrator1_adj_6558[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17567), .COUT(n17568), .S0(n150_adj_6314), 
          .S1(n147_adj_6313));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_12 (.A0(integrator2_adj_6559[45]), .B0(integrator1_adj_6558[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[46]), .B1(integrator1_adj_6558[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17566), .COUT(n17567), .S0(n156_adj_6316), 
          .S1(n153_adj_6315));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_10 (.A0(integrator2_adj_6559[43]), .B0(integrator1_adj_6558[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[44]), .B1(integrator1_adj_6558[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17565), .COUT(n17566), .S0(n162_adj_6318), 
          .S1(n159_adj_6317));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_8 (.A0(integrator2_adj_6559[41]), .B0(integrator1_adj_6558[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[42]), .B1(integrator1_adj_6558[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17564), .COUT(n17565), .S0(n168_adj_6320), 
          .S1(n165_adj_6319));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_6 (.A0(integrator2_adj_6559[39]), .B0(integrator1_adj_6558[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[40]), .B1(integrator1_adj_6558[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17563), .COUT(n17564), .S0(n174_adj_6322), 
          .S1(n171_adj_6321));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_4 (.A0(integrator2_adj_6559[37]), .B0(integrator1_adj_6558[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[38]), .B1(integrator1_adj_6558[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17562), .COUT(n17563), .S0(n180_adj_6324), 
          .S1(n177_adj_6323));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3588_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3588_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator2_adj_6559[36]), .B1(integrator1_adj_6558[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n17562), .S1(n183_adj_6325));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3588_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3588_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3588_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3588_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3783_add_4_37 (.A0(integrator2[70]), .B0(cout_adj_5296), 
          .C0(n81_adj_6246), .D0(integrator3[70]), .A1(integrator2[71]), 
          .B1(cout_adj_5296), .C1(n78_adj_6245), .D1(integrator3[71]), 
          .CIN(n17560), .S0(integrator3_71__N_1104[70]), .S1(integrator3_71__N_1104[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3783_add_4_35 (.A0(integrator2[68]), .B0(cout_adj_5296), 
          .C0(n87_adj_6248), .D0(integrator3[68]), .A1(integrator2[69]), 
          .B1(cout_adj_5296), .C1(n84_adj_6247), .D1(integrator3[69]), 
          .CIN(n17559), .COUT(n17560), .S0(integrator3_71__N_1104[68]), 
          .S1(integrator3_71__N_1104[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3783_add_4_33 (.A0(integrator2[66]), .B0(cout_adj_5296), 
          .C0(n93_adj_6250), .D0(integrator3[66]), .A1(integrator2[67]), 
          .B1(cout_adj_5296), .C1(n90_adj_6249), .D1(integrator3[67]), 
          .CIN(n17558), .COUT(n17559), .S0(integrator3_71__N_1104[66]), 
          .S1(integrator3_71__N_1104[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_33.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut (.A(led_0_6), .B(rx_byte[2]), .C(n19822), .D(rx_data_valid), 
         .Z(n18700)) /* synthesis lut_function=(!(A (D)+!A !(B (C+!(D))+!B !(D)))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h40ff;
    CCU2C _add_1_3504_add_4_14 (.A0(amdemod_out_d_11__N_2410[9]), .B0(square_sum[25]), 
          .C0(n30_adj_6282), .D0(n13890), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2410[10]), .D1(VCC_net), .CIN(n16714), 
          .COUT(n16715));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3504_add_4_14.INIT0 = 16'h596a;
    defparam _add_1_3504_add_4_14.INIT1 = 16'he1e1;
    defparam _add_1_3504_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3504_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3783_add_4_31 (.A0(integrator2[64]), .B0(cout_adj_5296), 
          .C0(n99_adj_6252), .D0(integrator3[64]), .A1(integrator2[65]), 
          .B1(cout_adj_5296), .C1(n96_adj_6251), .D1(integrator3[65]), 
          .CIN(n17557), .COUT(n17558), .S0(integrator3_71__N_1104[64]), 
          .S1(integrator3_71__N_1104[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3645_add_4_33 (.A0(integrator_tmp_adj_6556[66]), .B0(cout_adj_6512), 
          .C0(n93_adj_5766), .D0(n7_adj_5461), .A1(integrator_tmp_adj_6556[67]), 
          .B1(cout_adj_6512), .C1(n90_adj_5765), .D1(n6_adj_5460), .CIN(n17249), 
          .COUT(n17250), .S0(comb6_71__N_1993_adj_6589[66]), .S1(comb6_71__N_1993_adj_6589[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3504_add_4_12 (.A0(n19815), .B0(amdemod_out_d_11__N_2410[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2410[8]), 
          .B1(amdemod_out_d_11__N_2370[11]), .C1(amdemod_out_d_11__N_2363), 
          .D1(amdemod_out_d_11__N_2369[11]), .CIN(n16713), .COUT(n16714));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3504_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3504_add_4_12.INIT1 = 16'h656a;
    defparam _add_1_3504_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3504_add_4_12.INJECT1_1 = "NO";
    PFUMX mux_2476_i1 (.BLUT(n4060), .ALUT(n4070), .C0(led_0_6), .Z(n4076));
    CCU2C _add_1_3504_add_4_10 (.A0(n19813), .B0(amdemod_out_d_11__N_2410[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2410[6]), 
          .B1(amdemod_out_d_11__N_2380[14]), .C1(n19815), .D1(amdemod_out_d_11__N_2379[14]), 
          .CIN(n16712), .COUT(n16713));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3504_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3504_add_4_10.INIT1 = 16'h656a;
    defparam _add_1_3504_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3504_add_4_10.INJECT1_1 = "NO";
    LUT4 mux_1414_i1_3_lut (.A(phase_increment_1__63__N_19[37]), .B(phase_increment_1__63__N_20[37]), 
         .C(rx_byte[0]), .Z(n2650)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1414_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3504_add_4_8 (.A0(n19811), .B0(amdemod_out_d_11__N_2410[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2410[4]), 
          .B1(amdemod_out_d_11__N_2390[14]), .C1(n19813), .D1(amdemod_out_d_11__N_2389[14]), 
          .CIN(n16711), .COUT(n16712));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3504_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3504_add_4_8.INIT1 = 16'h656a;
    defparam _add_1_3504_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3504_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3798_add_4_22 (.A0(integrator3[55]), .B0(integrator2[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[56]), .B1(integrator2[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17725), .COUT(n17726), .S0(n126_adj_6261), 
          .S1(n123_adj_6260));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3783_add_4_29 (.A0(integrator2[62]), .B0(cout_adj_5296), 
          .C0(n105_adj_6254), .D0(integrator3[62]), .A1(integrator2[63]), 
          .B1(cout_adj_5296), .C1(n102_adj_6253), .D1(integrator3[63]), 
          .CIN(n17556), .COUT(n17557), .S0(integrator3_71__N_1104[62]), 
          .S1(integrator3_71__N_1104[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_29.INJECT1_1 = "NO";
    LUT4 mux_1449_i1_3_lut (.A(phase_increment_1__63__N_19[36]), .B(phase_increment_1__63__N_20[36]), 
         .C(rx_byte[0]), .Z(n2697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1449_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3798_add_4_20 (.A0(integrator3[53]), .B0(integrator2[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[54]), .B1(integrator2[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17724), .COUT(n17725), .S0(n132_adj_6263), 
          .S1(n129_adj_6262));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3783_add_4_27 (.A0(integrator2[60]), .B0(cout_adj_5296), 
          .C0(n111_adj_6256), .D0(integrator3[60]), .A1(integrator2[61]), 
          .B1(cout_adj_5296), .C1(n108_adj_6255), .D1(integrator3[61]), 
          .CIN(n17555), .COUT(n17556), .S0(integrator3_71__N_1104[60]), 
          .S1(integrator3_71__N_1104[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3783_add_4_25 (.A0(integrator2[58]), .B0(cout_adj_5296), 
          .C0(n117_adj_6258), .D0(integrator3[58]), .A1(integrator2[59]), 
          .B1(cout_adj_5296), .C1(n114_adj_6257), .D1(integrator3[59]), 
          .CIN(n17554), .COUT(n17555), .S0(integrator3_71__N_1104[58]), 
          .S1(integrator3_71__N_1104[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3504_add_4_6 (.A0(n19809), .B0(amdemod_out_d_11__N_2410[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2410[2]), 
          .B1(amdemod_out_d_11__N_2400[14]), .C1(n19811), .D1(amdemod_out_d_11__N_2399[14]), 
          .CIN(n16710), .COUT(n16711));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3504_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3504_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_3504_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3504_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3504_add_4_4 (.A0(n19808), .B0(square_sum[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_out_d_11__N_2410[0]), .B1(amdemod_out_d_11__N_2410[14]), 
          .C1(n19809), .D1(amdemod_out_d_11__N_2409[14]), .CIN(n16709), 
          .COUT(n16710));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3504_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3504_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_3504_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3504_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3783_add_4_23 (.A0(integrator2[56]), .B0(cout_adj_5296), 
          .C0(n123_adj_6260), .D0(integrator3[56]), .A1(integrator2[57]), 
          .B1(cout_adj_5296), .C1(n120_adj_6259), .D1(integrator3[57]), 
          .CIN(n17553), .COUT(n17554), .S0(integrator3_71__N_1104[56]), 
          .S1(integrator3_71__N_1104[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_23.INJECT1_1 = "NO";
    LUT4 i4877_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[62]), 
         .Z(n1465)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4877_2_lut_2_lut.init = 16'h4444;
    PFUMX i8538 (.BLUT(n19542), .ALUT(n19541), .C0(rx_byte[2]), .Z(n19543));
    CCU2C _add_1_3783_add_4_21 (.A0(integrator2[54]), .B0(cout_adj_5296), 
          .C0(n129_adj_6262), .D0(integrator3[54]), .A1(integrator2[55]), 
          .B1(cout_adj_5296), .C1(n126_adj_6261), .D1(integrator3[55]), 
          .CIN(n17552), .COUT(n17553), .S0(integrator3_71__N_1104[54]), 
          .S1(integrator3_71__N_1104[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_21.INJECT1_1 = "NO";
    LUT4 mux_1367_i1_3_lut (.A(phase_increment_1__63__N_16[38]), .B(phase_increment_1__63__N_18[38]), 
         .C(rx_byte[0]), .Z(n2588)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1367_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3783_add_4_19 (.A0(integrator2[52]), .B0(cout_adj_5296), 
          .C0(n135_adj_6264), .D0(integrator3[52]), .A1(integrator2[53]), 
          .B1(cout_adj_5296), .C1(n132_adj_6263), .D1(integrator3[53]), 
          .CIN(n17551), .COUT(n17552), .S0(integrator3_71__N_1104[52]), 
          .S1(integrator3_71__N_1104[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_19.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_10__bdd_2_lut_8537_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[10]), .Z(n19541)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_10__bdd_2_lut_8537_2_lut.init = 16'h4444;
    CCU2C _add_1_3504_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16709));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3504_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3504_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3504_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3504_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3783_add_4_17 (.A0(integrator2[50]), .B0(cout_adj_5296), 
          .C0(n141_adj_6266), .D0(integrator3[50]), .A1(integrator2[51]), 
          .B1(cout_adj_5296), .C1(n138_adj_6265), .D1(integrator3[51]), 
          .CIN(n17550), .COUT(n17551), .S0(integrator3_71__N_1104[50]), 
          .S1(integrator3_71__N_1104[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3798_add_4_18 (.A0(integrator3[51]), .B0(integrator2[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[52]), .B1(integrator2[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17723), .COUT(n17724), .S0(n138_adj_6265), 
          .S1(n135_adj_6264));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3567_add_4_37 (.A0(integrator3[70]), .B0(cout_adj_5327), 
          .C0(n81_adj_6094), .D0(integrator4[70]), .A1(integrator3[71]), 
          .B1(cout_adj_5327), .C1(n78_adj_6093), .D1(integrator4[71]), 
          .CIN(n16707), .S0(integrator4_71__N_1176[70]), .S1(integrator4_71__N_1176[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3567_add_4_35 (.A0(integrator3[68]), .B0(cout_adj_5327), 
          .C0(n87_adj_6096), .D0(integrator4[68]), .A1(integrator3[69]), 
          .B1(cout_adj_5327), .C1(n84_adj_6095), .D1(integrator4[69]), 
          .CIN(n16706), .COUT(n16707), .S0(integrator4_71__N_1176[68]), 
          .S1(integrator4_71__N_1176[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_35.INJECT1_1 = "NO";
    FD1S3AX rx_byte_i7 (.D(rx_byte1[7]), .CK(clk_80mhz), .Q(rx_byte[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam rx_byte_i7.GSR = "ENABLED";
    CCU2C _add_1_3783_add_4_15 (.A0(integrator2[48]), .B0(cout_adj_5296), 
          .C0(n147_adj_6268), .D0(integrator3[48]), .A1(integrator2[49]), 
          .B1(cout_adj_5296), .C1(n144_adj_6267), .D1(integrator3[49]), 
          .CIN(n17549), .COUT(n17550), .S0(integrator3_71__N_1104[48]), 
          .S1(integrator3_71__N_1104[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3783_add_4_13 (.A0(integrator2[46]), .B0(cout_adj_5296), 
          .C0(n153_adj_6270), .D0(integrator3[46]), .A1(integrator2[47]), 
          .B1(cout_adj_5296), .C1(n150_adj_6269), .D1(integrator3[47]), 
          .CIN(n17548), .COUT(n17549), .S0(integrator3_71__N_1104[46]), 
          .S1(integrator3_71__N_1104[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3567_add_4_33 (.A0(integrator3[66]), .B0(cout_adj_5327), 
          .C0(n93_adj_6098), .D0(integrator4[66]), .A1(integrator3[67]), 
          .B1(cout_adj_5327), .C1(n90_adj_6097), .D1(integrator4[67]), 
          .CIN(n16705), .COUT(n16706), .S0(integrator4_71__N_1176[66]), 
          .S1(integrator4_71__N_1176[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_33.INJECT1_1 = "NO";
    LUT4 i5004_4_lut_4_lut (.A(rx_byte[3]), .B(rx_byte[0]), .C(phase_increment_1__63__N_18[12]), 
         .D(phase_increment_1__63__N_16[12]), .Z(n3835)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(265[5] 289[6])
    defparam i5004_4_lut_4_lut.init = 16'hf7d5;
    CCU2C _add_1_3567_add_4_31 (.A0(integrator3[64]), .B0(cout_adj_5327), 
          .C0(n99_adj_6100), .D0(integrator4[64]), .A1(integrator3[65]), 
          .B1(cout_adj_5327), .C1(n96_adj_6099), .D1(integrator4[65]), 
          .CIN(n16704), .COUT(n16705), .S0(integrator4_71__N_1176[64]), 
          .S1(integrator4_71__N_1176[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3783_add_4_11 (.A0(integrator2[44]), .B0(cout_adj_5296), 
          .C0(n159_adj_6272), .D0(integrator3[44]), .A1(integrator2[45]), 
          .B1(cout_adj_5296), .C1(n156_adj_6271), .D1(integrator3[45]), 
          .CIN(n17547), .COUT(n17548), .S0(integrator3_71__N_1104[44]), 
          .S1(integrator3_71__N_1104[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3783_add_4_9 (.A0(integrator2[42]), .B0(cout_adj_5296), 
          .C0(n165_adj_6274), .D0(integrator3[42]), .A1(integrator2[43]), 
          .B1(cout_adj_5296), .C1(n162_adj_6273), .D1(integrator3[43]), 
          .CIN(n17546), .COUT(n17547), .S0(integrator3_71__N_1104[42]), 
          .S1(integrator3_71__N_1104[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3798_add_4_16 (.A0(integrator3[49]), .B0(integrator2[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[50]), .B1(integrator2[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17722), .COUT(n17723), .S0(n144_adj_6267), 
          .S1(n141_adj_6266));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_16.INJECT1_1 = "NO";
    LUT4 i4892_2_lut_2_lut (.A(led_0_6), .B(phase_increment_1__63__N_17[55]), 
         .Z(n1794)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i4892_2_lut_2_lut.init = 16'h4444;
    CCU2C _add_1_3798_add_4_14 (.A0(integrator3[47]), .B0(integrator2[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[48]), .B1(integrator2[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17721), .COUT(n17722), .S0(n150_adj_6269), 
          .S1(n147_adj_6268));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_14.INJECT1_1 = "NO";
    FD1S3AX square_sum_e3__i1 (.D(n126_adj_5600), .CK(cic_sine_clk), .Q(square_sum[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i1.GSR = "ENABLED";
    CCU2C _add_1_3783_add_4_7 (.A0(integrator2[40]), .B0(cout_adj_5296), 
          .C0(n171_adj_6276), .D0(integrator3[40]), .A1(integrator2[41]), 
          .B1(cout_adj_5296), .C1(n168_adj_6275), .D1(integrator3[41]), 
          .CIN(n17545), .COUT(n17546), .S0(integrator3_71__N_1104[40]), 
          .S1(integrator3_71__N_1104[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3798_add_4_12 (.A0(integrator3[45]), .B0(integrator2[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[46]), .B1(integrator2[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17720), .COUT(n17721), .S0(n156_adj_6271), 
          .S1(n153_adj_6270));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3645_add_4_31 (.A0(integrator_tmp_adj_6556[64]), .B0(cout_adj_6512), 
          .C0(n99_adj_5768), .D0(n9_adj_5463), .A1(integrator_tmp_adj_6556[65]), 
          .B1(cout_adj_6512), .C1(n96_adj_5767), .D1(n8_adj_5462), .CIN(n17248), 
          .COUT(n17249), .S0(comb6_71__N_1993_adj_6589[64]), .S1(comb6_71__N_1993_adj_6589[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_31.INJECT1_1 = "NO";
    LUT4 i4936_2_lut (.A(phase_increment_1__63__N_17[40]), .B(led_0_6), 
         .Z(n2499)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4936_2_lut.init = 16'heeee;
    CCU2C _add_1_3783_add_4_5 (.A0(integrator2[38]), .B0(cout_adj_5296), 
          .C0(n177_adj_6278), .D0(integrator3[38]), .A1(integrator2[39]), 
          .B1(cout_adj_5296), .C1(n174_adj_6277), .D1(integrator3[39]), 
          .CIN(n17544), .COUT(n17545), .S0(integrator3_71__N_1104[38]), 
          .S1(integrator3_71__N_1104[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_5.INJECT1_1 = "NO";
    LUT4 i4937_2_lut (.A(phase_increment_1__63__N_21[40]), .B(rx_byte[0]), 
         .Z(n2514)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4937_2_lut.init = 16'heeee;
    LUT4 i4991_4_lut (.A(phase_increment_1__63__N_16[17]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[17]), .D(rx_byte[0]), .Z(n3600)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4991_4_lut.init = 16'hc088;
    CCU2C _add_1_3645_add_4_29 (.A0(integrator_tmp_adj_6556[62]), .B0(cout_adj_6512), 
          .C0(n105_adj_5770), .D0(n11_adj_5465), .A1(integrator_tmp_adj_6556[63]), 
          .B1(cout_adj_6512), .C1(n102_adj_5769), .D1(n10_adj_5464), .CIN(n17247), 
          .COUT(n17248), .S0(comb6_71__N_1993_adj_6589[62]), .S1(comb6_71__N_1993_adj_6589[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_29.INJECT1_1 = "NO";
    LUT4 mux_924_i1_3_lut (.A(phase_increment_1__63__N_19[51]), .B(phase_increment_1__63__N_20[51]), 
         .C(rx_byte[0]), .Z(n1992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_924_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3783_add_4_3 (.A0(integrator2[36]), .B0(cout_adj_5296), 
          .C0(n183_adj_6280), .D0(integrator3[36]), .A1(integrator2[37]), 
          .B1(cout_adj_5296), .C1(n180_adj_6279), .D1(integrator3[37]), 
          .CIN(n17543), .COUT(n17544), .S0(integrator3_71__N_1104[36]), 
          .S1(integrator3_71__N_1104[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3783_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3783_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_3.INJECT1_1 = "NO";
    LUT4 mux_1344_i1_3_lut (.A(phase_increment_1__63__N_19[39]), .B(phase_increment_1__63__N_20[39]), 
         .C(rx_byte[0]), .Z(n2556)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1344_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3783_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5296), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17543));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3783_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3783_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3783_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3783_add_4_1.INJECT1_1 = "NO";
    LUT4 i4963_4_lut_4_lut (.A(rx_byte[3]), .B(rx_byte[0]), .C(phase_increment_1__63__N_18[29]), 
         .D(phase_increment_1__63__N_16[29]), .Z(n3036)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(265[5] 289[6])
    defparam i4963_4_lut_4_lut.init = 16'hf7d5;
    CCU2C _add_1_3645_add_4_27 (.A0(integrator_tmp_adj_6556[60]), .B0(cout_adj_6512), 
          .C0(n111_adj_5772), .D0(n13_adj_5467), .A1(integrator_tmp_adj_6556[61]), 
          .B1(cout_adj_6512), .C1(n108_adj_5771), .D1(n12_adj_5466), .CIN(n17246), 
          .COUT(n17247), .S0(comb6_71__N_1993_adj_6589[60]), .S1(comb6_71__N_1993_adj_6589[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_61 (.A0(\phase_increment[0] [63]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17539), .S0(phase_increment_1__63__N_17[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_61.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_61.INIT1 = 16'h0000;
    defparam _add_1_3591_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_61.INJECT1_1 = "NO";
    LUT4 mux_1379_i1_3_lut (.A(phase_increment_1__63__N_19[38]), .B(phase_increment_1__63__N_20[38]), 
         .C(rx_byte[0]), .Z(n2603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1379_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3591_add_4_59 (.A0(\phase_increment[0] [61]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [62]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17538), .COUT(n17539), .S0(phase_increment_1__63__N_17[61]), 
          .S1(phase_increment_1__63__N_17[62]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_59.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_59.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_57 (.A0(\phase_increment[0] [59]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [60]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17537), .COUT(n17538), .S0(phase_increment_1__63__N_17[59]), 
          .S1(phase_increment_1__63__N_17[60]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_57.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_57.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_57.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_25__bdd_2_lut_8495_2_lut (.A(led_0_6), 
         .B(phase_increment_1__63__N_17[25]), .Z(n19478)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam phase_increment_1__63__N_21_25__bdd_2_lut_8495_2_lut.init = 16'h4444;
    LUT4 i5031_3_lut_3_lut (.A(rx_byte[3]), .B(rx_byte[0]), .C(phase_increment_1__63__N_18[2]), 
         .Z(n4305)) /* synthesis lut_function=((B (C))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(265[5] 289[6])
    defparam i5031_3_lut_3_lut.init = 16'hd5d5;
    CCU2C _add_1_3591_add_4_55 (.A0(\phase_increment[0] [57]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [58]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17536), .COUT(n17537), .S0(phase_increment_1__63__N_17[57]), 
          .S1(phase_increment_1__63__N_17[58]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_55.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_55.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_3645_add_4_25 (.A0(integrator_tmp_adj_6556[58]), .B0(cout_adj_6512), 
          .C0(n117_adj_5774), .D0(n15_adj_5469), .A1(integrator_tmp_adj_6556[59]), 
          .B1(cout_adj_6512), .C1(n114_adj_5773), .D1(n14_adj_5468), .CIN(n17245), 
          .COUT(n17246), .S0(comb6_71__N_1993_adj_6589[58]), .S1(comb6_71__N_1993_adj_6589[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_25.INJECT1_1 = "NO";
    PFUMX mux_1113_i1 (.BLUT(n2237), .ALUT(n2243), .C0(n19302), .Z(n2246));
    CCU2C _add_1_3645_add_4_23 (.A0(integrator_tmp_adj_6556[56]), .B0(cout_adj_6512), 
          .C0(n123_adj_5776), .D0(n17_adj_5471), .A1(integrator_tmp_adj_6556[57]), 
          .B1(cout_adj_6512), .C1(n120_adj_5775), .D1(n16_adj_5470), .CIN(n17244), 
          .COUT(n17245), .S0(comb6_71__N_1993_adj_6589[56]), .S1(comb6_71__N_1993_adj_6589[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_23.INJECT1_1 = "NO";
    PFUMX i8529 (.BLUT(n19525), .ALUT(n19524), .C0(rx_byte[2]), .Z(n19526));
    CCU2C _add_1_3591_add_4_53 (.A0(\phase_increment[0] [55]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [56]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17535), .COUT(n17536), .S0(phase_increment_1__63__N_17[55]), 
          .S1(phase_increment_1__63__N_17[56]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_53.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_53.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_53.INJECT1_1 = "NO";
    LUT4 mux_652_i1_3_lut (.A(rx_byte[2]), .B(n1601), .C(rx_byte[3]), 
         .Z(n1626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_652_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3591_add_4_51 (.A0(\phase_increment[0] [53]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [54]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17534), .COUT(n17535), .S0(phase_increment_1__63__N_17[53]), 
          .S1(phase_increment_1__63__N_17[54]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_51.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_51.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_51.INJECT1_1 = "NO";
    LUT4 mux_2114_i1_3_lut (.A(phase_increment_1__63__N_19[17]), .B(phase_increment_1__63__N_20[17]), 
         .C(rx_byte[0]), .Z(n3590)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2114_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3591_add_4_49 (.A0(\phase_increment[0] [51]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [52]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17533), .COUT(n17534), .S0(phase_increment_1__63__N_17[51]), 
          .S1(phase_increment_1__63__N_17[52]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_49.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_49.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_47 (.A0(\phase_increment[0] [49]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [50]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17532), .COUT(n17533), .S0(phase_increment_1__63__N_17[49]), 
          .S1(phase_increment_1__63__N_17[50]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_47.INIT0 = 16'h555f;
    defparam _add_1_3591_add_4_47.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_47.INJECT1_1 = "NO";
    FD1S3AX rx_byte_i6 (.D(rx_byte1[6]), .CK(clk_80mhz), .Q(rx_byte[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam rx_byte_i6.GSR = "ENABLED";
    FD1S3AX rx_byte_i5 (.D(rx_byte1[5]), .CK(clk_80mhz), .Q(rx_byte[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam rx_byte_i5.GSR = "ENABLED";
    FD1S3AX rx_byte_i4 (.D(rx_byte1[4]), .CK(clk_80mhz), .Q(rx_byte[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam rx_byte_i4.GSR = "ENABLED";
    CCU2C _add_1_3591_add_4_45 (.A0(\phase_increment[0] [47]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [48]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17531), .COUT(n17532), .S0(phase_increment_1__63__N_17[47]), 
          .S1(phase_increment_1__63__N_17[48]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_45.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_45.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_45.INJECT1_1 = "NO";
    FD1S3AX rx_byte_i3 (.D(rx_byte1[3]), .CK(clk_80mhz), .Q(rx_byte[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam rx_byte_i3.GSR = "ENABLED";
    LUT4 mux_2604_i1_3_lut (.A(phase_increment_1__63__N_19[3]), .B(phase_increment_1__63__N_20[3]), 
         .C(rx_byte[0]), .Z(n4248)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2604_i1_3_lut.init = 16'hcaca;
    LUT4 mux_2367_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n3904), 
         .Z(n3929)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2367_i1_3_lut_3_lut.init = 16'hd1d1;
    FD1S3AX rx_byte_i2 (.D(rx_byte1[2]), .CK(clk_80mhz), .Q(rx_byte[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam rx_byte_i2.GSR = "ENABLED";
    CCU2C _add_1_3591_add_4_43 (.A0(\phase_increment[0] [45]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [46]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17530), .COUT(n17531), .S0(phase_increment_1__63__N_17[45]), 
          .S1(phase_increment_1__63__N_17[46]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_43.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_43.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_43.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_27__bdd_2_lut_8436 (.A(phase_increment_1__63__N_17[27]), 
         .B(led_0_6), .Z(n19416)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_27__bdd_2_lut_8436.init = 16'heeee;
    PFUMX mux_1078_i1 (.BLUT(n2190), .ALUT(n2196), .C0(n19295), .Z(n2199));
    CCU2C _add_1_3591_add_4_41 (.A0(\phase_increment[0] [43]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [44]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17529), .COUT(n17530), .S0(phase_increment_1__63__N_17[43]), 
          .S1(phase_increment_1__63__N_17[44]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_41.INIT0 = 16'h555f;
    defparam _add_1_3591_add_4_41.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_39 (.A0(\phase_increment[0] [41]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [42]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17528), .COUT(n17529), .S0(phase_increment_1__63__N_17[41]), 
          .S1(phase_increment_1__63__N_17[42]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_39.INIT0 = 16'h555f;
    defparam _add_1_3591_add_4_39.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_37 (.A0(\phase_increment[0] [39]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [40]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17527), .COUT(n17528), .S0(phase_increment_1__63__N_17[39]), 
          .S1(phase_increment_1__63__N_17[40]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_37.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_37.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_35 (.A0(\phase_increment[0] [37]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [38]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17526), .COUT(n17527), .S0(phase_increment_1__63__N_17[37]), 
          .S1(phase_increment_1__63__N_17[38]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_35.INIT0 = 16'h555f;
    defparam _add_1_3591_add_4_35.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_35.INJECT1_1 = "NO";
    LUT4 i4914_4_lut (.A(phase_increment_1__63__N_16[50]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[50]), .D(rx_byte[0]), .Z(n2049)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4914_4_lut.init = 16'hc088;
    CCU2C _add_1_3591_add_4_33 (.A0(\phase_increment[0] [35]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [36]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17525), .COUT(n17526), .S0(phase_increment_1__63__N_17[35]), 
          .S1(phase_increment_1__63__N_17[36]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_33.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_33.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_31 (.A0(\phase_increment[0] [33]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [34]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17524), .COUT(n17525), .S0(phase_increment_1__63__N_17[33]), 
          .S1(phase_increment_1__63__N_17[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_31.INIT0 = 16'h555f;
    defparam _add_1_3591_add_4_31.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_29 (.A0(\phase_increment[0] [31]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [32]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17523), .COUT(n17524), .S0(phase_increment_1__63__N_17[31]), 
          .S1(phase_increment_1__63__N_17[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_29.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_29.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_27 (.A0(\phase_increment[0] [29]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [30]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17522), .COUT(n17523), .S0(phase_increment_1__63__N_17[29]), 
          .S1(phase_increment_1__63__N_17[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_27.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_27.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_25 (.A0(\phase_increment[0] [27]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [28]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17521), .COUT(n17522), .S0(phase_increment_1__63__N_17[27]), 
          .S1(phase_increment_1__63__N_17[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_25.INIT0 = 16'h555f;
    defparam _add_1_3591_add_4_25.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_23 (.A0(\phase_increment[0] [25]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [26]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17520), .COUT(n17521), .S0(phase_increment_1__63__N_17[25]), 
          .S1(phase_increment_1__63__N_17[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_23.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_23.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_23.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_292 (.A(rx_byte[5]), .B(rx_byte[7]), .Z(n19831)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_292.init = 16'h2222;
    CCU2C _add_1_3591_add_4_21 (.A0(\phase_increment[0] [23]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [24]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17519), .COUT(n17520), .S0(phase_increment_1__63__N_17[23]), 
          .S1(phase_increment_1__63__N_17[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_21.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_21.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_21.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_286_3_lut (.A(rx_byte[5]), .B(rx_byte[7]), .C(rx_byte[6]), 
         .Z(n19825)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_rep_286_3_lut.init = 16'h2020;
    LUT4 i4938_4_lut (.A(phase_increment_1__63__N_16[40]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[40]), .D(rx_byte[0]), .Z(n2519)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4938_4_lut.init = 16'hc088;
    LUT4 mux_1309_i1_3_lut (.A(phase_increment_1__63__N_19[40]), .B(phase_increment_1__63__N_20[40]), 
         .C(rx_byte[0]), .Z(n2509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1309_i1_3_lut.init = 16'hcaca;
    LUT4 phase_increment_1__63__N_21_27__bdd_2_lut_8986 (.A(phase_increment_1__63__N_21[27]), 
         .B(rx_byte[0]), .Z(n19417)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_27__bdd_2_lut_8986.init = 16'heeee;
    LUT4 i1_2_lut_rep_283_3_lut_4_lut (.A(rx_byte[5]), .B(rx_byte[7]), .C(n26_adj_5299), 
         .D(rx_byte[6]), .Z(n19822)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_rep_283_3_lut_4_lut.init = 16'h2000;
    LUT4 mux_1694_i1_3_lut (.A(phase_increment_1__63__N_19[29]), .B(phase_increment_1__63__N_20[29]), 
         .C(rx_byte[0]), .Z(n3026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1694_i1_3_lut.init = 16'hcaca;
    LUT4 phase_increment_1__63__N_21_9__bdd_2_lut_8703 (.A(phase_increment_1__63__N_17[9]), 
         .B(led_0_6), .Z(n19760)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_9__bdd_2_lut_8703.init = 16'heeee;
    LUT4 phase_increment_1__63__N_21_9__bdd_2_lut_8799 (.A(phase_increment_1__63__N_21[9]), 
         .B(rx_byte[0]), .Z(n19761)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_9__bdd_2_lut_8799.init = 16'heeee;
    OB pwm_out_p_pad_1 (.I(pwm_out_p_c), .O(pwm_out_p[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(43[22:31])
    OB pwm_out_p_pad_0 (.I(pwm_out_p_c), .O(pwm_out_p[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(43[22:31])
    OB pwm_out_n_pad_3 (.I(GND_net), .O(pwm_out_n[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(44[22:31])
    OB pwm_out_n_pad_2 (.I(GND_net), .O(pwm_out_n[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(44[22:31])
    OB pwm_out_n_pad_1 (.I(GND_net), .O(pwm_out_n[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(44[22:31])
    OB pwm_out_n_pad_0 (.I(GND_net), .O(pwm_out_n[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(44[22:31])
    OB led_pad_7 (.I(GND_net), .O(led[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(45[22:25])
    FD1S3AX rx_byte_i1 (.D(rx_byte1[1]), .CK(clk_80mhz), .Q(led_0_6));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam rx_byte_i1.GSR = "ENABLED";
    LUT4 mux_1387_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n2588), 
         .Z(n2613)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1387_i1_3_lut_3_lut.init = 16'hd1d1;
    LUT4 phase_increment_1__63__N_21_47__bdd_2_lut_8834 (.A(phase_increment_1__63__N_21[47]), 
         .B(rx_byte[0]), .Z(n19554)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_47__bdd_2_lut_8834.init = 16'heeee;
    LUT4 phase_increment_1__63__N_21_60__bdd_2_lut_8725 (.A(led_0_6), .B(phase_increment_1__63__N_17[60]), 
         .Z(n19785)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_60__bdd_2_lut_8725.init = 16'heeee;
    CCU2C _add_1_3567_add_4_29 (.A0(integrator3[62]), .B0(cout_adj_5327), 
          .C0(n105_adj_6102), .D0(integrator4[62]), .A1(integrator3[63]), 
          .B1(cout_adj_5327), .C1(n102_adj_6101), .D1(integrator4[63]), 
          .CIN(n16703), .COUT(n16704), .S0(integrator4_71__N_1176[62]), 
          .S1(integrator4_71__N_1176[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_29.INJECT1_1 = "NO";
    L6MUX21 i8523 (.D0(n19519), .D1(n19516), .SD(n19822), .Z(n19520));
    CCU2C _add_1_3567_add_4_27 (.A0(integrator3[60]), .B0(cout_adj_5327), 
          .C0(n111_adj_6104), .D0(integrator4[60]), .A1(integrator3[61]), 
          .B1(cout_adj_5327), .C1(n108_adj_6103), .D1(integrator4[61]), 
          .CIN(n16702), .COUT(n16703), .S0(integrator4_71__N_1176[60]), 
          .S1(integrator4_71__N_1176[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3567_add_4_25 (.A0(integrator3[58]), .B0(cout_adj_5327), 
          .C0(n117_adj_6106), .D0(integrator4[58]), .A1(integrator3[59]), 
          .B1(cout_adj_5327), .C1(n114_adj_6105), .D1(integrator4[59]), 
          .CIN(n16701), .COUT(n16702), .S0(integrator4_71__N_1176[58]), 
          .S1(integrator4_71__N_1176[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3567_add_4_23 (.A0(integrator3[56]), .B0(cout_adj_5327), 
          .C0(n123_adj_6108), .D0(integrator4[56]), .A1(integrator3[57]), 
          .B1(cout_adj_5327), .C1(n120_adj_6107), .D1(integrator4[57]), 
          .CIN(n16700), .COUT(n16701), .S0(integrator4_71__N_1176[56]), 
          .S1(integrator4_71__N_1176[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_23.INJECT1_1 = "NO";
    LUT4 mux_2137_i1_3_lut (.A(phase_increment_1__63__N_16[16]), .B(phase_increment_1__63__N_18[16]), 
         .C(rx_byte[0]), .Z(n3622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2137_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3567_add_4_21 (.A0(integrator3[54]), .B0(cout_adj_5327), 
          .C0(n129_adj_6110), .D0(integrator4[54]), .A1(integrator3[55]), 
          .B1(cout_adj_5327), .C1(n126_adj_6109), .D1(integrator4[55]), 
          .CIN(n16699), .COUT(n16700), .S0(integrator4_71__N_1176[54]), 
          .S1(integrator4_71__N_1176[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_14 (.A0(integrator_d_tmp_adj_6557[11]), .B0(integrator_tmp_adj_6556[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[12]), 
          .B1(integrator_tmp_adj_6556[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17328), .COUT(n17329), .S0(comb6_71__N_1993_adj_6589[11]), 
          .S1(comb6_71__N_1993_adj_6589[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_19 (.A0(\phase_increment[0] [21]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [22]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17518), .COUT(n17519), .S0(phase_increment_1__63__N_17[21]), 
          .S1(phase_increment_1__63__N_17[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_19.INIT0 = 16'h555f;
    defparam _add_1_3591_add_4_19.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3567_add_4_19 (.A0(integrator3[52]), .B0(cout_adj_5327), 
          .C0(n135_adj_6112), .D0(integrator4[52]), .A1(integrator3[53]), 
          .B1(cout_adj_5327), .C1(n132_adj_6111), .D1(integrator4[53]), 
          .CIN(n16698), .COUT(n16699), .S0(integrator4_71__N_1176[52]), 
          .S1(integrator4_71__N_1176[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3567_add_4_17 (.A0(integrator3[50]), .B0(cout_adj_5327), 
          .C0(n141_adj_6114), .D0(integrator4[50]), .A1(integrator3[51]), 
          .B1(cout_adj_5327), .C1(n138_adj_6113), .D1(integrator4[51]), 
          .CIN(n16697), .COUT(n16698), .S0(integrator4_71__N_1176[50]), 
          .S1(integrator4_71__N_1176[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_4 (.A0(integrator_d_tmp_adj_6557[1]), .B0(integrator_tmp_adj_6556[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[2]), 
          .B1(integrator_tmp_adj_6556[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17323), .COUT(n17324), .S0(comb6_71__N_1993_adj_6589[1]), 
          .S1(comb6_71__N_1993_adj_6589[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_33 (.A0(comb7[66]), .B0(cout_adj_6543), .C0(n93_adj_5897), 
          .D0(n7_adj_5389), .A1(comb7[67]), .B1(cout_adj_6543), .C1(n90_adj_5896), 
          .D1(n6_adj_5388), .CIN(n17319), .COUT(n17320), .S0(comb8_71__N_2137[66]), 
          .S1(comb8_71__N_2137[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_6 (.A0(integrator_d_tmp_adj_6557[3]), .B0(integrator_tmp_adj_6556[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[4]), 
          .B1(integrator_tmp_adj_6556[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17324), .COUT(n17325), .S0(comb6_71__N_1993_adj_6589[3]), 
          .S1(comb6_71__N_1993_adj_6589[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_6.INJECT1_1 = "NO";
    LUT4 mux_862_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n1883), 
         .Z(n1908)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_862_i1_3_lut_3_lut.init = 16'hd1d1;
    CCU2C _add_1_3630_add_4_16 (.A0(integrator_d_tmp_adj_6557[13]), .B0(integrator_tmp_adj_6556[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[14]), 
          .B1(integrator_tmp_adj_6556[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17329), .COUT(n17330), .S0(comb6_71__N_1993_adj_6589[13]), 
          .S1(comb6_71__N_1993_adj_6589[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3630_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3630_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[0]), .B1(integrator_tmp_adj_6556[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n17323), .S1(comb6_71__N_1993_adj_6589[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3630_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3630_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3630_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3630_add_4_2.INJECT1_1 = "NO";
    PFUMX mux_969_i1 (.BLUT(n2044), .ALUT(n2029), .C0(rx_byte[2]), .Z(n2052));
    LUT4 i4865_4_lut (.A(phase_increment_1__63__N_16[61]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[61]), .D(rx_byte[0]), .Z(n1532)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4865_4_lut.init = 16'hc088;
    CCU2C _add_1_3567_add_4_15 (.A0(integrator3[48]), .B0(cout_adj_5327), 
          .C0(n147_adj_6116), .D0(integrator4[48]), .A1(integrator3[49]), 
          .B1(cout_adj_5327), .C1(n144_adj_6115), .D1(integrator4[49]), 
          .CIN(n16696), .COUT(n16697), .S0(integrator4_71__N_1176[48]), 
          .S1(integrator4_71__N_1176[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_15.INJECT1_1 = "NO";
    LUT4 n1554_bdd_3_lut_8728 (.A(n1554), .B(rx_byte[2]), .C(rx_byte[3]), 
         .Z(n19788)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n1554_bdd_3_lut_8728.init = 16'hacac;
    CCU2C _add_1_3567_add_4_13 (.A0(integrator3[46]), .B0(cout_adj_5327), 
          .C0(n153_adj_6118), .D0(integrator4[46]), .A1(integrator3[47]), 
          .B1(cout_adj_5327), .C1(n150_adj_6117), .D1(integrator4[47]), 
          .CIN(n16695), .COUT(n16696), .S0(integrator4_71__N_1176[46]), 
          .S1(integrator4_71__N_1176[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_13.INJECT1_1 = "NO";
    LUT4 n1554_bdd_3_lut (.A(phase_increment_1__63__N_19[60]), .B(phase_increment_1__63__N_20[60]), 
         .C(rx_byte[0]), .Z(n19789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1554_bdd_3_lut.init = 16'hcaca;
    LUT4 phase_increment_1__63__N_21_58__bdd_2_lut_8734 (.A(led_0_6), .B(phase_increment_1__63__N_17[58]), 
         .Z(n19792)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_58__bdd_2_lut_8734.init = 16'heeee;
    CCU2C _add_1_3798_add_4_10 (.A0(integrator3[43]), .B0(integrator2[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[44]), .B1(integrator2[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17719), .COUT(n17720), .S0(n162_adj_6273), 
          .S1(n159_adj_6272));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3567_add_4_11 (.A0(integrator3[44]), .B0(cout_adj_5327), 
          .C0(n159_adj_6120), .D0(integrator4[44]), .A1(integrator3[45]), 
          .B1(cout_adj_5327), .C1(n156_adj_6119), .D1(integrator4[45]), 
          .CIN(n16694), .COUT(n16695), .S0(integrator4_71__N_1176[44]), 
          .S1(integrator4_71__N_1176[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_11.INJECT1_1 = "NO";
    LUT4 n1648_bdd_3_lut_8737 (.A(n1648), .B(rx_byte[2]), .C(rx_byte[3]), 
         .Z(n19795)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n1648_bdd_3_lut_8737.init = 16'hacac;
    CCU2C _add_1_3567_add_4_9 (.A0(integrator3[42]), .B0(cout_adj_5327), 
          .C0(n165_adj_6122), .D0(integrator4[42]), .A1(integrator3[43]), 
          .B1(cout_adj_5327), .C1(n162_adj_6121), .D1(integrator4[43]), 
          .CIN(n16693), .COUT(n16694), .S0(integrator4_71__N_1176[42]), 
          .S1(integrator4_71__N_1176[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_27 (.A0(comb7[60]), .B0(cout_adj_6543), .C0(n111_adj_5903), 
          .D0(n13_adj_5395), .A1(comb7[61]), .B1(cout_adj_6543), .C1(n108_adj_5902), 
          .D1(n12_adj_5394), .CIN(n17316), .COUT(n17317), .S0(comb8_71__N_2137[60]), 
          .S1(comb8_71__N_2137[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3621_add_4_14 (.A0(comb_d9[11]), .B0(comb9[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[12]), .B1(comb9[12]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17390), .COUT(n17391));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_14.INJECT1_1 = "NO";
    LUT4 n1648_bdd_3_lut (.A(phase_increment_1__63__N_19[58]), .B(phase_increment_1__63__N_20[58]), 
         .C(rx_byte[0]), .Z(n19796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1648_bdd_3_lut.init = 16'hcaca;
    LUT4 i5008_2_lut (.A(phase_increment_1__63__N_21[11]), .B(rx_byte[0]), 
         .Z(n3877)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i5008_2_lut.init = 16'heeee;
    LUT4 i4926_2_lut (.A(phase_increment_1__63__N_17[44]), .B(led_0_6), 
         .Z(n2311)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4926_2_lut.init = 16'heeee;
    LUT4 mux_959_i1_3_lut (.A(phase_increment_1__63__N_19[50]), .B(phase_increment_1__63__N_20[50]), 
         .C(rx_byte[0]), .Z(n2039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_959_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3591_add_4_17 (.A0(\phase_increment[0] [19]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [20]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17517), .COUT(n17518), .S0(phase_increment_1__63__N_17[19]), 
          .S1(phase_increment_1__63__N_17[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_17.INIT0 = 16'h555f;
    defparam _add_1_3591_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3567_add_4_7 (.A0(integrator3[40]), .B0(cout_adj_5327), 
          .C0(n171_adj_6124), .D0(integrator4[40]), .A1(integrator3[41]), 
          .B1(cout_adj_5327), .C1(n168_adj_6123), .D1(integrator4[41]), 
          .CIN(n16692), .COUT(n16693), .S0(integrator4_71__N_1176[40]), 
          .S1(integrator4_71__N_1176[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_7.INJECT1_1 = "NO";
    LUT4 mux_1204_i1_3_lut (.A(phase_increment_1__63__N_19[43]), .B(phase_increment_1__63__N_20[43]), 
         .C(rx_byte[0]), .Z(n2368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1204_i1_3_lut.init = 16'hcaca;
    LUT4 mux_574_i1_3_lut (.A(phase_increment_1__63__N_19[61]), .B(phase_increment_1__63__N_20[61]), 
         .C(rx_byte[0]), .Z(n1522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_574_i1_3_lut.init = 16'hcaca;
    LUT4 i4875_4_lut (.A(phase_increment_1__63__N_16[62]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[62]), .D(rx_byte[0]), .Z(n1485)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4875_4_lut.init = 16'hc088;
    LUT4 mux_539_i1_3_lut (.A(phase_increment_1__63__N_19[62]), .B(phase_increment_1__63__N_20[62]), 
         .C(rx_byte[0]), .Z(n1475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_539_i1_3_lut.init = 16'hcaca;
    LUT4 phase_increment_1__63__N_21_54__bdd_2_lut_8439 (.A(phase_increment_1__63__N_17[54]), 
         .B(led_0_6), .Z(n19419)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_54__bdd_2_lut_8439.init = 16'heeee;
    LUT4 led_0_6_bdd_2_lut_8450 (.A(led_0_6), .B(phase_increment_1__63__N_17[20]), 
         .Z(n19429)) /* synthesis lut_function=(A+(B)) */ ;
    defparam led_0_6_bdd_2_lut_8450.init = 16'heeee;
    LUT4 phase_increment_1__63__N_21_54__bdd_2_lut_8482 (.A(phase_increment_1__63__N_21[54]), 
         .B(rx_byte[0]), .Z(n19420)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_54__bdd_2_lut_8482.init = 16'heeee;
    LUT4 mux_1239_i1_3_lut (.A(phase_increment_1__63__N_19[42]), .B(phase_increment_1__63__N_20[42]), 
         .C(rx_byte[0]), .Z(n2415)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1239_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3633_add_4_25 (.A0(comb7[58]), .B0(cout_adj_6543), .C0(n117_adj_5905), 
          .D0(n15_adj_5397), .A1(comb7[59]), .B1(cout_adj_6543), .C1(n114_adj_5904), 
          .D1(n14_adj_5396), .CIN(n17315), .COUT(n17316), .S0(comb8_71__N_2137[58]), 
          .S1(comb8_71__N_2137[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_25.INJECT1_1 = "NO";
    PFUMX mux_1148_i1 (.BLUT(n2284), .ALUT(n2290), .C0(n19300), .Z(n2293));
    CCU2C _add_1_3621_add_4_12 (.A0(comb_d9[9]), .B0(comb9[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[10]), .B1(comb9[10]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17389), .COUT(n17390));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_12.INJECT1_1 = "NO";
    PFUMX i8521 (.BLUT(n19518), .ALUT(n19517), .C0(led_0_6), .Z(n19519));
    LUT4 i6779_2_lut (.A(q_squared[0]), .B(i_squared[0]), .Z(n126_adj_5600)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i6779_2_lut.init = 16'h6666;
    LUT4 i4935_4_lut (.A(phase_increment_1__63__N_16[41]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[41]), .D(rx_byte[0]), .Z(n2472)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4935_4_lut.init = 16'hc088;
    CCU2C _add_1_3567_add_4_5 (.A0(integrator3[38]), .B0(cout_adj_5327), 
          .C0(n177_adj_6126), .D0(integrator4[38]), .A1(integrator3[39]), 
          .B1(cout_adj_5327), .C1(n174_adj_6125), .D1(integrator4[39]), 
          .CIN(n16691), .COUT(n16692), .S0(integrator4_71__N_1176[38]), 
          .S1(integrator4_71__N_1176[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_5.INJECT1_1 = "NO";
    LUT4 mux_1274_i1_3_lut (.A(phase_increment_1__63__N_19[41]), .B(phase_increment_1__63__N_20[41]), 
         .C(rx_byte[0]), .Z(n2462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1274_i1_3_lut.init = 16'hcaca;
    LUT4 i4976_2_lut (.A(phase_increment_1__63__N_17[22]), .B(led_0_6), 
         .Z(n3345)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4976_2_lut.init = 16'heeee;
    LUT4 i1_3_lut (.A(rx_byte[3]), .B(rx_byte[2]), .C(rx_byte[4]), .Z(n18533)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut.init = 16'h1010;
    CCU2C _add_1_3591_add_4_15 (.A0(\phase_increment[0] [17]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [18]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17516), .COUT(n17517), .S0(phase_increment_1__63__N_17[17]), 
          .S1(phase_increment_1__63__N_17[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_15.INJECT1_1 = "NO";
    LUT4 i4977_2_lut (.A(phase_increment_1__63__N_21[22]), .B(rx_byte[0]), 
         .Z(n3360)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4977_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_240 (.A(n19823), .B(n18533), .C(n19831), .D(rx_byte[6]), 
         .Z(cic_gain_7__N_544[1])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_4_lut_adj_240.init = 16'h0080;
    LUT4 led_0_6_bdd_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[20]), 
         .Z(n19430)) /* synthesis lut_function=(A+(B)) */ ;
    defparam led_0_6_bdd_2_lut.init = 16'heeee;
    LUT4 mux_1772_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n3105), 
         .Z(n3130)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1772_i1_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i1_3_lut_rep_280_4_lut (.A(rx_byte[6]), .B(n19831), .C(n45), 
         .D(n26_adj_5299), .Z(n19819)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_3_lut_rep_280_4_lut.init = 16'h8880;
    LUT4 mux_1737_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n3058), 
         .Z(n3083)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1737_i1_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_2402_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n3951), 
         .Z(n3976)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2402_i1_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i6782_2_lut (.A(mix_sinewave[0]), .B(integrator1[0]), .Z(integrator1_71__N_960[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i6782_2_lut.init = 16'h6666;
    CCU2C _add_1_3633_add_4_23 (.A0(comb7[56]), .B0(cout_adj_6543), .C0(n123_adj_5907), 
          .D0(n17_adj_5399), .A1(comb7[57]), .B1(cout_adj_6543), .C1(n120_adj_5906), 
          .D1(n16_adj_5398), .CIN(n17314), .COUT(n17315), .S0(comb8_71__N_2137[56]), 
          .S1(comb8_71__N_2137[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_23.INJECT1_1 = "NO";
    LUT4 mux_1422_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n2635), 
         .Z(n2660)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1422_i1_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i6759_2_lut (.A(integrator2_adj_6559[0]), .B(integrator1_adj_6558[0]), 
         .Z(integrator2_71__N_1032_adj_6574[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i6759_2_lut.init = 16'h6666;
    CCU2C _add_1_3621_add_4_10 (.A0(comb_d9[7]), .B0(comb9[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[8]), .B1(comb9[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17388), .COUT(n17389));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3621_add_4_8 (.A0(comb_d9[5]), .B0(comb9[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[6]), .B1(comb9[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17387), .COUT(n17388));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_8.INJECT1_1 = "NO";
    LUT4 i4882_4_lut (.A(phase_increment_1__63__N_16[63]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[63]), .D(rx_byte[0]), .Z(n1438)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4882_4_lut.init = 16'hc088;
    LUT4 i6758_2_lut (.A(integrator3_adj_6560[0]), .B(integrator2_adj_6559[0]), 
         .Z(integrator3_71__N_1104_adj_6575[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i6758_2_lut.init = 16'h6666;
    LUT4 mux_504_i1_3_lut (.A(phase_increment_1__63__N_19[63]), .B(phase_increment_1__63__N_20[63]), 
         .C(rx_byte[0]), .Z(n1428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_504_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1134_i1_3_lut (.A(phase_increment_1__63__N_19[45]), .B(phase_increment_1__63__N_20[45]), 
         .C(rx_byte[0]), .Z(n2274)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1134_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3591_add_4_13 (.A0(\phase_increment[0] [15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [16]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17515), .COUT(n17516), .S0(phase_increment_1__63__N_17[15]), 
          .S1(phase_increment_1__63__N_17[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_13.INIT0 = 16'h555f;
    defparam _add_1_3591_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_13.INJECT1_1 = "NO";
    LUT4 i6757_2_lut (.A(integrator4_adj_6561[0]), .B(integrator3_adj_6560[0]), 
         .Z(integrator4_71__N_1176_adj_6576[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i6757_2_lut.init = 16'h6666;
    LUT4 mux_994_i1_3_lut (.A(phase_increment_1__63__N_19[49]), .B(phase_increment_1__63__N_20[49]), 
         .C(rx_byte[0]), .Z(n2086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_994_i1_3_lut.init = 16'hcaca;
    LUT4 i6756_2_lut (.A(integrator5_adj_6562[0]), .B(integrator4_adj_6561[0]), 
         .Z(integrator5_71__N_1248_adj_6577[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i6756_2_lut.init = 16'h6666;
    PFUMX mux_1743_i1 (.BLUT(n3083), .ALUT(n3089), .C0(n19301), .Z(n3092));
    PFUMX mux_2056_i1 (.BLUT(n3496), .ALUT(n3506), .C0(led_0_6), .Z(n3512));
    LUT4 i4928_4_lut (.A(phase_increment_1__63__N_16[44]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[44]), .D(rx_byte[0]), .Z(n2331)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4928_4_lut.init = 16'hc088;
    LUT4 mux_1169_i1_3_lut (.A(phase_increment_1__63__N_19[44]), .B(phase_increment_1__63__N_20[44]), 
         .C(rx_byte[0]), .Z(n2321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1169_i1_3_lut.init = 16'hcaca;
    LUT4 i8341_rep_191_2_lut_3_lut_4_lut (.A(rx_byte[6]), .B(n19831), .C(led_0_6), 
         .D(n26_adj_5299), .Z(n19295)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i8341_rep_191_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i4986_4_lut (.A(phase_increment_1__63__N_16[19]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[19]), .D(rx_byte[0]), .Z(n3506)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4986_4_lut.init = 16'hc088;
    LUT4 mux_1212_i1_3_lut (.A(rx_byte[2]), .B(n2353), .C(rx_byte[3]), 
         .Z(n2378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1212_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1247_i1_3_lut (.A(rx_byte[2]), .B(n2400), .C(rx_byte[3]), 
         .Z(n2425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1247_i1_3_lut.init = 16'hcaca;
    LUT4 phase_increment_1__63__N_21_18__bdd_2_lut_8517 (.A(led_0_6), .B(phase_increment_1__63__N_17[18]), 
         .Z(n19514)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_18__bdd_2_lut_8517.init = 16'heeee;
    LUT4 mux_2394_i1_3_lut (.A(phase_increment_1__63__N_19[9]), .B(phase_increment_1__63__N_20[9]), 
         .C(rx_byte[0]), .Z(n3966)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2394_i1_3_lut.init = 16'hcaca;
    LUT4 i4916_2_lut (.A(phase_increment_1__63__N_21[49]), .B(rx_byte[0]), 
         .Z(n2091)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4916_2_lut.init = 16'heeee;
    PFUMX i8518 (.BLUT(n19515), .ALUT(n19514), .C0(rx_byte[2]), .Z(n19516));
    LUT4 mux_2044_i1_3_lut (.A(phase_increment_1__63__N_19[19]), .B(phase_increment_1__63__N_20[19]), 
         .C(rx_byte[0]), .Z(n3496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2044_i1_3_lut.init = 16'hcaca;
    LUT4 phase_increment_1__63__N_21_34__bdd_2_lut (.A(phase_increment_1__63__N_21[34]), 
         .B(rx_byte[0]), .Z(n19625)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_34__bdd_2_lut.init = 16'heeee;
    CCU2C _add_1_3621_add_4_6 (.A0(comb_d9[3]), .B0(comb9[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[4]), .B1(comb9[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17386), .COUT(n17387));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_6.INJECT1_1 = "NO";
    LUT4 i8341_rep_195_2_lut_3_lut_4_lut (.A(rx_byte[6]), .B(n19831), .C(led_0_6), 
         .D(n26_adj_5299), .Z(n19299)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i8341_rep_195_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 mux_1904_i1_3_lut (.A(phase_increment_1__63__N_19[23]), .B(phase_increment_1__63__N_20[23]), 
         .C(rx_byte[0]), .Z(n3308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1904_i1_3_lut.init = 16'hcaca;
    LUT4 i8341_rep_193_2_lut_3_lut_4_lut (.A(rx_byte[6]), .B(n19831), .C(led_0_6), 
         .D(n26_adj_5299), .Z(n19297)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i8341_rep_193_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 phase_increment_1__63__N_21_46__bdd_2_lut_8542 (.A(phase_increment_1__63__N_17[46]), 
         .B(led_0_6), .Z(n19550)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_46__bdd_2_lut_8542.init = 16'heeee;
    CCU2C _add_1_3591_add_4_11 (.A0(\phase_increment[0] [13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17514), .COUT(n17515), .S0(phase_increment_1__63__N_17[13]), 
          .S1(phase_increment_1__63__N_17[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_11.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_11.INJECT1_1 = "NO";
    LUT4 i4115_2_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n45), .D(rx_data_valid), 
         .Z(clk_80mhz_enable_235)) /* synthesis lut_function=(A (B (D))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(265[5] 289[6])
    defparam i4115_2_lut_4_lut.init = 16'hc800;
    LUT4 i8341_rep_197_2_lut_3_lut_4_lut (.A(rx_byte[6]), .B(n19831), .C(led_0_6), 
         .D(n26_adj_5299), .Z(n19301)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i8341_rep_197_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i6751_2_lut (.A(mix_cosinewave[0]), .B(integrator1_adj_6558[0]), 
         .Z(integrator1_71__N_960_adj_6573[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i6751_2_lut.init = 16'h6666;
    LUT4 mux_1064_i1_3_lut (.A(phase_increment_1__63__N_19[47]), .B(phase_increment_1__63__N_20[47]), 
         .C(rx_byte[0]), .Z(n2180)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1064_i1_3_lut.init = 16'hcaca;
    LUT4 n3528_bdd_3_lut_8520 (.A(n3528), .B(rx_byte[2]), .C(rx_byte[3]), 
         .Z(n19517)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n3528_bdd_3_lut_8520.init = 16'hacac;
    LUT4 n3528_bdd_3_lut (.A(phase_increment_1__63__N_19[18]), .B(phase_increment_1__63__N_20[18]), 
         .C(rx_byte[0]), .Z(n19518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3528_bdd_3_lut.init = 16'hcaca;
    LUT4 i8341_rep_194_2_lut_3_lut_4_lut (.A(rx_byte[6]), .B(n19831), .C(led_0_6), 
         .D(n26_adj_5299), .Z(n19298)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i8341_rep_194_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i8341_rep_190_2_lut_3_lut_4_lut (.A(rx_byte[6]), .B(n19831), .C(led_0_6), 
         .D(n26_adj_5299), .Z(n19294)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i8341_rep_190_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 mux_1099_i1_3_lut (.A(phase_increment_1__63__N_19[46]), .B(phase_increment_1__63__N_20[46]), 
         .C(rx_byte[0]), .Z(n2227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1099_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1612_i1_3_lut (.A(phase_increment_1__63__N_16[31]), .B(phase_increment_1__63__N_18[31]), 
         .C(rx_byte[0]), .Z(n2917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1612_i1_3_lut.init = 16'hcaca;
    LUT4 i8341_rep_198_2_lut_3_lut_4_lut (.A(rx_byte[6]), .B(n19831), .C(led_0_6), 
         .D(n26_adj_5299), .Z(n19302)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i8341_rep_198_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i8341_rep_196_2_lut_3_lut_4_lut (.A(rx_byte[6]), .B(n19831), .C(led_0_6), 
         .D(n26_adj_5299), .Z(n19300)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i8341_rep_196_2_lut_3_lut_4_lut.init = 16'h8f0f;
    PFUMX mux_1004_i1 (.BLUT(n2091), .ALUT(n2076), .C0(rx_byte[2]), .Z(n2099));
    LUT4 i8380_2_lut_3_lut_4_lut (.A(rx_byte[6]), .B(n19831), .C(led_0_6), 
         .D(n26_adj_5299), .Z(n19134)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i8380_2_lut_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_1037_i1_3_lut (.A(rx_byte[2]), .B(n2118), .C(rx_byte[3]), 
         .Z(n2143)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1037_i1_3_lut.init = 16'hcaca;
    LUT4 i5020_4_lut (.A(phase_increment_1__63__N_16[7]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[7]), .D(rx_byte[0]), .Z(n4070)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i5020_4_lut.init = 16'hc088;
    CCU2C _add_1_3567_add_4_3 (.A0(integrator3[36]), .B0(cout_adj_5327), 
          .C0(n183_adj_6128), .D0(integrator4[36]), .A1(integrator3[37]), 
          .B1(cout_adj_5327), .C1(n180_adj_6127), .D1(integrator4[37]), 
          .CIN(n16690), .COUT(n16691), .S0(integrator4_71__N_1176[36]), 
          .S1(integrator4_71__N_1176[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3567_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3567_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_31 (.A0(comb7[64]), .B0(cout_adj_6543), .C0(n99_adj_5899), 
          .D0(n9_adj_5391), .A1(comb7[65]), .B1(cout_adj_6543), .C1(n96_adj_5898), 
          .D1(n8_adj_5390), .CIN(n17318), .COUT(n17319), .S0(comb8_71__N_2137[64]), 
          .S1(comb8_71__N_2137[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_31.INJECT1_1 = "NO";
    PFUMX mux_1253_i1 (.BLUT(n2425), .ALUT(n2431), .C0(n19298), .Z(n2434));
    LUT4 mux_1107_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n2212), 
         .Z(n2237)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1107_i1_3_lut_3_lut.init = 16'hd1d1;
    CCU2C _add_1_3591_add_4_9 (.A0(\phase_increment[0] [11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17513), .COUT(n17514), .S0(phase_increment_1__63__N_17[11]), 
          .S1(phase_increment_1__63__N_17[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_9.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_9.INJECT1_1 = "NO";
    LUT4 mux_2157_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n3622), 
         .Z(n3647)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2157_i1_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i4978_4_lut (.A(phase_increment_1__63__N_16[22]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[22]), .D(rx_byte[0]), .Z(n3365)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4978_4_lut.init = 16'hc088;
    LUT4 n1836_bdd_3_lut_8442 (.A(n1836), .B(rx_byte[2]), .C(rx_byte[3]), 
         .Z(n19422)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n1836_bdd_3_lut_8442.init = 16'hacac;
    LUT4 mux_2464_i1_3_lut (.A(phase_increment_1__63__N_19[7]), .B(phase_increment_1__63__N_20[7]), 
         .C(rx_byte[0]), .Z(n4060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2464_i1_3_lut.init = 16'hcaca;
    LUT4 i4913_2_lut (.A(phase_increment_1__63__N_21[50]), .B(rx_byte[0]), 
         .Z(n2044)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4913_2_lut.init = 16'heeee;
    LUT4 phase_increment_1__63__N_16_20__bdd_3_lut_8453 (.A(phase_increment_1__63__N_16[20]), 
         .B(rx_byte[0]), .C(phase_increment_1__63__N_18[20]), .Z(n19432)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam phase_increment_1__63__N_16_20__bdd_3_lut_8453.init = 16'he2e2;
    PFUMX mux_1218_i1 (.BLUT(n2378), .ALUT(n2384), .C0(n19298), .Z(n2387));
    LUT4 mux_1029_i1_3_lut (.A(phase_increment_1__63__N_19[48]), .B(phase_increment_1__63__N_20[48]), 
         .C(rx_byte[0]), .Z(n2133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1029_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1912_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n3293), 
         .Z(n3318)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1912_i1_3_lut_3_lut.init = 16'hd1d1;
    CCU2C _add_1_3621_add_4_4 (.A0(comb_d9[1]), .B0(comb9[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[2]), .B1(comb9[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17385), .COUT(n17386));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_4.INJECT1_1 = "NO";
    LUT4 mux_1332_i1_3_lut (.A(phase_increment_1__63__N_16[39]), .B(phase_increment_1__63__N_18[39]), 
         .C(rx_byte[0]), .Z(n2541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1332_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1072_i1_3_lut (.A(rx_byte[2]), .B(n2165), .C(rx_byte[3]), 
         .Z(n2190)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1072_i1_3_lut.init = 16'hcaca;
    LUT4 i8341_rep_192_2_lut_3_lut_4_lut (.A(rx_byte[6]), .B(n19831), .C(led_0_6), 
         .D(n26_adj_5299), .Z(n19296)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i8341_rep_192_2_lut_3_lut_4_lut.init = 16'h8f0f;
    CCU2C _add_1_3591_add_4_7 (.A0(\phase_increment[0] [9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17512), .COUT(n17513), .S0(phase_increment_1__63__N_17[9]), 
          .S1(phase_increment_1__63__N_17[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_3591_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_7.INJECT1_1 = "NO";
    PFUMX mux_1181_i1 (.BLUT(n2321), .ALUT(n2331), .C0(led_0_6), .Z(n2337));
    LUT4 phase_increment_1__63__N_16_20__bdd_3_lut (.A(phase_increment_1__63__N_19[20]), 
         .B(phase_increment_1__63__N_20[20]), .C(rx_byte[0]), .Z(n19434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam phase_increment_1__63__N_16_20__bdd_3_lut.init = 16'hcaca;
    LUT4 mux_932_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n1977), 
         .Z(n2002)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_932_i1_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_1142_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n2259), 
         .Z(n2284)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1142_i1_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_807_i1_3_lut (.A(phase_increment_1__63__N_16[54]), .B(phase_increment_1__63__N_18[54]), 
         .C(rx_byte[0]), .Z(n1836)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_807_i1_3_lut.init = 16'hcaca;
    LUT4 mux_2684_i1_4_lut (.A(phase_increment_1__63__N_21[1]), .B(led_0_6), 
         .C(rx_byte[2]), .D(rx_byte[0]), .Z(n4355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2684_i1_4_lut.init = 16'hcfca;
    PFUMX i8513 (.BLUT(n19508), .ALUT(n19507), .C0(rx_byte[2]), .Z(n19509));
    PFUMX i8440 (.BLUT(n19420), .ALUT(n19419), .C0(rx_byte[2]), .Z(n19421));
    LUT4 mux_1087_i1_3_lut (.A(phase_increment_1__63__N_16[46]), .B(phase_increment_1__63__N_18[46]), 
         .C(rx_byte[0]), .Z(n2212)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1087_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3591_add_4_5 (.A0(\phase_increment[0] [7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17511), .COUT(n17512), .S0(phase_increment_1__63__N_17[7]), 
          .S1(phase_increment_1__63__N_17[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_3591_add_4_5.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_5.INJECT1_1 = "NO";
    LUT4 mux_2639_i1_3_lut (.A(phase_increment_1__63__N_19[2]), .B(phase_increment_1__63__N_20[2]), 
         .C(rx_byte[0]), .Z(n4295)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2639_i1_3_lut.init = 16'hcaca;
    LUT4 mux_854_i1_3_lut (.A(phase_increment_1__63__N_19[53]), .B(phase_increment_1__63__N_20[53]), 
         .C(rx_byte[0]), .Z(n1898)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_854_i1_3_lut.init = 16'hcaca;
    LUT4 mux_2359_i1_3_lut (.A(phase_increment_1__63__N_19[10]), .B(phase_increment_1__63__N_20[10]), 
         .C(rx_byte[0]), .Z(n3919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2359_i1_3_lut.init = 16'hcaca;
    LUT4 i6762_2_lut (.A(\phase_increment[1] [0]), .B(phase_accumulator_adj_6545[0]), 
         .Z(n321)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i6762_2_lut.init = 16'h6666;
    LUT4 i4887_2_lut (.A(phase_increment_1__63__N_21[57]), .B(rx_byte[0]), 
         .Z(n1715)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4887_2_lut.init = 16'heeee;
    CCU2C _add_1_3798_add_4_8 (.A0(integrator3[41]), .B0(integrator2[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[42]), .B1(integrator2[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17718), .COUT(n17719), .S0(n168_adj_6275), 
          .S1(n165_adj_6274));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_8.INJECT1_1 = "NO";
    LUT4 mux_1052_i1_3_lut (.A(phase_increment_1__63__N_16[47]), .B(phase_increment_1__63__N_18[47]), 
         .C(rx_byte[0]), .Z(n2165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1052_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3591_add_4_3 (.A0(\phase_increment[0] [5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17510), .COUT(n17511), .S0(phase_increment_1__63__N_17[5]), 
          .S1(phase_increment_1__63__N_17[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_3.INIT0 = 16'h555f;
    defparam _add_1_3591_add_4_3.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3567_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5327), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16690));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3567_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3567_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3567_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3567_add_4_1.INJECT1_1 = "NO";
    LUT4 mux_1352_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n2541), 
         .Z(n2566)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1352_i1_3_lut_3_lut.init = 16'hd1d1;
    PFUMX mux_1706_i1 (.BLUT(n3026), .ALUT(n3036), .C0(led_0_6), .Z(n3042));
    LUT4 mux_1457_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n2682), 
         .Z(n2707)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1457_i1_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_2577_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n4186), 
         .Z(n4211)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2577_i1_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i5018_2_lut (.A(phase_increment_1__63__N_17[7]), .B(led_0_6), .Z(n4050)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i5018_2_lut.init = 16'heeee;
    PFUMX mux_1949_i1 (.BLUT(n3360), .ALUT(n3345), .C0(rx_byte[2]), .Z(n3368));
    CCU2C _add_1_3534_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16686), .S0(cout_adj_5269));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_3534_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_3534_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_cout.INJECT1_1 = "NO";
    PFUMX mux_1286_i1 (.BLUT(n2462), .ALUT(n2472), .C0(led_0_6), .Z(n2478));
    PFUMX mux_2334_i1 (.BLUT(n3877), .ALUT(n3862), .C0(rx_byte[2]), .Z(n3885));
    CCU2C _add_1_3534_add_4_36 (.A0(integrator2_adj_6559[34]), .B0(integrator1_adj_6558[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[35]), .B1(integrator1_adj_6558[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16685), .COUT(n16686), .S0(integrator2_71__N_1032_adj_6574[34]), 
          .S1(integrator2_71__N_1032_adj_6574[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_34 (.A0(integrator2_adj_6559[32]), .B0(integrator1_adj_6558[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[33]), .B1(integrator1_adj_6558[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16684), .COUT(n16685), .S0(integrator2_71__N_1032_adj_6574[32]), 
          .S1(integrator2_71__N_1032_adj_6574[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_34.INJECT1_1 = "NO";
    FD1S3AX _add_1_3507_i7 (.D(cout_adj_5314), .CK(clk_80mhz), .Q(pwm_out_c));
    defparam _add_1_3507_i7.GSR = "ENABLED";
    CCU2C _add_1_3798_add_4_6 (.A0(integrator3[39]), .B0(integrator2[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[40]), .B1(integrator2[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17717), .COUT(n17718), .S0(n174_adj_6277), 
          .S1(n171_adj_6276));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3798_add_4_4 (.A0(integrator3[37]), .B0(integrator2[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[38]), .B1(integrator2[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17716), .COUT(n17717), .S0(n180_adj_6279), 
          .S1(n177_adj_6278));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3798_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_32 (.A0(integrator2_adj_6559[30]), .B0(integrator1_adj_6558[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[31]), .B1(integrator1_adj_6558[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16683), .COUT(n16684), .S0(integrator2_71__N_1032_adj_6574[30]), 
          .S1(integrator2_71__N_1032_adj_6574[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3798_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator3[36]), .B1(integrator2[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17716), .S1(n183_adj_6280));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3798_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3798_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3798_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3798_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3591_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\phase_increment[0] [4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17510), .S1(phase_increment_1__63__N_17[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(283[40:79])
    defparam _add_1_3591_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3591_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3591_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3591_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_38 (.A0(comb_d9_adj_6570[35]), .B0(comb9_adj_6569[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17715), .S1(cout_adj_6281));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3801_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_36 (.A0(comb_d9_adj_6570[33]), .B0(comb9_adj_6569[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[34]), .B1(comb9_adj_6569[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17714), .COUT(n17715));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_36.INJECT1_1 = "NO";
    LUT4 mux_1939_i1_3_lut (.A(phase_increment_1__63__N_19[22]), .B(phase_increment_1__63__N_20[22]), 
         .C(rx_byte[0]), .Z(n3355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1939_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3801_add_4_34 (.A0(comb_d9_adj_6570[31]), .B0(comb9_adj_6569[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[32]), .B1(comb9_adj_6569[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17713), .COUT(n17714));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_32 (.A0(comb_d9_adj_6570[29]), .B0(comb9_adj_6569[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[30]), .B1(comb9_adj_6569[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17712), .COUT(n17713));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_30 (.A0(integrator2_adj_6559[28]), .B0(integrator1_adj_6558[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[29]), .B1(integrator1_adj_6558[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16682), .COUT(n16683), .S0(integrator2_71__N_1032_adj_6574[28]), 
          .S1(integrator2_71__N_1032_adj_6574[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_30.INJECT1_1 = "NO";
    LUT4 i4891_2_lut (.A(phase_increment_1__63__N_21[55]), .B(rx_byte[0]), 
         .Z(n1809)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4891_2_lut.init = 16'heeee;
    CCU2C _add_1_3594_add_4_13 (.A0(sine_table_value[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17509), .S0(n28_adj_6326));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[48:65])
    defparam _add_1_3594_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_3594_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_3594_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3594_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3645_add_4_21 (.A0(integrator_tmp_adj_6556[54]), .B0(cout_adj_6512), 
          .C0(n129_adj_5778), .D0(n19_adj_5473), .A1(integrator_tmp_adj_6556[55]), 
          .B1(cout_adj_6512), .C1(n126_adj_5777), .D1(n18_adj_5472), .CIN(n17243), 
          .COUT(n17244), .S0(comb6_71__N_1993_adj_6589[54]), .S1(comb6_71__N_1993_adj_6589[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_28 (.A0(integrator2_adj_6559[26]), .B0(integrator1_adj_6558[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[27]), .B1(integrator1_adj_6558[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16681), .COUT(n16682), .S0(integrator2_71__N_1032_adj_6574[26]), 
          .S1(integrator2_71__N_1032_adj_6574[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3645_add_4_19 (.A0(integrator_tmp_adj_6556[52]), .B0(cout_adj_6512), 
          .C0(n135_adj_5780), .D0(n21_adj_5475), .A1(integrator_tmp_adj_6556[53]), 
          .B1(cout_adj_6512), .C1(n132_adj_5779), .D1(n20_adj_5474), .CIN(n17242), 
          .COUT(n17243), .S0(comb6_71__N_1993_adj_6589[52]), .S1(comb6_71__N_1993_adj_6589[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_19.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_5__bdd_4_lut (.A(phase_increment_1__63__N_21[5]), 
         .B(rx_byte[0]), .C(n19426), .D(rx_byte[2]), .Z(n19806)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam phase_increment_1__63__N_21_5__bdd_4_lut.init = 16'hf0ee;
    LUT4 mux_1492_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n2729), 
         .Z(n2754)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1492_i1_3_lut_3_lut.init = 16'hd1d1;
    CCU2C _add_1_3645_add_4_17 (.A0(integrator_tmp_adj_6556[50]), .B0(cout_adj_6512), 
          .C0(n141_adj_5782), .D0(n23_adj_5477), .A1(integrator_tmp_adj_6556[51]), 
          .B1(cout_adj_6512), .C1(n138_adj_5781), .D1(n22_adj_5476), .CIN(n17241), 
          .COUT(n17242), .S0(comb6_71__N_1993_adj_6589[50]), .S1(comb6_71__N_1993_adj_6589[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3645_add_4_15 (.A0(integrator_tmp_adj_6556[48]), .B0(cout_adj_6512), 
          .C0(n147_adj_5784), .D0(n25_adj_5479), .A1(integrator_tmp_adj_6556[49]), 
          .B1(cout_adj_6512), .C1(n144_adj_5783), .D1(n24_adj_5478), .CIN(n17240), 
          .COUT(n17241), .S0(comb6_71__N_1993_adj_6589[48]), .S1(comb6_71__N_1993_adj_6589[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3645_add_4_13 (.A0(integrator_tmp_adj_6556[46]), .B0(cout_adj_6512), 
          .C0(n153_adj_5786), .D0(n27_adj_5481), .A1(integrator_tmp_adj_6556[47]), 
          .B1(cout_adj_6512), .C1(n150_adj_5785), .D1(n26_adj_5480), .CIN(n17239), 
          .COUT(n17240), .S0(comb6_71__N_1993_adj_6589[46]), .S1(comb6_71__N_1993_adj_6589[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_30 (.A0(comb_d9_adj_6570[27]), .B0(comb9_adj_6569[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[28]), .B1(comb9_adj_6569[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17711), .COUT(n17712));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3594_add_4_11 (.A0(sine_table_value[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(sine_table_value[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17508), .COUT(n17509), .S0(n34_adj_6328), 
          .S1(n31_adj_6327));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[48:65])
    defparam _add_1_3594_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_3594_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_3594_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3594_add_4_11.INJECT1_1 = "NO";
    LUT4 n1836_bdd_3_lut (.A(phase_increment_1__63__N_19[54]), .B(phase_increment_1__63__N_20[54]), 
         .C(rx_byte[0]), .Z(n19423)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1836_bdd_3_lut.init = 16'hcaca;
    CCU2C _add_1_3801_add_4_28 (.A0(comb_d9_adj_6570[25]), .B0(comb9_adj_6569[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[26]), .B1(comb9_adj_6569[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17710), .COUT(n17711));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_26 (.A0(comb_d9_adj_6570[23]), .B0(comb9_adj_6569[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[24]), .B1(comb9_adj_6569[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17709), .COUT(n17710));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3645_add_4_11 (.A0(integrator_tmp_adj_6556[44]), .B0(cout_adj_6512), 
          .C0(n159_adj_5788), .D0(n29_adj_5483), .A1(integrator_tmp_adj_6556[45]), 
          .B1(cout_adj_6512), .C1(n156_adj_5787), .D1(n28_adj_5482), .CIN(n17238), 
          .COUT(n17239), .S0(comb6_71__N_1993_adj_6589[44]), .S1(comb6_71__N_1993_adj_6589[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3594_add_4_9 (.A0(sine_table_value[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(sine_table_value[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17507), .COUT(n17508), .S0(n40_adj_6330), 
          .S1(n37_adj_6329));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[48:65])
    defparam _add_1_3594_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_3594_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_3594_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3594_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3645_add_4_9 (.A0(integrator_tmp_adj_6556[42]), .B0(cout_adj_6512), 
          .C0(n165_adj_5790), .D0(n31_adj_5485), .A1(integrator_tmp_adj_6556[43]), 
          .B1(cout_adj_6512), .C1(n162_adj_5789), .D1(n30_adj_5484), .CIN(n17237), 
          .COUT(n17238), .S0(comb6_71__N_1993_adj_6589[42]), .S1(comb6_71__N_1993_adj_6589[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3645_add_4_7 (.A0(integrator_tmp_adj_6556[40]), .B0(cout_adj_6512), 
          .C0(n171_adj_5792), .D0(n33_adj_5487), .A1(integrator_tmp_adj_6556[41]), 
          .B1(cout_adj_6512), .C1(n168_adj_5791), .D1(n32_adj_5486), .CIN(n17236), 
          .COUT(n17237), .S0(comb6_71__N_1993_adj_6589[40]), .S1(comb6_71__N_1993_adj_6589[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_7.INJECT1_1 = "NO";
    LUT4 mux_2417_i1_3_lut (.A(phase_increment_1__63__N_16[8]), .B(phase_increment_1__63__N_18[8]), 
         .C(rx_byte[0]), .Z(n3998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2417_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1632_i1_3_lut_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n2917), 
         .Z(n2942)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1632_i1_3_lut_3_lut.init = 16'hd1d1;
    CCU2C _add_1_3645_add_4_5 (.A0(integrator_tmp_adj_6556[38]), .B0(cout_adj_6512), 
          .C0(n177_adj_5794), .D0(n35_adj_5489), .A1(integrator_tmp_adj_6556[39]), 
          .B1(cout_adj_6512), .C1(n174_adj_5793), .D1(n34_adj_5488), .CIN(n17235), 
          .COUT(n17236), .S0(comb6_71__N_1993_adj_6589[38]), .S1(comb6_71__N_1993_adj_6589[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_5.INJECT1_1 = "NO";
    PFUMX i8437 (.BLUT(n19417), .ALUT(n19416), .C0(rx_byte[2]), .Z(n19418));
    CCU2C _add_1_3645_add_4_3 (.A0(integrator_tmp_adj_6556[36]), .B0(cout_adj_6512), 
          .C0(n183_adj_5796), .D0(n37_adj_5491), .A1(integrator_tmp_adj_6556[37]), 
          .B1(cout_adj_6512), .C1(n180_adj_5795), .D1(n36_adj_5490), .CIN(n17234), 
          .COUT(n17235), .S0(comb6_71__N_1993_adj_6589[36]), .S1(comb6_71__N_1993_adj_6589[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3645_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3645_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3645_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_6512), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17234));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3645_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3645_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3645_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3645_add_4_1.INJECT1_1 = "NO";
    LUT4 n1424_bdd_3_lut_8475_3_lut (.A(rx_byte[2]), .B(rx_byte[3]), .C(n19432), 
         .Z(n19433)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam n1424_bdd_3_lut_8475_3_lut.init = 16'hd1d1;
    CCU2C _add_1_3594_add_4_7 (.A0(sine_table_value[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(sine_table_value[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17506), .COUT(n17507), .S0(n46_adj_6332), 
          .S1(n43_adj_6331));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[48:65])
    defparam _add_1_3594_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_3594_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_3594_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3594_add_4_7.INJECT1_1 = "NO";
    LUT4 mux_842_i1_3_lut (.A(phase_increment_1__63__N_16[53]), .B(phase_increment_1__63__N_18[53]), 
         .C(rx_byte[0]), .Z(n1883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_842_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3801_add_4_24 (.A0(comb_d9_adj_6570[21]), .B0(comb9_adj_6569[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[22]), .B1(comb9_adj_6569[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17708), .COUT(n17709));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_37 (.A0(comb6_adj_6563[70]), .B0(cout_adj_5627), 
          .C0(n81_adj_5726), .D0(n3_adj_5493), .A1(comb6_adj_6563[71]), 
          .B1(cout_adj_5627), .C1(n78_adj_5725), .D1(n2_adj_5492), .CIN(n17229), 
          .S0(comb7_71__N_2065_adj_6590[70]), .S1(comb7_71__N_2065_adj_6590[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_37.INJECT1_1 = "NO";
    LUT4 i4995_2_lut (.A(phase_increment_1__63__N_21[15]), .B(rx_byte[0]), 
         .Z(n3689)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4995_2_lut.init = 16'heeee;
    LUT4 i4905_2_lut (.A(phase_increment_1__63__N_17[56]), .B(led_0_6), 
         .Z(n1747)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4905_2_lut.init = 16'heeee;
    CCU2C _add_1_3594_add_4_5 (.A0(sine_table_value[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(sine_table_value[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17505), .COUT(n17506), .S0(n52_adj_6334), 
          .S1(n49_adj_6333));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[48:65])
    defparam _add_1_3594_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_3594_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_3594_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3594_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_35 (.A0(comb6_adj_6563[68]), .B0(cout_adj_5627), 
          .C0(n87_adj_5728), .D0(n5_adj_5495), .A1(comb6_adj_6563[69]), 
          .B1(cout_adj_5627), .C1(n84_adj_5727), .D1(n4_adj_5494), .CIN(n17228), 
          .COUT(n17229), .S0(comb7_71__N_2065_adj_6590[68]), .S1(comb7_71__N_2065_adj_6590[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_35.INJECT1_1 = "NO";
    LUT4 n2776_bdd_3_lut_8595 (.A(n2776), .B(rx_byte[2]), .C(rx_byte[3]), 
         .Z(n19627)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n2776_bdd_3_lut_8595.init = 16'hacac;
    CCU2C _add_1_3801_add_4_22 (.A0(comb_d9_adj_6570[19]), .B0(comb9_adj_6569[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[20]), .B1(comb9_adj_6569[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17707), .COUT(n17708));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_33 (.A0(comb6_adj_6563[66]), .B0(cout_adj_5627), 
          .C0(n93_adj_5730), .D0(n7_adj_5497), .A1(comb6_adj_6563[67]), 
          .B1(cout_adj_5627), .C1(n90_adj_5729), .D1(n6_adj_5496), .CIN(n17227), 
          .COUT(n17228), .S0(comb7_71__N_2065_adj_6590[66]), .S1(comb7_71__N_2065_adj_6590[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3594_add_4_3 (.A0(sine_table_value[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(sine_table_value[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17504), .COUT(n17505), .S0(n58_adj_6336), 
          .S1(n55_adj_6335));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[48:65])
    defparam _add_1_3594_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_3594_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_3594_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3594_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_31 (.A0(comb6_adj_6563[64]), .B0(cout_adj_5627), 
          .C0(n99_adj_5732), .D0(n9_adj_5499), .A1(comb6_adj_6563[65]), 
          .B1(cout_adj_5627), .C1(n96_adj_5731), .D1(n8_adj_5498), .CIN(n17226), 
          .COUT(n17227), .S0(comb7_71__N_2065_adj_6590[64]), .S1(comb7_71__N_2065_adj_6590[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_31.INJECT1_1 = "NO";
    PFUMX mux_1179_i1 (.BLUT(n2326), .ALUT(n2311), .C0(rx_byte[2]), .Z(n2334));
    CCU2C _add_1_3648_add_4_29 (.A0(comb6_adj_6563[62]), .B0(cout_adj_5627), 
          .C0(n105_adj_5734), .D0(n11_adj_5501), .A1(comb6_adj_6563[63]), 
          .B1(cout_adj_5627), .C1(n102_adj_5733), .D1(n10_adj_5500), .CIN(n17225), 
          .COUT(n17226), .S0(comb7_71__N_2065_adj_6590[62]), .S1(comb7_71__N_2065_adj_6590[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_27 (.A0(comb6_adj_6563[60]), .B0(cout_adj_5627), 
          .C0(n111_adj_5736), .D0(n13_adj_5503), .A1(comb6_adj_6563[61]), 
          .B1(cout_adj_5627), .C1(n108_adj_5735), .D1(n12_adj_5502), .CIN(n17224), 
          .COUT(n17225), .S0(comb7_71__N_2065_adj_6590[60]), .S1(comb7_71__N_2065_adj_6590[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_25 (.A0(comb6_adj_6563[58]), .B0(cout_adj_5627), 
          .C0(n117_adj_5738), .D0(n15_adj_5505), .A1(comb6_adj_6563[59]), 
          .B1(cout_adj_5627), .C1(n114_adj_5737), .D1(n14_adj_5504), .CIN(n17223), 
          .COUT(n17224), .S0(comb7_71__N_2065_adj_6590[58]), .S1(comb7_71__N_2065_adj_6590[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_23 (.A0(comb6_adj_6563[56]), .B0(cout_adj_5627), 
          .C0(n123_adj_5740), .D0(n17_adj_5507), .A1(comb6_adj_6563[57]), 
          .B1(cout_adj_5627), .C1(n120_adj_5739), .D1(n16_adj_5506), .CIN(n17222), 
          .COUT(n17223), .S0(comb7_71__N_2065_adj_6590[56]), .S1(comb7_71__N_2065_adj_6590[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_23.INJECT1_1 = "NO";
    LUT4 n2776_bdd_3_lut (.A(phase_increment_1__63__N_19[34]), .B(phase_increment_1__63__N_20[34]), 
         .C(rx_byte[0]), .Z(n19628)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n2776_bdd_3_lut.init = 16'hcaca;
    CCU2C _add_1_3648_add_4_21 (.A0(comb6_adj_6563[54]), .B0(cout_adj_5627), 
          .C0(n129_adj_5742), .D0(n19_adj_5509), .A1(comb6_adj_6563[55]), 
          .B1(cout_adj_5627), .C1(n126_adj_5741), .D1(n18_adj_5508), .CIN(n17221), 
          .COUT(n17222), .S0(comb7_71__N_2065_adj_6590[54]), .S1(comb7_71__N_2065_adj_6590[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_19 (.A0(comb6_adj_6563[52]), .B0(cout_adj_5627), 
          .C0(n135_adj_5744), .D0(n21_adj_5511), .A1(comb6_adj_6563[53]), 
          .B1(cout_adj_5627), .C1(n132_adj_5743), .D1(n20_adj_5510), .CIN(n17220), 
          .COUT(n17221), .S0(comb7_71__N_2065_adj_6590[52]), .S1(comb7_71__N_2065_adj_6590[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_17 (.A0(comb6_adj_6563[50]), .B0(cout_adj_5627), 
          .C0(n141_adj_5746), .D0(n23_adj_5513), .A1(comb6_adj_6563[51]), 
          .B1(cout_adj_5627), .C1(n138_adj_5745), .D1(n22_adj_5512), .CIN(n17219), 
          .COUT(n17220), .S0(comb7_71__N_2065_adj_6590[50]), .S1(comb7_71__N_2065_adj_6590[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_17.INJECT1_1 = "NO";
    L6MUX21 i8740 (.D0(n19797), .D1(n19794), .SD(n19822), .Z(n19798));
    LUT4 phase_increment_1__63__N_21_8__bdd_2_lut_8699 (.A(phase_increment_1__63__N_21[8]), 
         .B(rx_byte[0]), .Z(n19441)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_8__bdd_2_lut_8699.init = 16'heeee;
    CCU2C _add_1_3534_add_4_26 (.A0(integrator2_adj_6559[24]), .B0(integrator1_adj_6558[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[25]), .B1(integrator1_adj_6558[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16680), .COUT(n16681), .S0(integrator2_71__N_1032_adj_6574[24]), 
          .S1(integrator2_71__N_1032_adj_6574[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_15 (.A0(comb6_adj_6563[48]), .B0(cout_adj_5627), 
          .C0(n147_adj_5748), .D0(n25_adj_5515), .A1(comb6_adj_6563[49]), 
          .B1(cout_adj_5627), .C1(n144_adj_5747), .D1(n24_adj_5514), .CIN(n17218), 
          .COUT(n17219), .S0(comb7_71__N_2065_adj_6590[48]), .S1(comb7_71__N_2065_adj_6590[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_15.INJECT1_1 = "NO";
    PFUMX i8738 (.BLUT(n19796), .ALUT(n19795), .C0(led_0_6), .Z(n19797));
    CCU2C _add_1_3648_add_4_13 (.A0(comb6_adj_6563[46]), .B0(cout_adj_5627), 
          .C0(n153_adj_5750), .D0(n27_adj_5517), .A1(comb6_adj_6563[47]), 
          .B1(cout_adj_5627), .C1(n150_adj_5749), .D1(n26_adj_5516), .CIN(n17217), 
          .COUT(n17218), .S0(comb7_71__N_2065_adj_6590[46]), .S1(comb7_71__N_2065_adj_6590[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3594_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(sine_table_value[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17504), .S1(n61_adj_6337));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[48:65])
    defparam _add_1_3594_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3594_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_3594_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3594_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_24 (.A0(integrator2_adj_6559[22]), .B0(integrator1_adj_6558[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[23]), .B1(integrator1_adj_6558[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16679), .COUT(n16680), .S0(integrator2_71__N_1032_adj_6574[22]), 
          .S1(integrator2_71__N_1032_adj_6574[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_11 (.A0(comb6_adj_6563[44]), .B0(cout_adj_5627), 
          .C0(n159_adj_5752), .D0(n29_adj_5519), .A1(comb6_adj_6563[45]), 
          .B1(cout_adj_5627), .C1(n156_adj_5751), .D1(n28_adj_5518), .CIN(n17216), 
          .COUT(n17217), .S0(comb7_71__N_2065_adj_6590[44]), .S1(comb7_71__N_2065_adj_6590[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_11.INJECT1_1 = "NO";
    LUT4 i5019_2_lut (.A(phase_increment_1__63__N_21[7]), .B(rx_byte[0]), 
         .Z(n4065)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i5019_2_lut.init = 16'heeee;
    CCU2C _add_1_3534_add_4_22 (.A0(integrator2_adj_6559[20]), .B0(integrator1_adj_6558[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[21]), .B1(integrator1_adj_6558[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16678), .COUT(n16679), .S0(integrator2_71__N_1032_adj_6574[20]), 
          .S1(integrator2_71__N_1032_adj_6574[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_20 (.A0(integrator2_adj_6559[18]), .B0(integrator1_adj_6558[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[19]), .B1(integrator1_adj_6558[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16677), .COUT(n16678), .S0(integrator2_71__N_1032_adj_6574[18]), 
          .S1(integrator2_71__N_1032_adj_6574[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_20.INJECT1_1 = "NO";
    OB pwm_out_p_pad_2 (.I(pwm_out_p_c), .O(pwm_out_p[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(43[22:31])
    CCU2C _add_1_3534_add_4_18 (.A0(integrator2_adj_6559[16]), .B0(integrator1_adj_6558[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[17]), .B1(integrator1_adj_6558[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16676), .COUT(n16677), .S0(integrator2_71__N_1032_adj_6574[16]), 
          .S1(integrator2_71__N_1032_adj_6574[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_18.INJECT1_1 = "NO";
    OB diff_out_pad (.I(diff_out_c), .O(diff_out));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(41[22:30])
    CCU2C _add_1_3534_add_4_16 (.A0(integrator2_adj_6559[14]), .B0(integrator1_adj_6558[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[15]), .B1(integrator1_adj_6558[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16675), .COUT(n16676), .S0(integrator2_71__N_1032_adj_6574[14]), 
          .S1(integrator2_71__N_1032_adj_6574[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_14 (.A0(integrator2_adj_6559[12]), .B0(integrator1_adj_6558[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[13]), .B1(integrator1_adj_6558[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16674), .COUT(n16675), .S0(integrator2_71__N_1032_adj_6574[12]), 
          .S1(integrator2_71__N_1032_adj_6574[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_12 (.A0(integrator2_adj_6559[10]), .B0(integrator1_adj_6558[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[11]), .B1(integrator1_adj_6558[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16673), .COUT(n16674), .S0(integrator2_71__N_1032_adj_6574[10]), 
          .S1(integrator2_71__N_1032_adj_6574[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_10 (.A0(integrator2_adj_6559[8]), .B0(integrator1_adj_6558[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[9]), .B1(integrator1_adj_6558[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16672), .COUT(n16673), .S0(integrator2_71__N_1032_adj_6574[8]), 
          .S1(integrator2_71__N_1032_adj_6574[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_8 (.A0(integrator2_adj_6559[6]), .B0(integrator1_adj_6558[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[7]), .B1(integrator1_adj_6558[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16671), .COUT(n16672), .S0(integrator2_71__N_1032_adj_6574[6]), 
          .S1(integrator2_71__N_1032_adj_6574[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_6 (.A0(integrator2_adj_6559[4]), .B0(integrator1_adj_6558[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[5]), .B1(integrator1_adj_6558[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16670), .COUT(n16671), .S0(integrator2_71__N_1032_adj_6574[4]), 
          .S1(integrator2_71__N_1032_adj_6574[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_4 (.A0(integrator2_adj_6559[2]), .B0(integrator1_adj_6558[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[3]), .B1(integrator1_adj_6558[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16669), .COUT(n16670), .S0(integrator2_71__N_1032_adj_6574[2]), 
          .S1(integrator2_71__N_1032_adj_6574[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3534_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3534_add_4_2 (.A0(integrator2_adj_6559[0]), .B0(integrator1_adj_6558[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6559[1]), .B1(integrator1_adj_6558[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16669), .S1(integrator2_71__N_1032_adj_6574[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3534_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_3534_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3534_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3534_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_38 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16667), .S0(n78_adj_5268));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3570_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_36 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16666), .COUT(n16667), .S0(n84_adj_5266), 
          .S1(n81_adj_5267));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_34 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16665), .COUT(n16666), .S0(n90_adj_5264), 
          .S1(n87_adj_5265));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_32 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16664), .COUT(n16665), .S0(n96), 
          .S1(n93));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_30 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16663), .COUT(n16664), .S0(n102), 
          .S1(n99));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_28 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16662), .COUT(n16663), .S0(n108), 
          .S1(n105));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_26 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16661), .COUT(n16662), .S0(n114), 
          .S1(n111));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_24 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16660), .COUT(n16661), .S0(n120), 
          .S1(n117));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_22 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16659), .COUT(n16660), .S0(n126), 
          .S1(n123));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_20 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16658), .COUT(n16659), .S0(n132), 
          .S1(n129));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_18 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16657), .COUT(n16658), .S0(n138), 
          .S1(n135));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_16 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16656), .COUT(n16657), .S0(n144), 
          .S1(n141_adj_4975));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_14 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16655), .COUT(n16656), .S0(n150), 
          .S1(n147));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_12 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16654), .COUT(n16655), .S0(n156), 
          .S1(n153));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_10 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16653), .COUT(n16654), .S0(n162), 
          .S1(n159));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_8 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16652), .COUT(n16653), .S0(n168), 
          .S1(n165));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_6 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16651), .COUT(n16652), .S0(n174), 
          .S1(n171));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_4 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16650), .COUT(n16651), .S0(n180), 
          .S1(n177));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3570_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3570_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16650), .S1(n183));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3570_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3570_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3570_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3570_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3507_add_4_12 (.A0(count_adj_6635[9]), .B0(data_in_reg[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16649), .S1(cout_adj_5314));
    defparam _add_1_3507_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3507_add_4_12.INIT1 = 16'h0000;
    defparam _add_1_3507_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3507_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3507_add_4_10 (.A0(count_adj_6635[7]), .B0(data_in_reg[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(count_adj_6635[8]), .B1(data_in_reg[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16648), .COUT(n16649));
    defparam _add_1_3507_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3507_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3507_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3507_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3507_add_4_8 (.A0(count_adj_6635[5]), .B0(data_in_reg[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(count_adj_6635[6]), .B1(data_in_reg[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16647), .COUT(n16648));
    defparam _add_1_3507_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3507_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3507_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3507_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3507_add_4_6 (.A0(count_adj_6635[3]), .B0(data_in_reg[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(count_adj_6635[4]), .B1(data_in_reg[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16646), .COUT(n16647));
    defparam _add_1_3507_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3507_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3507_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3507_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3507_add_4_4 (.A0(count_adj_6635[1]), .B0(data_in_reg[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(count_adj_6635[2]), .B1(data_in_reg[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16645), .COUT(n16646));
    defparam _add_1_3507_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3507_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3507_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3507_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3507_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_6635[0]), .B1(data_in_reg[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16645));
    defparam _add_1_3507_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3507_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3507_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3507_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16644), .S0(cout));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_3537_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_3537_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_36 (.A0(integrator3_adj_6560[34]), .B0(integrator2_adj_6559[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[35]), .B1(integrator2_adj_6559[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16643), .COUT(n16644), .S0(integrator3_71__N_1104_adj_6575[34]), 
          .S1(integrator3_71__N_1104_adj_6575[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_34 (.A0(integrator3_adj_6560[32]), .B0(integrator2_adj_6559[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[33]), .B1(integrator2_adj_6559[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16642), .COUT(n16643), .S0(integrator3_71__N_1104_adj_6575[32]), 
          .S1(integrator3_71__N_1104_adj_6575[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_32 (.A0(integrator3_adj_6560[30]), .B0(integrator2_adj_6559[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[31]), .B1(integrator2_adj_6559[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16641), .COUT(n16642), .S0(integrator3_71__N_1104_adj_6575[30]), 
          .S1(integrator3_71__N_1104_adj_6575[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_30 (.A0(integrator3_adj_6560[28]), .B0(integrator2_adj_6559[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[29]), .B1(integrator2_adj_6559[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16640), .COUT(n16641), .S0(integrator3_71__N_1104_adj_6575[28]), 
          .S1(integrator3_71__N_1104_adj_6575[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_28 (.A0(integrator3_adj_6560[26]), .B0(integrator2_adj_6559[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[27]), .B1(integrator2_adj_6559[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16639), .COUT(n16640), .S0(integrator3_71__N_1104_adj_6575[26]), 
          .S1(integrator3_71__N_1104_adj_6575[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_26 (.A0(integrator3_adj_6560[24]), .B0(integrator2_adj_6559[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[25]), .B1(integrator2_adj_6559[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16638), .COUT(n16639), .S0(integrator3_71__N_1104_adj_6575[24]), 
          .S1(integrator3_71__N_1104_adj_6575[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_24 (.A0(integrator3_adj_6560[22]), .B0(integrator2_adj_6559[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[23]), .B1(integrator2_adj_6559[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16637), .COUT(n16638), .S0(integrator3_71__N_1104_adj_6575[22]), 
          .S1(integrator3_71__N_1104_adj_6575[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_22 (.A0(integrator3_adj_6560[20]), .B0(integrator2_adj_6559[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[21]), .B1(integrator2_adj_6559[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16636), .COUT(n16637), .S0(integrator3_71__N_1104_adj_6575[20]), 
          .S1(integrator3_71__N_1104_adj_6575[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_20 (.A0(integrator3_adj_6560[18]), .B0(integrator2_adj_6559[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[19]), .B1(integrator2_adj_6559[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16635), .COUT(n16636), .S0(integrator3_71__N_1104_adj_6575[18]), 
          .S1(integrator3_71__N_1104_adj_6575[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_18 (.A0(integrator3_adj_6560[16]), .B0(integrator2_adj_6559[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[17]), .B1(integrator2_adj_6559[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16634), .COUT(n16635), .S0(integrator3_71__N_1104_adj_6575[16]), 
          .S1(integrator3_71__N_1104_adj_6575[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_16 (.A0(integrator3_adj_6560[14]), .B0(integrator2_adj_6559[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[15]), .B1(integrator2_adj_6559[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16633), .COUT(n16634), .S0(integrator3_71__N_1104_adj_6575[14]), 
          .S1(integrator3_71__N_1104_adj_6575[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_14 (.A0(integrator3_adj_6560[12]), .B0(integrator2_adj_6559[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[13]), .B1(integrator2_adj_6559[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16632), .COUT(n16633), .S0(integrator3_71__N_1104_adj_6575[12]), 
          .S1(integrator3_71__N_1104_adj_6575[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_12 (.A0(integrator3_adj_6560[10]), .B0(integrator2_adj_6559[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[11]), .B1(integrator2_adj_6559[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16631), .COUT(n16632), .S0(integrator3_71__N_1104_adj_6575[10]), 
          .S1(integrator3_71__N_1104_adj_6575[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_10 (.A0(integrator3_adj_6560[8]), .B0(integrator2_adj_6559[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[9]), .B1(integrator2_adj_6559[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16630), .COUT(n16631), .S0(integrator3_71__N_1104_adj_6575[8]), 
          .S1(integrator3_71__N_1104_adj_6575[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_8 (.A0(integrator3_adj_6560[6]), .B0(integrator2_adj_6559[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[7]), .B1(integrator2_adj_6559[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16629), .COUT(n16630), .S0(integrator3_71__N_1104_adj_6575[6]), 
          .S1(integrator3_71__N_1104_adj_6575[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_6 (.A0(integrator3_adj_6560[4]), .B0(integrator2_adj_6559[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[5]), .B1(integrator2_adj_6559[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16628), .COUT(n16629), .S0(integrator3_71__N_1104_adj_6575[4]), 
          .S1(integrator3_71__N_1104_adj_6575[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_4 (.A0(integrator3_adj_6560[2]), .B0(integrator2_adj_6559[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[3]), .B1(integrator2_adj_6559[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16627), .COUT(n16628), .S0(integrator3_71__N_1104_adj_6575[2]), 
          .S1(integrator3_71__N_1104_adj_6575[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3537_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3537_add_4_2 (.A0(integrator3_adj_6560[0]), .B0(integrator2_adj_6559[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[1]), .B1(integrator2_adj_6559[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16627), .S1(integrator3_71__N_1104_adj_6575[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3537_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_3537_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3537_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3537_add_4_2.INJECT1_1 = "NO";
    PFUMX i8735 (.BLUT(n19793), .ALUT(n19792), .C0(rx_byte[2]), .Z(n19794));
    CCU2C _add_1_3717_add_4_38 (.A0(comb_d7[71]), .B0(comb7[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16625), .S0(n78_adj_5892));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3717_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_36 (.A0(comb_d7[69]), .B0(comb7[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[70]), .B1(comb7[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16624), .COUT(n16625), .S0(n84_adj_5894), 
          .S1(n81_adj_5893));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_34 (.A0(comb_d7[67]), .B0(comb7[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[68]), .B1(comb7[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16623), .COUT(n16624), .S0(n90_adj_5896), 
          .S1(n87_adj_5895));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_32 (.A0(comb_d7[65]), .B0(comb7[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[66]), .B1(comb7[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16622), .COUT(n16623), .S0(n96_adj_5898), 
          .S1(n93_adj_5897));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_30 (.A0(comb_d7[63]), .B0(comb7[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[64]), .B1(comb7[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16621), .COUT(n16622), .S0(n102_adj_5900), 
          .S1(n99_adj_5899));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_28 (.A0(comb_d7[61]), .B0(comb7[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[62]), .B1(comb7[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16620), .COUT(n16621), .S0(n108_adj_5902), 
          .S1(n105_adj_5901));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_26 (.A0(comb_d7[59]), .B0(comb7[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[60]), .B1(comb7[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16619), .COUT(n16620), .S0(n114_adj_5904), 
          .S1(n111_adj_5903));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_24 (.A0(comb_d7[57]), .B0(comb7[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[58]), .B1(comb7[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16618), .COUT(n16619), .S0(n120_adj_5906), 
          .S1(n117_adj_5905));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_22 (.A0(comb_d7[55]), .B0(comb7[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[56]), .B1(comb7[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16617), .COUT(n16618), .S0(n126_adj_5908), 
          .S1(n123_adj_5907));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_20 (.A0(comb_d7[53]), .B0(comb7[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[54]), .B1(comb7[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16616), .COUT(n16617), .S0(n132_adj_5910), 
          .S1(n129_adj_5909));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_18 (.A0(comb_d7[51]), .B0(comb7[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[52]), .B1(comb7[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16615), .COUT(n16616), .S0(n138_adj_5912), 
          .S1(n135_adj_5911));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_16 (.A0(comb_d7[49]), .B0(comb7[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[50]), .B1(comb7[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16614), .COUT(n16615), .S0(n144_adj_5914), 
          .S1(n141_adj_5913));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_14 (.A0(comb_d7[47]), .B0(comb7[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[48]), .B1(comb7[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16613), .COUT(n16614), .S0(n150_adj_5916), 
          .S1(n147_adj_5915));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_12 (.A0(comb_d7[45]), .B0(comb7[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[46]), .B1(comb7[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16612), .COUT(n16613), .S0(n156_adj_5918), 
          .S1(n153_adj_5917));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_10 (.A0(comb_d7[43]), .B0(comb7[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[44]), .B1(comb7[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16611), .COUT(n16612), .S0(n162_adj_5920), 
          .S1(n159_adj_5919));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_8 (.A0(comb_d7[41]), .B0(comb7[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[42]), .B1(comb7[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16610), .COUT(n16611), .S0(n168_adj_5922), 
          .S1(n165_adj_5921));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_6 (.A0(comb_d7[39]), .B0(comb7[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[40]), .B1(comb7[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16609), .COUT(n16610), .S0(n174_adj_5924), 
          .S1(n171_adj_5923));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_4 (.A0(comb_d7[37]), .B0(comb7[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[38]), .B1(comb7[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16608), .COUT(n16609), .S0(n180_adj_5926), 
          .S1(n177_adj_5925));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3717_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3717_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[36]), .B1(comb7[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16608), .S1(n183_adj_5927));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3717_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3717_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3717_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3717_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_38 (.A0(comb_d6[71]), .B0(comb6[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16607), .S0(n78_adj_5928));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3720_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_36 (.A0(comb_d6[69]), .B0(comb6[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[70]), .B1(comb6[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16606), .COUT(n16607), .S0(n84_adj_5930), 
          .S1(n81_adj_5929));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_34 (.A0(comb_d6[67]), .B0(comb6[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[68]), .B1(comb6[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16605), .COUT(n16606), .S0(n90_adj_5932), 
          .S1(n87_adj_5931));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_32 (.A0(comb_d6[65]), .B0(comb6[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[66]), .B1(comb6[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16604), .COUT(n16605), .S0(n96_adj_5934), 
          .S1(n93_adj_5933));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_30 (.A0(comb_d6[63]), .B0(comb6[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[64]), .B1(comb6[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16603), .COUT(n16604), .S0(n102_adj_5936), 
          .S1(n99_adj_5935));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_28 (.A0(comb_d6[61]), .B0(comb6[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[62]), .B1(comb6[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16602), .COUT(n16603), .S0(n108_adj_5938), 
          .S1(n105_adj_5937));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_26 (.A0(comb_d6[59]), .B0(comb6[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[60]), .B1(comb6[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16601), .COUT(n16602), .S0(n114_adj_5940), 
          .S1(n111_adj_5939));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_24 (.A0(comb_d6[57]), .B0(comb6[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[58]), .B1(comb6[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16600), .COUT(n16601), .S0(n120_adj_5942), 
          .S1(n117_adj_5941));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_22 (.A0(comb_d6[55]), .B0(comb6[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[56]), .B1(comb6[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16599), .COUT(n16600), .S0(n126_adj_5944), 
          .S1(n123_adj_5943));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_20 (.A0(comb_d6[53]), .B0(comb6[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[54]), .B1(comb6[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16598), .COUT(n16599), .S0(n132_adj_5946), 
          .S1(n129_adj_5945));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_18 (.A0(comb_d6[51]), .B0(comb6[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[52]), .B1(comb6[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16597), .COUT(n16598), .S0(n138_adj_5948), 
          .S1(n135_adj_5947));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_18.INJECT1_1 = "NO";
    L6MUX21 i8731 (.D0(n19790), .D1(n19787), .SD(n19822), .Z(n19791));
    PFUMX i8729 (.BLUT(n19789), .ALUT(n19788), .C0(led_0_6), .Z(n19790));
    PFUMX i8726 (.BLUT(n19786), .ALUT(n19785), .C0(rx_byte[2]), .Z(n19787));
    CCU2C _add_1_3720_add_4_16 (.A0(comb_d6[49]), .B0(comb6[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[50]), .B1(comb6[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16596), .COUT(n16597), .S0(n144_adj_5950), 
          .S1(n141_adj_5949));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_14 (.A0(comb_d6[47]), .B0(comb6[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[48]), .B1(comb6[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16595), .COUT(n16596), .S0(n150_adj_5952), 
          .S1(n147_adj_5951));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_12 (.A0(comb_d6[45]), .B0(comb6[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[46]), .B1(comb6[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16594), .COUT(n16595), .S0(n156_adj_5954), 
          .S1(n153_adj_5953));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_10 (.A0(comb_d6[43]), .B0(comb6[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[44]), .B1(comb6[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16593), .COUT(n16594), .S0(n162_adj_5956), 
          .S1(n159_adj_5955));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_8 (.A0(comb_d6[41]), .B0(comb6[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[42]), .B1(comb6[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16592), .COUT(n16593), .S0(n168_adj_5958), 
          .S1(n165_adj_5957));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_6 (.A0(comb_d6[39]), .B0(comb6[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[40]), .B1(comb6[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16591), .COUT(n16592), .S0(n174_adj_5960), 
          .S1(n171_adj_5959));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_4 (.A0(comb_d6[37]), .B0(comb6[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[38]), .B1(comb6[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16590), .COUT(n16591), .S0(n180_adj_5962), 
          .S1(n177_adj_5961));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3720_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3720_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[36]), .B1(comb6[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16590), .S1(n183_adj_5963));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3720_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3720_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3720_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3720_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3723_add_4_16 (.A0(amdemod_out_d_11__N_2567), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2564), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16588), .S1(amdemod_out_d_11__N_2379[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3723_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_3723_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3723_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3723_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3723_add_4_14 (.A0(amdemod_out_d_11__N_2573), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2570), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16587), .COUT(n16588), .S0(amdemod_out_d_11__N_2379[11]), 
          .S1(amdemod_out_d_11__N_2379[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3723_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_3723_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_3723_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3723_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3723_add_4_12 (.A0(amdemod_out_d_11__N_2579), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2576), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16586), .COUT(n16587), .S0(amdemod_out_d_11__N_2379[9]), 
          .S1(amdemod_out_d_11__N_2379[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3723_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_3723_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_3723_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3723_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3723_add_4_10 (.A0(amdemod_out_d_11__N_2585), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2582), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16585), .COUT(n16586), .S0(amdemod_out_d_11__N_2379[7]), 
          .S1(amdemod_out_d_11__N_2379[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3723_add_4_10.INIT0 = 16'h555f;
    defparam _add_1_3723_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_3723_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3723_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3723_add_4_8 (.A0(square_sum[25]), .B0(n19824), .C0(amdemod_out_d_11__N_2591), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(amdemod_out_d_11__N_2588), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16584), .COUT(n16585), .S0(amdemod_out_d_11__N_2379[5]), 
          .S1(amdemod_out_d_11__N_2379[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3723_add_4_8.INIT0 = 16'he1e1;
    defparam _add_1_3723_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3723_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3723_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3723_add_4_6 (.A0(amdemod_out_d_11__N_2597), .B0(amdemod_out_d_11__N_2370[11]), 
          .C0(amdemod_out_d_11__N_2363), .D0(amdemod_out_d_11__N_2369[11]), 
          .A1(amdemod_out_d_11__N_2594), .B1(square_sum[25]), .C1(n30_adj_6282), 
          .D1(n13890), .CIN(n16583), .COUT(n16584), .S0(amdemod_out_d_11__N_2379[3]), 
          .S1(amdemod_out_d_11__N_2379[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3723_add_4_6.INIT0 = 16'h656a;
    defparam _add_1_3723_add_4_6.INIT1 = 16'h596a;
    defparam _add_1_3723_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3723_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3723_add_4_4 (.A0(n19815), .B0(square_sum[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19815), .B1(amdemod_out_d_11__N_2600), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16582), .COUT(n16583), .S0(amdemod_out_d_11__N_2379[1]), 
          .S1(amdemod_out_d_11__N_2379[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3723_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3723_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3723_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3723_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3723_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16582), .S1(amdemod_out_d_11__N_2379[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3723_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3723_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3723_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3723_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_38 (.A0(integrator_d_tmp[71]), .B0(integrator_tmp[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16581), .S0(n78_adj_5964));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3726_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_36 (.A0(integrator_d_tmp[69]), .B0(integrator_tmp[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[70]), .B1(integrator_tmp[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16580), .COUT(n16581), .S0(n84_adj_5966), 
          .S1(n81_adj_5965));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_34 (.A0(integrator_d_tmp[67]), .B0(integrator_tmp[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[68]), .B1(integrator_tmp[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16579), .COUT(n16580), .S0(n90_adj_5968), 
          .S1(n87_adj_5967));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_32 (.A0(integrator_d_tmp[65]), .B0(integrator_tmp[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[66]), .B1(integrator_tmp[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16578), .COUT(n16579), .S0(n96_adj_5970), 
          .S1(n93_adj_5969));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_30 (.A0(integrator_d_tmp[63]), .B0(integrator_tmp[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[64]), .B1(integrator_tmp[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16577), .COUT(n16578), .S0(n102_adj_5972), 
          .S1(n99_adj_5971));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_28 (.A0(integrator_d_tmp[61]), .B0(integrator_tmp[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[62]), .B1(integrator_tmp[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16576), .COUT(n16577), .S0(n108_adj_5974), 
          .S1(n105_adj_5973));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_26 (.A0(integrator_d_tmp[59]), .B0(integrator_tmp[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[60]), .B1(integrator_tmp[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16575), .COUT(n16576), .S0(n114_adj_5976), 
          .S1(n111_adj_5975));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_24 (.A0(integrator_d_tmp[57]), .B0(integrator_tmp[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[58]), .B1(integrator_tmp[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16574), .COUT(n16575), .S0(n120_adj_5978), 
          .S1(n117_adj_5977));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_22 (.A0(integrator_d_tmp[55]), .B0(integrator_tmp[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[56]), .B1(integrator_tmp[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16573), .COUT(n16574), .S0(n126_adj_5980), 
          .S1(n123_adj_5979));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_20 (.A0(integrator_d_tmp[53]), .B0(integrator_tmp[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[54]), .B1(integrator_tmp[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16572), .COUT(n16573), .S0(n132_adj_5982), 
          .S1(n129_adj_5981));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_18 (.A0(integrator_d_tmp[51]), .B0(integrator_tmp[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[52]), .B1(integrator_tmp[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16571), .COUT(n16572), .S0(n138_adj_5984), 
          .S1(n135_adj_5983));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_16 (.A0(integrator_d_tmp[49]), .B0(integrator_tmp[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[50]), .B1(integrator_tmp[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16570), .COUT(n16571), .S0(n144_adj_5986), 
          .S1(n141_adj_5985));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_14 (.A0(integrator_d_tmp[47]), .B0(integrator_tmp[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[48]), .B1(integrator_tmp[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16569), .COUT(n16570), .S0(n150_adj_5988), 
          .S1(n147_adj_5987));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_12 (.A0(integrator_d_tmp[45]), .B0(integrator_tmp[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[46]), .B1(integrator_tmp[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16568), .COUT(n16569), .S0(n156_adj_5990), 
          .S1(n153_adj_5989));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_10 (.A0(integrator_d_tmp[43]), .B0(integrator_tmp[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[44]), .B1(integrator_tmp[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16567), .COUT(n16568), .S0(n162_adj_5992), 
          .S1(n159_adj_5991));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_8 (.A0(integrator_d_tmp[41]), .B0(integrator_tmp[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[42]), .B1(integrator_tmp[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16566), .COUT(n16567), .S0(n168_adj_5994), 
          .S1(n165_adj_5993));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_6 (.A0(integrator_d_tmp[39]), .B0(integrator_tmp[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[40]), .B1(integrator_tmp[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16565), .COUT(n16566), .S0(n174_adj_5996), 
          .S1(n171_adj_5995));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_4 (.A0(integrator_d_tmp[37]), .B0(integrator_tmp[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[38]), .B1(integrator_tmp[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16564), .COUT(n16565), .S0(n180_adj_5998), 
          .S1(n177_adj_5997));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3726_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3726_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator_d_tmp[36]), .B1(integrator_tmp[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16564), .S1(n183_adj_5999));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3726_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3726_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3726_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3726_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3729_add_4_16 (.A0(amdemod_out_d_11__N_2645), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2642), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16562), .S1(amdemod_out_d_11__N_2389[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3729_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_3729_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3729_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3729_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3729_add_4_14 (.A0(amdemod_out_d_11__N_2651), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2648), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16561), .COUT(n16562), .S0(amdemod_out_d_11__N_2389[11]), 
          .S1(amdemod_out_d_11__N_2389[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3729_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_3729_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_3729_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3729_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3729_add_4_12 (.A0(amdemod_out_d_11__N_2657), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2654), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16560), .COUT(n16561), .S0(amdemod_out_d_11__N_2389[9]), 
          .S1(amdemod_out_d_11__N_2389[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3729_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_3729_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_3729_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3729_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3729_add_4_10 (.A0(square_sum[25]), .B0(n19824), .C0(amdemod_out_d_11__N_2663), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(amdemod_out_d_11__N_2660), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16559), .COUT(n16560), .S0(amdemod_out_d_11__N_2389[7]), 
          .S1(amdemod_out_d_11__N_2389[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3729_add_4_10.INIT0 = 16'he1e1;
    defparam _add_1_3729_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3729_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3729_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3729_add_4_8 (.A0(amdemod_out_d_11__N_2669), .B0(amdemod_out_d_11__N_2370[11]), 
          .C0(amdemod_out_d_11__N_2363), .D0(amdemod_out_d_11__N_2369[11]), 
          .A1(amdemod_out_d_11__N_2666), .B1(square_sum[25]), .C1(n30_adj_6282), 
          .D1(n13890), .CIN(n16558), .COUT(n16559), .S0(amdemod_out_d_11__N_2389[5]), 
          .S1(amdemod_out_d_11__N_2389[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3729_add_4_8.INIT0 = 16'h656a;
    defparam _add_1_3729_add_4_8.INIT1 = 16'h596a;
    defparam _add_1_3729_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3729_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3729_add_4_6 (.A0(amdemod_out_d_11__N_2675), .B0(amdemod_out_d_11__N_2380[14]), 
          .C0(n19815), .D0(amdemod_out_d_11__N_2379[14]), .A1(n19815), 
          .B1(amdemod_out_d_11__N_2672), .C1(GND_net), .D1(VCC_net), .CIN(n16557), 
          .COUT(n16558), .S0(amdemod_out_d_11__N_2389[3]), .S1(amdemod_out_d_11__N_2389[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3729_add_4_6.INIT0 = 16'h656a;
    defparam _add_1_3729_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3729_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3729_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3729_add_4_4 (.A0(n19813), .B0(square_sum[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19813), .B1(amdemod_out_d_11__N_2678), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16556), .COUT(n16557), .S0(amdemod_out_d_11__N_2389[1]), 
          .S1(amdemod_out_d_11__N_2389[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3729_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3729_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3729_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3729_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3729_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16556), .S1(amdemod_out_d_11__N_2389[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3729_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3729_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3729_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3729_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3732_add_4_16 (.A0(amdemod_out_d_11__N_2723), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2720), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16554), .S1(amdemod_out_d_11__N_2399[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3732_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_3732_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3732_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3732_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3732_add_4_14 (.A0(amdemod_out_d_11__N_2729), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2726), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16553), .COUT(n16554), .S0(amdemod_out_d_11__N_2399[11]), 
          .S1(amdemod_out_d_11__N_2399[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3732_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_3732_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_3732_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3732_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3732_add_4_12 (.A0(square_sum[25]), .B0(n19824), .C0(amdemod_out_d_11__N_2735), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(amdemod_out_d_11__N_2732), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16552), .COUT(n16553), .S0(amdemod_out_d_11__N_2399[9]), 
          .S1(amdemod_out_d_11__N_2399[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3732_add_4_12.INIT0 = 16'he1e1;
    defparam _add_1_3732_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3732_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3732_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3732_add_4_10 (.A0(amdemod_out_d_11__N_2741), .B0(amdemod_out_d_11__N_2370[11]), 
          .C0(amdemod_out_d_11__N_2363), .D0(amdemod_out_d_11__N_2369[11]), 
          .A1(amdemod_out_d_11__N_2738), .B1(square_sum[25]), .C1(n30_adj_6282), 
          .D1(n13890), .CIN(n16551), .COUT(n16552), .S0(amdemod_out_d_11__N_2399[7]), 
          .S1(amdemod_out_d_11__N_2399[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3732_add_4_10.INIT0 = 16'h656a;
    defparam _add_1_3732_add_4_10.INIT1 = 16'h596a;
    defparam _add_1_3732_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3732_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3732_add_4_8 (.A0(amdemod_out_d_11__N_2747), .B0(amdemod_out_d_11__N_2380[14]), 
          .C0(n19815), .D0(amdemod_out_d_11__N_2379[14]), .A1(n19815), 
          .B1(amdemod_out_d_11__N_2744), .C1(GND_net), .D1(VCC_net), .CIN(n16550), 
          .COUT(n16551), .S0(amdemod_out_d_11__N_2399[5]), .S1(amdemod_out_d_11__N_2399[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3732_add_4_8.INIT0 = 16'h656a;
    defparam _add_1_3732_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3732_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3732_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3732_add_4_6 (.A0(amdemod_out_d_11__N_2753), .B0(amdemod_out_d_11__N_2390[14]), 
          .C0(n19813), .D0(amdemod_out_d_11__N_2389[14]), .A1(n19813), 
          .B1(amdemod_out_d_11__N_2750), .C1(GND_net), .D1(VCC_net), .CIN(n16549), 
          .COUT(n16550), .S0(amdemod_out_d_11__N_2399[3]), .S1(amdemod_out_d_11__N_2399[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3732_add_4_6.INIT0 = 16'h656a;
    defparam _add_1_3732_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3732_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3732_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3732_add_4_4 (.A0(n19811), .B0(square_sum[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19811), .B1(amdemod_out_d_11__N_2756), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16548), .COUT(n16549), .S0(amdemod_out_d_11__N_2399[1]), 
          .S1(amdemod_out_d_11__N_2399[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3732_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3732_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3732_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3732_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3732_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16548), .S1(amdemod_out_d_11__N_2399[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3732_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3732_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3732_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3732_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_38 (.A0(integrator5[71]), .B0(integrator4[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16547), .S0(n78_adj_6000));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3735_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_36 (.A0(integrator5[69]), .B0(integrator4[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[70]), .B1(integrator4[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16546), .COUT(n16547), .S0(n84_adj_6002), 
          .S1(n81_adj_6001));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_34 (.A0(integrator5[67]), .B0(integrator4[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[68]), .B1(integrator4[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16545), .COUT(n16546), .S0(n90_adj_6004), 
          .S1(n87_adj_6003));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_32 (.A0(integrator5[65]), .B0(integrator4[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[66]), .B1(integrator4[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16544), .COUT(n16545), .S0(n96_adj_6006), 
          .S1(n93_adj_6005));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_30 (.A0(integrator5[63]), .B0(integrator4[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[64]), .B1(integrator4[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16543), .COUT(n16544), .S0(n102_adj_6008), 
          .S1(n99_adj_6007));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_28 (.A0(integrator5[61]), .B0(integrator4[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[62]), .B1(integrator4[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16542), .COUT(n16543), .S0(n108_adj_6010), 
          .S1(n105_adj_6009));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_26 (.A0(integrator5[59]), .B0(integrator4[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[60]), .B1(integrator4[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16541), .COUT(n16542), .S0(n114_adj_6012), 
          .S1(n111_adj_6011));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_24 (.A0(integrator5[57]), .B0(integrator4[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[58]), .B1(integrator4[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16540), .COUT(n16541), .S0(n120_adj_6014), 
          .S1(n117_adj_6013));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_22 (.A0(integrator5[55]), .B0(integrator4[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[56]), .B1(integrator4[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16539), .COUT(n16540), .S0(n126_adj_6016), 
          .S1(n123_adj_6015));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_20 (.A0(integrator5[53]), .B0(integrator4[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[54]), .B1(integrator4[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16538), .COUT(n16539), .S0(n132_adj_6018), 
          .S1(n129_adj_6017));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_18 (.A0(integrator5[51]), .B0(integrator4[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[52]), .B1(integrator4[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16537), .COUT(n16538), .S0(n138_adj_6020), 
          .S1(n135_adj_6019));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_16 (.A0(integrator5[49]), .B0(integrator4[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[50]), .B1(integrator4[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16536), .COUT(n16537), .S0(n144_adj_6022), 
          .S1(n141_adj_6021));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_14 (.A0(integrator5[47]), .B0(integrator4[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[48]), .B1(integrator4[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16535), .COUT(n16536), .S0(n150_adj_6024), 
          .S1(n147_adj_6023));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_12 (.A0(integrator5[45]), .B0(integrator4[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[46]), .B1(integrator4[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16534), .COUT(n16535), .S0(n156_adj_6026), 
          .S1(n153_adj_6025));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_10 (.A0(integrator5[43]), .B0(integrator4[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[44]), .B1(integrator4[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16533), .COUT(n16534), .S0(n162_adj_6028), 
          .S1(n159_adj_6027));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_8 (.A0(integrator5[41]), .B0(integrator4[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[42]), .B1(integrator4[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16532), .COUT(n16533), .S0(n168_adj_6030), 
          .S1(n165_adj_6029));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_6 (.A0(integrator5[39]), .B0(integrator4[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[40]), .B1(integrator4[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16531), .COUT(n16532), .S0(n174_adj_6032), 
          .S1(n171_adj_6031));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_4 (.A0(integrator5[37]), .B0(integrator4[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[38]), .B1(integrator4[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16530), .COUT(n16531), .S0(n180_adj_6034), 
          .S1(n177_adj_6033));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3735_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3735_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[36]), .B1(integrator4[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16530), .S1(n183_adj_6035));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3735_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3735_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3735_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3735_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3738_add_4_15 (.A0(amdemod_out_d_11__N_2400[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2400[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16528), .S1(n34_adj_6036));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3738_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3738_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3738_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3738_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3738_add_4_13 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2400[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2400[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16527), .COUT(n16528), 
          .S0(n43_adj_6038), .S1(n40_adj_6037));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3738_add_4_13.INIT0 = 16'h666a;
    defparam _add_1_3738_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3738_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3738_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3738_add_4_11 (.A0(amdemod_out_d_11__N_2363), .B0(amdemod_out_d_11__N_2400[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2400[8]), .D1(VCC_net), .CIN(n16526), 
          .COUT(n16527), .S0(n49_adj_6040), .S1(n46_adj_6039));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3738_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_3738_add_4_11.INIT1 = 16'h1e1e;
    defparam _add_1_3738_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3738_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3738_add_4_9 (.A0(n19815), .B0(amdemod_out_d_11__N_2400[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(n19816), .B1(amdemod_out_d_11__N_2400[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16525), .COUT(n16526), .S0(n55_adj_6042), 
          .S1(n52_adj_6041));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3738_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_3738_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_3738_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3738_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3738_add_4_7 (.A0(n19813), .B0(amdemod_out_d_11__N_2400[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(n19814), .B1(amdemod_out_d_11__N_2400[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16524), .COUT(n16525), .S0(n61_adj_6044), 
          .S1(n58_adj_6043));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3738_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_3738_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_3738_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3738_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3738_add_4_5 (.A0(n19811), .B0(amdemod_out_d_11__N_2400[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n19812), .B1(amdemod_out_d_11__N_2400[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16523), .COUT(n16524), .S0(n67_adj_6046), 
          .S1(n64_adj_6045));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3738_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3738_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_3738_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3738_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3738_add_4_3 (.A0(square_sum[5]), .B0(amdemod_out_d_11__N_2400[14]), 
          .C0(n19811), .D0(amdemod_out_d_11__N_2399[14]), .A1(n19810), 
          .B1(amdemod_out_d_11__N_2400[0]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16522), .COUT(n16523), .S0(n73), .S1(n70_adj_6047));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3738_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_3738_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3738_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3738_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3738_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16522), .S1(n76_adj_6048));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3738_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3738_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3738_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3738_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3741_add_4_15 (.A0(amdemod_out_d_11__N_2399[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2399[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16520), .S1(n34_adj_6049));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3741_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3741_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3741_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3741_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3741_add_4_13 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2399[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2399[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16519), .COUT(n16520), 
          .S0(n43_adj_6051), .S1(n40_adj_6050));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3741_add_4_13.INIT0 = 16'h666a;
    defparam _add_1_3741_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3741_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3741_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3741_add_4_11 (.A0(amdemod_out_d_11__N_2363), .B0(amdemod_out_d_11__N_2399[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2399[8]), .D1(VCC_net), .CIN(n16518), 
          .COUT(n16519), .S0(n49_adj_6053), .S1(n46_adj_6052));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3741_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_3741_add_4_11.INIT1 = 16'h1e1e;
    defparam _add_1_3741_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3741_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3741_add_4_9 (.A0(n19815), .B0(amdemod_out_d_11__N_2399[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(n19816), .B1(amdemod_out_d_11__N_2399[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16517), .COUT(n16518), .S0(n55_adj_6055), 
          .S1(n52_adj_6054));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3741_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_3741_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_3741_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3741_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3741_add_4_7 (.A0(n19813), .B0(amdemod_out_d_11__N_2399[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(n19814), .B1(amdemod_out_d_11__N_2399[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16516), .COUT(n16517), .S0(n61_adj_6057), 
          .S1(n58_adj_6056));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3741_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_3741_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_3741_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3741_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3741_add_4_5 (.A0(n19811), .B0(amdemod_out_d_11__N_2399[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n19812), .B1(amdemod_out_d_11__N_2399[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16515), .COUT(n16516), .S0(n67_adj_6059), 
          .S1(n64_adj_6058));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3741_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3741_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_3741_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3741_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3741_add_4_3 (.A0(square_sum[5]), .B0(amdemod_out_d_11__N_2400[14]), 
          .C0(n19811), .D0(amdemod_out_d_11__N_2399[14]), .A1(n19810), 
          .B1(amdemod_out_d_11__N_2399[0]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16514), .COUT(n16515), .S0(n73_adj_6061), .S1(n70_adj_6060));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3741_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_3741_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3741_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3741_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3741_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16514), .S1(n76_adj_6062));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3741_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3741_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3741_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3741_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3744_add_4_15 (.A0(amdemod_out_d_11__N_2390[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2390[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16512), .S1(n34_adj_6063));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3744_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3744_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3744_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3744_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3744_add_4_13 (.A0(amdemod_out_d_11__N_2390[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2390[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16511), .COUT(n16512), 
          .S0(n43_adj_6065), .S1(n40_adj_6064));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3744_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3744_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3744_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3744_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3744_add_4_11 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2390[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2390[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16510), .COUT(n16511), 
          .S0(n49_adj_6067), .S1(n46_adj_6066));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3744_add_4_11.INIT0 = 16'h666a;
    defparam _add_1_3744_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3744_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3744_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3744_add_4_9 (.A0(amdemod_out_d_11__N_2363), .B0(amdemod_out_d_11__N_2390[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2390[6]), .D1(VCC_net), .CIN(n16509), 
          .COUT(n16510), .S0(n55_adj_6069), .S1(n52_adj_6068));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3744_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_3744_add_4_9.INIT1 = 16'h1e1e;
    defparam _add_1_3744_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3744_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3744_add_4_7 (.A0(n19815), .B0(amdemod_out_d_11__N_2390[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(n19816), .B1(amdemod_out_d_11__N_2390[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16508), .COUT(n16509), .S0(n61_adj_6071), 
          .S1(n58_adj_6070));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3744_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_3744_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_3744_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3744_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3744_add_4_5 (.A0(n19813), .B0(amdemod_out_d_11__N_2390[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n19814), .B1(amdemod_out_d_11__N_2390[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16507), .COUT(n16508), .S0(n67_adj_6073), 
          .S1(n64_adj_6072));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3744_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3744_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_3744_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3744_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3744_add_4_3 (.A0(square_sum[9]), .B0(amdemod_out_d_11__N_2390[14]), 
          .C0(n19813), .D0(amdemod_out_d_11__N_2389[14]), .A1(n19812), 
          .B1(amdemod_out_d_11__N_2390[0]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16506), .COUT(n16507), .S0(n73_adj_6075), .S1(n70_adj_6074));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3744_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_3744_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3744_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3744_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3744_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16506), .S1(n76_adj_6076));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3744_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3744_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3744_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3744_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3747_add_4_15 (.A0(amdemod_out_d_11__N_2389[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2389[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16504), .S1(n34_adj_6077));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3747_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3747_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3747_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3747_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3747_add_4_13 (.A0(amdemod_out_d_11__N_2389[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2389[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16503), .COUT(n16504), 
          .S0(n43_adj_6079), .S1(n40_adj_6078));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3747_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3747_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3747_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3747_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3747_add_4_11 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2389[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2389[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16502), .COUT(n16503), 
          .S0(n49_adj_6081), .S1(n46_adj_6080));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3747_add_4_11.INIT0 = 16'h666a;
    defparam _add_1_3747_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3747_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3747_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3747_add_4_9 (.A0(amdemod_out_d_11__N_2363), .B0(amdemod_out_d_11__N_2389[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2389[6]), .D1(VCC_net), .CIN(n16501), 
          .COUT(n16502), .S0(n55_adj_6083), .S1(n52_adj_6082));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3747_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_3747_add_4_9.INIT1 = 16'h1e1e;
    defparam _add_1_3747_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3747_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3747_add_4_7 (.A0(n19815), .B0(amdemod_out_d_11__N_2389[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(n19816), .B1(amdemod_out_d_11__N_2389[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16500), .COUT(n16501), .S0(n61_adj_6085), 
          .S1(n58_adj_6084));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3747_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_3747_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_3747_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3747_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3747_add_4_5 (.A0(n19813), .B0(amdemod_out_d_11__N_2389[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n19814), .B1(amdemod_out_d_11__N_2389[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16499), .COUT(n16500), .S0(n67_adj_6087), 
          .S1(n64_adj_6086));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3747_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3747_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_3747_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3747_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3747_add_4_3 (.A0(square_sum[9]), .B0(amdemod_out_d_11__N_2390[14]), 
          .C0(n19813), .D0(amdemod_out_d_11__N_2389[14]), .A1(n19812), 
          .B1(amdemod_out_d_11__N_2389[0]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16498), .COUT(n16499), .S0(n73_adj_6089), .S1(n70_adj_6088));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3747_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_3747_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3747_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3747_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3747_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16498), .S1(n76_adj_6090));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3747_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3747_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3747_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3747_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16497), .S0(cout_adj_6091));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_3540_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_3540_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_36 (.A0(integrator4_adj_6561[34]), .B0(integrator3_adj_6560[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[35]), .B1(integrator3_adj_6560[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16496), .COUT(n16497), .S0(integrator4_71__N_1176_adj_6576[34]), 
          .S1(integrator4_71__N_1176_adj_6576[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_34 (.A0(integrator4_adj_6561[32]), .B0(integrator3_adj_6560[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[33]), .B1(integrator3_adj_6560[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16495), .COUT(n16496), .S0(integrator4_71__N_1176_adj_6576[32]), 
          .S1(integrator4_71__N_1176_adj_6576[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_32 (.A0(integrator4_adj_6561[30]), .B0(integrator3_adj_6560[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[31]), .B1(integrator3_adj_6560[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16494), .COUT(n16495), .S0(integrator4_71__N_1176_adj_6576[30]), 
          .S1(integrator4_71__N_1176_adj_6576[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_30 (.A0(integrator4_adj_6561[28]), .B0(integrator3_adj_6560[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[29]), .B1(integrator3_adj_6560[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16493), .COUT(n16494), .S0(integrator4_71__N_1176_adj_6576[28]), 
          .S1(integrator4_71__N_1176_adj_6576[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_28 (.A0(integrator4_adj_6561[26]), .B0(integrator3_adj_6560[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[27]), .B1(integrator3_adj_6560[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16492), .COUT(n16493), .S0(integrator4_71__N_1176_adj_6576[26]), 
          .S1(integrator4_71__N_1176_adj_6576[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_26 (.A0(integrator4_adj_6561[24]), .B0(integrator3_adj_6560[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[25]), .B1(integrator3_adj_6560[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16491), .COUT(n16492), .S0(integrator4_71__N_1176_adj_6576[24]), 
          .S1(integrator4_71__N_1176_adj_6576[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_24 (.A0(integrator4_adj_6561[22]), .B0(integrator3_adj_6560[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[23]), .B1(integrator3_adj_6560[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16490), .COUT(n16491), .S0(integrator4_71__N_1176_adj_6576[22]), 
          .S1(integrator4_71__N_1176_adj_6576[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_22 (.A0(integrator4_adj_6561[20]), .B0(integrator3_adj_6560[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[21]), .B1(integrator3_adj_6560[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16489), .COUT(n16490), .S0(integrator4_71__N_1176_adj_6576[20]), 
          .S1(integrator4_71__N_1176_adj_6576[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_20 (.A0(integrator4_adj_6561[18]), .B0(integrator3_adj_6560[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[19]), .B1(integrator3_adj_6560[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16488), .COUT(n16489), .S0(integrator4_71__N_1176_adj_6576[18]), 
          .S1(integrator4_71__N_1176_adj_6576[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_18 (.A0(integrator4_adj_6561[16]), .B0(integrator3_adj_6560[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[17]), .B1(integrator3_adj_6560[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16487), .COUT(n16488), .S0(integrator4_71__N_1176_adj_6576[16]), 
          .S1(integrator4_71__N_1176_adj_6576[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_16 (.A0(integrator4_adj_6561[14]), .B0(integrator3_adj_6560[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[15]), .B1(integrator3_adj_6560[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16486), .COUT(n16487), .S0(integrator4_71__N_1176_adj_6576[14]), 
          .S1(integrator4_71__N_1176_adj_6576[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_14 (.A0(integrator4_adj_6561[12]), .B0(integrator3_adj_6560[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[13]), .B1(integrator3_adj_6560[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16485), .COUT(n16486), .S0(integrator4_71__N_1176_adj_6576[12]), 
          .S1(integrator4_71__N_1176_adj_6576[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_12 (.A0(integrator4_adj_6561[10]), .B0(integrator3_adj_6560[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[11]), .B1(integrator3_adj_6560[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16484), .COUT(n16485), .S0(integrator4_71__N_1176_adj_6576[10]), 
          .S1(integrator4_71__N_1176_adj_6576[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_10 (.A0(integrator4_adj_6561[8]), .B0(integrator3_adj_6560[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[9]), .B1(integrator3_adj_6560[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16483), .COUT(n16484), .S0(integrator4_71__N_1176_adj_6576[8]), 
          .S1(integrator4_71__N_1176_adj_6576[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_8 (.A0(integrator4_adj_6561[6]), .B0(integrator3_adj_6560[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[7]), .B1(integrator3_adj_6560[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16482), .COUT(n16483), .S0(integrator4_71__N_1176_adj_6576[6]), 
          .S1(integrator4_71__N_1176_adj_6576[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_6 (.A0(integrator4_adj_6561[4]), .B0(integrator3_adj_6560[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[5]), .B1(integrator3_adj_6560[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16481), .COUT(n16482), .S0(integrator4_71__N_1176_adj_6576[4]), 
          .S1(integrator4_71__N_1176_adj_6576[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_4 (.A0(integrator4_adj_6561[2]), .B0(integrator3_adj_6560[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[3]), .B1(integrator3_adj_6560[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16480), .COUT(n16481), .S0(integrator4_71__N_1176_adj_6576[2]), 
          .S1(integrator4_71__N_1176_adj_6576[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3540_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3540_add_4_2 (.A0(integrator4_adj_6561[0]), .B0(integrator3_adj_6560[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[1]), .B1(integrator3_adj_6560[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16480), .S1(integrator4_71__N_1176_adj_6576[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3540_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_3540_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3540_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3540_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16478), .S0(cout_adj_6092));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_3543_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_3543_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_36 (.A0(integrator5_adj_6562[34]), .B0(integrator4_adj_6561[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[35]), .B1(integrator4_adj_6561[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16477), .COUT(n16478), .S0(integrator5_71__N_1248_adj_6577[34]), 
          .S1(integrator5_71__N_1248_adj_6577[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_34 (.A0(integrator5_adj_6562[32]), .B0(integrator4_adj_6561[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[33]), .B1(integrator4_adj_6561[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16476), .COUT(n16477), .S0(integrator5_71__N_1248_adj_6577[32]), 
          .S1(integrator5_71__N_1248_adj_6577[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_32 (.A0(integrator5_adj_6562[30]), .B0(integrator4_adj_6561[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[31]), .B1(integrator4_adj_6561[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16475), .COUT(n16476), .S0(integrator5_71__N_1248_adj_6577[30]), 
          .S1(integrator5_71__N_1248_adj_6577[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_30 (.A0(integrator5_adj_6562[28]), .B0(integrator4_adj_6561[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[29]), .B1(integrator4_adj_6561[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16474), .COUT(n16475), .S0(integrator5_71__N_1248_adj_6577[28]), 
          .S1(integrator5_71__N_1248_adj_6577[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_28 (.A0(integrator5_adj_6562[26]), .B0(integrator4_adj_6561[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[27]), .B1(integrator4_adj_6561[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16473), .COUT(n16474), .S0(integrator5_71__N_1248_adj_6577[26]), 
          .S1(integrator5_71__N_1248_adj_6577[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_26 (.A0(integrator5_adj_6562[24]), .B0(integrator4_adj_6561[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[25]), .B1(integrator4_adj_6561[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16472), .COUT(n16473), .S0(integrator5_71__N_1248_adj_6577[24]), 
          .S1(integrator5_71__N_1248_adj_6577[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_24 (.A0(integrator5_adj_6562[22]), .B0(integrator4_adj_6561[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[23]), .B1(integrator4_adj_6561[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16471), .COUT(n16472), .S0(integrator5_71__N_1248_adj_6577[22]), 
          .S1(integrator5_71__N_1248_adj_6577[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_22 (.A0(integrator5_adj_6562[20]), .B0(integrator4_adj_6561[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[21]), .B1(integrator4_adj_6561[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16470), .COUT(n16471), .S0(integrator5_71__N_1248_adj_6577[20]), 
          .S1(integrator5_71__N_1248_adj_6577[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_20 (.A0(integrator5_adj_6562[18]), .B0(integrator4_adj_6561[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[19]), .B1(integrator4_adj_6561[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16469), .COUT(n16470), .S0(integrator5_71__N_1248_adj_6577[18]), 
          .S1(integrator5_71__N_1248_adj_6577[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_18 (.A0(integrator5_adj_6562[16]), .B0(integrator4_adj_6561[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[17]), .B1(integrator4_adj_6561[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16468), .COUT(n16469), .S0(integrator5_71__N_1248_adj_6577[16]), 
          .S1(integrator5_71__N_1248_adj_6577[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_16 (.A0(integrator5_adj_6562[14]), .B0(integrator4_adj_6561[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[15]), .B1(integrator4_adj_6561[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16467), .COUT(n16468), .S0(integrator5_71__N_1248_adj_6577[14]), 
          .S1(integrator5_71__N_1248_adj_6577[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_14 (.A0(integrator5_adj_6562[12]), .B0(integrator4_adj_6561[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[13]), .B1(integrator4_adj_6561[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16466), .COUT(n16467), .S0(integrator5_71__N_1248_adj_6577[12]), 
          .S1(integrator5_71__N_1248_adj_6577[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_12 (.A0(integrator5_adj_6562[10]), .B0(integrator4_adj_6561[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[11]), .B1(integrator4_adj_6561[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16465), .COUT(n16466), .S0(integrator5_71__N_1248_adj_6577[10]), 
          .S1(integrator5_71__N_1248_adj_6577[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_10 (.A0(integrator5_adj_6562[8]), .B0(integrator4_adj_6561[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[9]), .B1(integrator4_adj_6561[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16464), .COUT(n16465), .S0(integrator5_71__N_1248_adj_6577[8]), 
          .S1(integrator5_71__N_1248_adj_6577[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_8 (.A0(integrator5_adj_6562[6]), .B0(integrator4_adj_6561[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[7]), .B1(integrator4_adj_6561[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16463), .COUT(n16464), .S0(integrator5_71__N_1248_adj_6577[6]), 
          .S1(integrator5_71__N_1248_adj_6577[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_6 (.A0(integrator5_adj_6562[4]), .B0(integrator4_adj_6561[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[5]), .B1(integrator4_adj_6561[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16462), .COUT(n16463), .S0(integrator5_71__N_1248_adj_6577[4]), 
          .S1(integrator5_71__N_1248_adj_6577[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3543_add_4_4 (.A0(integrator5_adj_6562[2]), .B0(integrator4_adj_6561[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[3]), .B1(integrator4_adj_6561[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16461), .COUT(n16462), .S0(integrator5_71__N_1248_adj_6577[2]), 
          .S1(integrator5_71__N_1248_adj_6577[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3543_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_4.INJECT1_1 = "NO";
    PFUMX i8707 (.BLUT(n19764), .ALUT(n19763), .C0(rx_byte[2]), .Z(n19765));
    PFUMX i8704 (.BLUT(n19761), .ALUT(n19760), .C0(rx_byte[2]), .Z(n19762));
    CCU2C _add_1_3543_add_4_2 (.A0(integrator5_adj_6562[0]), .B0(integrator4_adj_6561[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[1]), .B1(integrator4_adj_6561[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16461), .S1(integrator5_71__N_1248_adj_6577[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3543_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_3543_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3543_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3543_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16459), .S0(cout_adj_5318));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_3510_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_3510_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_36 (.A0(integrator2[34]), .B0(integrator1[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[35]), .B1(integrator1[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16458), .COUT(n16459), .S0(integrator2_71__N_1032[34]), 
          .S1(integrator2_71__N_1032[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_34 (.A0(integrator2[32]), .B0(integrator1[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[33]), .B1(integrator1[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16457), .COUT(n16458), .S0(integrator2_71__N_1032[32]), 
          .S1(integrator2_71__N_1032[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_32 (.A0(integrator2[30]), .B0(integrator1[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[31]), .B1(integrator1[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16456), .COUT(n16457), .S0(integrator2_71__N_1032[30]), 
          .S1(integrator2_71__N_1032[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_30 (.A0(integrator2[28]), .B0(integrator1[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[29]), .B1(integrator1[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16455), .COUT(n16456), .S0(integrator2_71__N_1032[28]), 
          .S1(integrator2_71__N_1032[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_28 (.A0(integrator2[26]), .B0(integrator1[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[27]), .B1(integrator1[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16454), .COUT(n16455), .S0(integrator2_71__N_1032[26]), 
          .S1(integrator2_71__N_1032[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_26 (.A0(integrator2[24]), .B0(integrator1[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[25]), .B1(integrator1[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16453), .COUT(n16454), .S0(integrator2_71__N_1032[24]), 
          .S1(integrator2_71__N_1032[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_24 (.A0(integrator2[22]), .B0(integrator1[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[23]), .B1(integrator1[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16452), .COUT(n16453), .S0(integrator2_71__N_1032[22]), 
          .S1(integrator2_71__N_1032[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_22 (.A0(integrator2[20]), .B0(integrator1[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[21]), .B1(integrator1[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16451), .COUT(n16452), .S0(integrator2_71__N_1032[20]), 
          .S1(integrator2_71__N_1032[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_20 (.A0(integrator2[18]), .B0(integrator1[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[19]), .B1(integrator1[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16450), .COUT(n16451), .S0(integrator2_71__N_1032[18]), 
          .S1(integrator2_71__N_1032[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_18 (.A0(integrator2[16]), .B0(integrator1[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[17]), .B1(integrator1[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16449), .COUT(n16450), .S0(integrator2_71__N_1032[16]), 
          .S1(integrator2_71__N_1032[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_16 (.A0(integrator2[14]), .B0(integrator1[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[15]), .B1(integrator1[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16448), .COUT(n16449), .S0(integrator2_71__N_1032[14]), 
          .S1(integrator2_71__N_1032[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_14 (.A0(integrator2[12]), .B0(integrator1[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[13]), .B1(integrator1[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16447), .COUT(n16448), .S0(integrator2_71__N_1032[12]), 
          .S1(integrator2_71__N_1032[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_12 (.A0(integrator2[10]), .B0(integrator1[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[11]), .B1(integrator1[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16446), .COUT(n16447), .S0(integrator2_71__N_1032[10]), 
          .S1(integrator2_71__N_1032[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_10 (.A0(integrator2[8]), .B0(integrator1[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[9]), .B1(integrator1[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16445), .COUT(n16446), .S0(integrator2_71__N_1032[8]), 
          .S1(integrator2_71__N_1032[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_8 (.A0(integrator2[6]), .B0(integrator1[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[7]), .B1(integrator1[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16444), .COUT(n16445), .S0(integrator2_71__N_1032[6]), 
          .S1(integrator2_71__N_1032[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_6 (.A0(integrator2[4]), .B0(integrator1[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[5]), .B1(integrator1[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16443), .COUT(n16444), .S0(integrator2_71__N_1032[4]), 
          .S1(integrator2_71__N_1032[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_4 (.A0(integrator2[2]), .B0(integrator1[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[3]), .B1(integrator1[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16442), .COUT(n16443), .S0(integrator2_71__N_1032[2]), 
          .S1(integrator2_71__N_1032[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3510_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3510_add_4_2 (.A0(integrator2[0]), .B0(integrator1[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[1]), .B1(integrator1[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16442), .S1(integrator2_71__N_1032[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3510_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_3510_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3510_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3510_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16440), .S0(cout_adj_5296));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_3513_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_3513_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_36 (.A0(integrator3[34]), .B0(integrator2[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[35]), .B1(integrator2[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16439), .COUT(n16440), .S0(integrator3_71__N_1104[34]), 
          .S1(integrator3_71__N_1104[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_34 (.A0(integrator3[32]), .B0(integrator2[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[33]), .B1(integrator2[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16438), .COUT(n16439), .S0(integrator3_71__N_1104[32]), 
          .S1(integrator3_71__N_1104[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_32 (.A0(integrator3[30]), .B0(integrator2[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[31]), .B1(integrator2[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16437), .COUT(n16438), .S0(integrator3_71__N_1104[30]), 
          .S1(integrator3_71__N_1104[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_30 (.A0(integrator3[28]), .B0(integrator2[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[29]), .B1(integrator2[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16436), .COUT(n16437), .S0(integrator3_71__N_1104[28]), 
          .S1(integrator3_71__N_1104[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_28 (.A0(integrator3[26]), .B0(integrator2[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[27]), .B1(integrator2[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16435), .COUT(n16436), .S0(integrator3_71__N_1104[26]), 
          .S1(integrator3_71__N_1104[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_26 (.A0(integrator3[24]), .B0(integrator2[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[25]), .B1(integrator2[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16434), .COUT(n16435), .S0(integrator3_71__N_1104[24]), 
          .S1(integrator3_71__N_1104[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_24 (.A0(integrator3[22]), .B0(integrator2[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[23]), .B1(integrator2[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16433), .COUT(n16434), .S0(integrator3_71__N_1104[22]), 
          .S1(integrator3_71__N_1104[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_22 (.A0(integrator3[20]), .B0(integrator2[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[21]), .B1(integrator2[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16432), .COUT(n16433), .S0(integrator3_71__N_1104[20]), 
          .S1(integrator3_71__N_1104[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_20 (.A0(integrator3[18]), .B0(integrator2[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[19]), .B1(integrator2[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16431), .COUT(n16432), .S0(integrator3_71__N_1104[18]), 
          .S1(integrator3_71__N_1104[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_18 (.A0(integrator3[16]), .B0(integrator2[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[17]), .B1(integrator2[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16430), .COUT(n16431), .S0(integrator3_71__N_1104[16]), 
          .S1(integrator3_71__N_1104[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_16 (.A0(integrator3[14]), .B0(integrator2[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[15]), .B1(integrator2[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16429), .COUT(n16430), .S0(integrator3_71__N_1104[14]), 
          .S1(integrator3_71__N_1104[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_14 (.A0(integrator3[12]), .B0(integrator2[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[13]), .B1(integrator2[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16428), .COUT(n16429), .S0(integrator3_71__N_1104[12]), 
          .S1(integrator3_71__N_1104[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_12 (.A0(integrator3[10]), .B0(integrator2[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[11]), .B1(integrator2[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16427), .COUT(n16428), .S0(integrator3_71__N_1104[10]), 
          .S1(integrator3_71__N_1104[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_10 (.A0(integrator3[8]), .B0(integrator2[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[9]), .B1(integrator2[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16426), .COUT(n16427), .S0(integrator3_71__N_1104[8]), 
          .S1(integrator3_71__N_1104[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_8 (.A0(integrator3[6]), .B0(integrator2[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[7]), .B1(integrator2[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16425), .COUT(n16426), .S0(integrator3_71__N_1104[6]), 
          .S1(integrator3_71__N_1104[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_6 (.A0(integrator3[4]), .B0(integrator2[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[5]), .B1(integrator2[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16424), .COUT(n16425), .S0(integrator3_71__N_1104[4]), 
          .S1(integrator3_71__N_1104[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_4 (.A0(integrator3[2]), .B0(integrator2[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[3]), .B1(integrator2[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16423), .COUT(n16424), .S0(integrator3_71__N_1104[2]), 
          .S1(integrator3_71__N_1104[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3513_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3513_add_4_2 (.A0(integrator3[0]), .B0(integrator2[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[1]), .B1(integrator2[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16423), .S1(integrator3_71__N_1104[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3513_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_3513_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3513_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3513_add_4_2.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_0__bdd_4_lut_8558 (.A(phase_increment_1__63__N_21[0]), 
         .B(rx_byte[2]), .C(led_0_6), .D(rx_byte[0]), .Z(n19574)) /* synthesis lut_function=(!((B (C)+!B (D))+!A)) */ ;
    defparam phase_increment_1__63__N_21_0__bdd_4_lut_8558.init = 16'h082a;
    CCU2C _add_1_3672_add_4_38 (.A0(comb_d9_adj_6570[71]), .B0(comb9_adj_6569[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16421), .S0(n78_adj_5612));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3672_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_36 (.A0(comb_d9_adj_6570[69]), .B0(comb9_adj_6569[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[70]), .B1(comb9_adj_6569[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16420), .COUT(n16421), .S0(n84_adj_5614), 
          .S1(n81_adj_5613));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_34 (.A0(comb_d9_adj_6570[67]), .B0(comb9_adj_6569[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[68]), .B1(comb9_adj_6569[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16419), .COUT(n16420), .S0(n90_adj_5616), 
          .S1(n87_adj_5615));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_32 (.A0(comb_d9_adj_6570[65]), .B0(comb9_adj_6569[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[66]), .B1(comb9_adj_6569[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16418), .COUT(n16419), .S0(n96_adj_5618), 
          .S1(n93_adj_5617));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_30 (.A0(comb_d9_adj_6570[63]), .B0(comb9_adj_6569[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[64]), .B1(comb9_adj_6569[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16417), .COUT(n16418), .S0(n102_adj_5620), 
          .S1(n99_adj_5619));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_28 (.A0(comb_d9_adj_6570[61]), .B0(comb9_adj_6569[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[62]), .B1(comb9_adj_6569[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16416), .COUT(n16417), .S0(n108_adj_5622), 
          .S1(n105_adj_5621));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_26 (.A0(comb_d9_adj_6570[59]), .B0(comb9_adj_6569[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[60]), .B1(comb9_adj_6569[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16415), .COUT(n16416), .S0(n114_adj_5624), 
          .S1(n111_adj_5623));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_24 (.A0(comb_d9_adj_6570[57]), .B0(comb9_adj_6569[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[58]), .B1(comb9_adj_6569[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16414), .COUT(n16415), .S0(n120_adj_5626), 
          .S1(n117_adj_5625));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_22 (.A0(comb_d9_adj_6570[55]), .B0(comb9_adj_6569[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[56]), .B1(comb9_adj_6569[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16413), .COUT(n16414));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_20 (.A0(comb_d9_adj_6570[53]), .B0(comb9_adj_6569[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[54]), .B1(comb9_adj_6569[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16412), .COUT(n16413));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_18 (.A0(comb_d9_adj_6570[51]), .B0(comb9_adj_6569[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[52]), .B1(comb9_adj_6569[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16411), .COUT(n16412));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_16 (.A0(comb_d9_adj_6570[49]), .B0(comb9_adj_6569[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[50]), .B1(comb9_adj_6569[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16410), .COUT(n16411));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_14 (.A0(comb_d9_adj_6570[47]), .B0(comb9_adj_6569[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[48]), .B1(comb9_adj_6569[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16409), .COUT(n16410));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_12 (.A0(comb_d9_adj_6570[45]), .B0(comb9_adj_6569[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[46]), .B1(comb9_adj_6569[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16408), .COUT(n16409));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_10 (.A0(comb_d9_adj_6570[43]), .B0(comb9_adj_6569[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[44]), .B1(comb9_adj_6569[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16407), .COUT(n16408));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_8 (.A0(comb_d9_adj_6570[41]), .B0(comb9_adj_6569[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[42]), .B1(comb9_adj_6569[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16406), .COUT(n16407));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_6 (.A0(comb_d9_adj_6570[39]), .B0(comb9_adj_6569[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[40]), .B1(comb9_adj_6569[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16405), .COUT(n16406));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_4 (.A0(comb_d9_adj_6570[37]), .B0(comb9_adj_6569[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[38]), .B1(comb9_adj_6569[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16404), .COUT(n16405));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3672_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3672_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9_adj_6570[36]), .B1(comb9_adj_6569[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16404));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3672_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3672_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3672_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3672_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16403), .S0(cout_adj_5327));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_3516_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_3516_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_36 (.A0(integrator4[34]), .B0(integrator3[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[35]), .B1(integrator3[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16402), .COUT(n16403), .S0(integrator4_71__N_1176[34]), 
          .S1(integrator4_71__N_1176[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_34 (.A0(integrator4[32]), .B0(integrator3[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[33]), .B1(integrator3[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16401), .COUT(n16402), .S0(integrator4_71__N_1176[32]), 
          .S1(integrator4_71__N_1176[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_32 (.A0(integrator4[30]), .B0(integrator3[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[31]), .B1(integrator3[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16400), .COUT(n16401), .S0(integrator4_71__N_1176[30]), 
          .S1(integrator4_71__N_1176[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_30 (.A0(integrator4[28]), .B0(integrator3[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[29]), .B1(integrator3[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16399), .COUT(n16400), .S0(integrator4_71__N_1176[28]), 
          .S1(integrator4_71__N_1176[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_28 (.A0(integrator4[26]), .B0(integrator3[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[27]), .B1(integrator3[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16398), .COUT(n16399), .S0(integrator4_71__N_1176[26]), 
          .S1(integrator4_71__N_1176[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_26 (.A0(integrator4[24]), .B0(integrator3[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[25]), .B1(integrator3[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16397), .COUT(n16398), .S0(integrator4_71__N_1176[24]), 
          .S1(integrator4_71__N_1176[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_24 (.A0(integrator4[22]), .B0(integrator3[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[23]), .B1(integrator3[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16396), .COUT(n16397), .S0(integrator4_71__N_1176[22]), 
          .S1(integrator4_71__N_1176[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_22 (.A0(integrator4[20]), .B0(integrator3[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[21]), .B1(integrator3[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16395), .COUT(n16396), .S0(integrator4_71__N_1176[20]), 
          .S1(integrator4_71__N_1176[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_20 (.A0(integrator4[18]), .B0(integrator3[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[19]), .B1(integrator3[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16394), .COUT(n16395), .S0(integrator4_71__N_1176[18]), 
          .S1(integrator4_71__N_1176[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_18 (.A0(integrator4[16]), .B0(integrator3[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[17]), .B1(integrator3[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16393), .COUT(n16394), .S0(integrator4_71__N_1176[16]), 
          .S1(integrator4_71__N_1176[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_16 (.A0(integrator4[14]), .B0(integrator3[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[15]), .B1(integrator3[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16392), .COUT(n16393), .S0(integrator4_71__N_1176[14]), 
          .S1(integrator4_71__N_1176[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_14 (.A0(integrator4[12]), .B0(integrator3[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[13]), .B1(integrator3[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16391), .COUT(n16392), .S0(integrator4_71__N_1176[12]), 
          .S1(integrator4_71__N_1176[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_12 (.A0(integrator4[10]), .B0(integrator3[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[11]), .B1(integrator3[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16390), .COUT(n16391), .S0(integrator4_71__N_1176[10]), 
          .S1(integrator4_71__N_1176[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_10 (.A0(integrator4[8]), .B0(integrator3[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[9]), .B1(integrator3[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16389), .COUT(n16390), .S0(integrator4_71__N_1176[8]), 
          .S1(integrator4_71__N_1176[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_8 (.A0(integrator4[6]), .B0(integrator3[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[7]), .B1(integrator3[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16388), .COUT(n16389), .S0(integrator4_71__N_1176[6]), 
          .S1(integrator4_71__N_1176[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_6 (.A0(integrator4[4]), .B0(integrator3[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[5]), .B1(integrator3[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16387), .COUT(n16388), .S0(integrator4_71__N_1176[4]), 
          .S1(integrator4_71__N_1176[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_4 (.A0(integrator4[2]), .B0(integrator3[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[3]), .B1(integrator3[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16386), .COUT(n16387), .S0(integrator4_71__N_1176[2]), 
          .S1(integrator4_71__N_1176[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3516_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3516_add_4_2 (.A0(integrator4[0]), .B0(integrator3[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[1]), .B1(integrator3[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16386), .S1(integrator4_71__N_1176[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3516_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_3516_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3516_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3516_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16384), .S0(cout_adj_5293));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_3519_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_3519_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_36 (.A0(integrator5[34]), .B0(integrator4[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[35]), .B1(integrator4[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16383), .COUT(n16384), .S0(integrator5_71__N_1248[34]), 
          .S1(integrator5_71__N_1248[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_34 (.A0(integrator5[32]), .B0(integrator4[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[33]), .B1(integrator4[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16382), .COUT(n16383), .S0(integrator5_71__N_1248[32]), 
          .S1(integrator5_71__N_1248[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_32 (.A0(integrator5[30]), .B0(integrator4[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[31]), .B1(integrator4[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16381), .COUT(n16382), .S0(integrator5_71__N_1248[30]), 
          .S1(integrator5_71__N_1248[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_30 (.A0(integrator5[28]), .B0(integrator4[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[29]), .B1(integrator4[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16380), .COUT(n16381), .S0(integrator5_71__N_1248[28]), 
          .S1(integrator5_71__N_1248[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_28 (.A0(integrator5[26]), .B0(integrator4[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[27]), .B1(integrator4[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16379), .COUT(n16380), .S0(integrator5_71__N_1248[26]), 
          .S1(integrator5_71__N_1248[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_26 (.A0(integrator5[24]), .B0(integrator4[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[25]), .B1(integrator4[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16378), .COUT(n16379), .S0(integrator5_71__N_1248[24]), 
          .S1(integrator5_71__N_1248[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_24 (.A0(integrator5[22]), .B0(integrator4[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[23]), .B1(integrator4[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16377), .COUT(n16378), .S0(integrator5_71__N_1248[22]), 
          .S1(integrator5_71__N_1248[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_22 (.A0(integrator5[20]), .B0(integrator4[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[21]), .B1(integrator4[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16376), .COUT(n16377), .S0(integrator5_71__N_1248[20]), 
          .S1(integrator5_71__N_1248[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_20 (.A0(integrator5[18]), .B0(integrator4[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[19]), .B1(integrator4[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16375), .COUT(n16376), .S0(integrator5_71__N_1248[18]), 
          .S1(integrator5_71__N_1248[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_18 (.A0(integrator5[16]), .B0(integrator4[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[17]), .B1(integrator4[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16374), .COUT(n16375), .S0(integrator5_71__N_1248[16]), 
          .S1(integrator5_71__N_1248[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_16 (.A0(integrator5[14]), .B0(integrator4[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[15]), .B1(integrator4[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16373), .COUT(n16374), .S0(integrator5_71__N_1248[14]), 
          .S1(integrator5_71__N_1248[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_14 (.A0(integrator5[12]), .B0(integrator4[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[13]), .B1(integrator4[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16372), .COUT(n16373), .S0(integrator5_71__N_1248[12]), 
          .S1(integrator5_71__N_1248[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_12 (.A0(integrator5[10]), .B0(integrator4[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[11]), .B1(integrator4[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16371), .COUT(n16372), .S0(integrator5_71__N_1248[10]), 
          .S1(integrator5_71__N_1248[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_10 (.A0(integrator5[8]), .B0(integrator4[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[9]), .B1(integrator4[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16370), .COUT(n16371), .S0(integrator5_71__N_1248[8]), 
          .S1(integrator5_71__N_1248[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_8 (.A0(integrator5[6]), .B0(integrator4[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[7]), .B1(integrator4[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16369), .COUT(n16370), .S0(integrator5_71__N_1248[6]), 
          .S1(integrator5_71__N_1248[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_6 (.A0(integrator5[4]), .B0(integrator4[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[5]), .B1(integrator4[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16368), .COUT(n16369), .S0(integrator5_71__N_1248[4]), 
          .S1(integrator5_71__N_1248[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_4 (.A0(integrator5[2]), .B0(integrator4[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[3]), .B1(integrator4[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16367), .COUT(n16368), .S0(integrator5_71__N_1248[2]), 
          .S1(integrator5_71__N_1248[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3519_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3519_add_4_2 (.A0(integrator5[0]), .B0(integrator4[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[1]), .B1(integrator4[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16367), .S1(integrator5_71__N_1248[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3519_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_3519_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3519_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3519_add_4_2.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_0__bdd_3_lut (.A(phase_increment_1__63__N_21[0]), 
         .B(phase_increment_1__63__N_18[0]), .C(rx_byte[0]), .Z(n19575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam phase_increment_1__63__N_21_0__bdd_3_lut.init = 16'hcaca;
    CCU2C _add_1_3522_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16365), .S0(cout_adj_5328));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_3522_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_3522_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_36 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16364), .COUT(n16365), .S0(integrator1_71__N_960_adj_6573[34]), 
          .S1(integrator1_71__N_960_adj_6573[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_34 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16363), .COUT(n16364), .S0(integrator1_71__N_960_adj_6573[32]), 
          .S1(integrator1_71__N_960_adj_6573[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_32 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16362), .COUT(n16363), .S0(integrator1_71__N_960_adj_6573[30]), 
          .S1(integrator1_71__N_960_adj_6573[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_30 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16361), .COUT(n16362), .S0(integrator1_71__N_960_adj_6573[28]), 
          .S1(integrator1_71__N_960_adj_6573[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_28 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16360), .COUT(n16361), .S0(integrator1_71__N_960_adj_6573[26]), 
          .S1(integrator1_71__N_960_adj_6573[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_26 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16359), .COUT(n16360), .S0(integrator1_71__N_960_adj_6573[24]), 
          .S1(integrator1_71__N_960_adj_6573[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_24 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16358), .COUT(n16359), .S0(integrator1_71__N_960_adj_6573[22]), 
          .S1(integrator1_71__N_960_adj_6573[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_22 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16357), .COUT(n16358), .S0(integrator1_71__N_960_adj_6573[20]), 
          .S1(integrator1_71__N_960_adj_6573[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_20 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16356), .COUT(n16357), .S0(integrator1_71__N_960_adj_6573[18]), 
          .S1(integrator1_71__N_960_adj_6573[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_18 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16355), .COUT(n16356), .S0(integrator1_71__N_960_adj_6573[16]), 
          .S1(integrator1_71__N_960_adj_6573[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_16 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16354), .COUT(n16355), .S0(integrator1_71__N_960_adj_6573[14]), 
          .S1(integrator1_71__N_960_adj_6573[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_14 (.A0(mix_cosinewave[11]), .B0(integrator1_adj_6558[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16353), .COUT(n16354), .S0(integrator1_71__N_960_adj_6573[12]), 
          .S1(integrator1_71__N_960_adj_6573[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_12 (.A0(mix_cosinewave[10]), .B0(integrator1_adj_6558[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[11]), .B1(integrator1_adj_6558[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16352), .COUT(n16353), .S0(integrator1_71__N_960_adj_6573[10]), 
          .S1(integrator1_71__N_960_adj_6573[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_10 (.A0(mix_cosinewave[8]), .B0(integrator1_adj_6558[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[9]), .B1(integrator1_adj_6558[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16351), .COUT(n16352), .S0(integrator1_71__N_960_adj_6573[8]), 
          .S1(integrator1_71__N_960_adj_6573[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_8 (.A0(mix_cosinewave[6]), .B0(integrator1_adj_6558[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[7]), .B1(integrator1_adj_6558[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16350), .COUT(n16351), .S0(integrator1_71__N_960_adj_6573[6]), 
          .S1(integrator1_71__N_960_adj_6573[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_6 (.A0(mix_cosinewave[4]), .B0(integrator1_adj_6558[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[5]), .B1(integrator1_adj_6558[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16349), .COUT(n16350), .S0(integrator1_71__N_960_adj_6573[4]), 
          .S1(integrator1_71__N_960_adj_6573[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_4 (.A0(mix_cosinewave[2]), .B0(integrator1_adj_6558[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[3]), .B1(integrator1_adj_6558[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16348), .COUT(n16349), .S0(integrator1_71__N_960_adj_6573[2]), 
          .S1(integrator1_71__N_960_adj_6573[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3522_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3522_add_4_2 (.A0(mix_cosinewave[0]), .B0(integrator1_adj_6558[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(mix_cosinewave[1]), .B1(integrator1_adj_6558[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16348), .S1(integrator1_71__N_960_adj_6573[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3522_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_3522_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3522_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3522_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_37 (.A0(integrator4_adj_6561[70]), .B0(cout_adj_6092), 
          .C0(n81_adj_6475), .D0(integrator5_adj_6562[70]), .A1(integrator4_adj_6561[71]), 
          .B1(cout_adj_6092), .C1(n78_adj_6474), .D1(integrator5_adj_6562[71]), 
          .CIN(n16345), .S0(integrator5_71__N_1248_adj_6577[70]), .S1(integrator5_71__N_1248_adj_6577[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_35 (.A0(integrator4_adj_6561[68]), .B0(cout_adj_6092), 
          .C0(n87_adj_6477), .D0(integrator5_adj_6562[68]), .A1(integrator4_adj_6561[69]), 
          .B1(cout_adj_6092), .C1(n84_adj_6476), .D1(integrator5_adj_6562[69]), 
          .CIN(n16344), .COUT(n16345), .S0(integrator5_71__N_1248_adj_6577[68]), 
          .S1(integrator5_71__N_1248_adj_6577[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_33 (.A0(integrator4_adj_6561[66]), .B0(cout_adj_6092), 
          .C0(n93_adj_6479), .D0(integrator5_adj_6562[66]), .A1(integrator4_adj_6561[67]), 
          .B1(cout_adj_6092), .C1(n90_adj_6478), .D1(integrator5_adj_6562[67]), 
          .CIN(n16343), .COUT(n16344), .S0(integrator5_71__N_1248_adj_6577[66]), 
          .S1(integrator5_71__N_1248_adj_6577[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_31 (.A0(integrator4_adj_6561[64]), .B0(cout_adj_6092), 
          .C0(n99_adj_6481), .D0(integrator5_adj_6562[64]), .A1(integrator4_adj_6561[65]), 
          .B1(cout_adj_6092), .C1(n96_adj_6480), .D1(integrator5_adj_6562[65]), 
          .CIN(n16342), .COUT(n16343), .S0(integrator5_71__N_1248_adj_6577[64]), 
          .S1(integrator5_71__N_1248_adj_6577[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_29 (.A0(integrator4_adj_6561[62]), .B0(cout_adj_6092), 
          .C0(n105_adj_6483), .D0(integrator5_adj_6562[62]), .A1(integrator4_adj_6561[63]), 
          .B1(cout_adj_6092), .C1(n102_adj_6482), .D1(integrator5_adj_6562[63]), 
          .CIN(n16341), .COUT(n16342), .S0(integrator5_71__N_1248_adj_6577[62]), 
          .S1(integrator5_71__N_1248_adj_6577[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_27 (.A0(integrator4_adj_6561[60]), .B0(cout_adj_6092), 
          .C0(n111_adj_6485), .D0(integrator5_adj_6562[60]), .A1(integrator4_adj_6561[61]), 
          .B1(cout_adj_6092), .C1(n108_adj_6484), .D1(integrator5_adj_6562[61]), 
          .CIN(n16340), .COUT(n16341), .S0(integrator5_71__N_1248_adj_6577[60]), 
          .S1(integrator5_71__N_1248_adj_6577[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_25 (.A0(integrator4_adj_6561[58]), .B0(cout_adj_6092), 
          .C0(n117_adj_6487), .D0(integrator5_adj_6562[58]), .A1(integrator4_adj_6561[59]), 
          .B1(cout_adj_6092), .C1(n114_adj_6486), .D1(integrator5_adj_6562[59]), 
          .CIN(n16339), .COUT(n16340), .S0(integrator5_71__N_1248_adj_6577[58]), 
          .S1(integrator5_71__N_1248_adj_6577[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_23 (.A0(integrator4_adj_6561[56]), .B0(cout_adj_6092), 
          .C0(n123_adj_6489), .D0(integrator5_adj_6562[56]), .A1(integrator4_adj_6561[57]), 
          .B1(cout_adj_6092), .C1(n120_adj_6488), .D1(integrator5_adj_6562[57]), 
          .CIN(n16338), .COUT(n16339), .S0(integrator5_71__N_1248_adj_6577[56]), 
          .S1(integrator5_71__N_1248_adj_6577[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_21 (.A0(integrator4_adj_6561[54]), .B0(cout_adj_6092), 
          .C0(n129_adj_6491), .D0(integrator5_adj_6562[54]), .A1(integrator4_adj_6561[55]), 
          .B1(cout_adj_6092), .C1(n126_adj_6490), .D1(integrator5_adj_6562[55]), 
          .CIN(n16337), .COUT(n16338), .S0(integrator5_71__N_1248_adj_6577[54]), 
          .S1(integrator5_71__N_1248_adj_6577[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_19 (.A0(integrator4_adj_6561[52]), .B0(cout_adj_6092), 
          .C0(n135_adj_6493), .D0(integrator5_adj_6562[52]), .A1(integrator4_adj_6561[53]), 
          .B1(cout_adj_6092), .C1(n132_adj_6492), .D1(integrator5_adj_6562[53]), 
          .CIN(n16336), .COUT(n16337), .S0(integrator5_71__N_1248_adj_6577[52]), 
          .S1(integrator5_71__N_1248_adj_6577[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_17 (.A0(integrator4_adj_6561[50]), .B0(cout_adj_6092), 
          .C0(n141_adj_6495), .D0(integrator5_adj_6562[50]), .A1(integrator4_adj_6561[51]), 
          .B1(cout_adj_6092), .C1(n138_adj_6494), .D1(integrator5_adj_6562[51]), 
          .CIN(n16335), .COUT(n16336), .S0(integrator5_71__N_1248_adj_6577[50]), 
          .S1(integrator5_71__N_1248_adj_6577[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_15 (.A0(integrator4_adj_6561[48]), .B0(cout_adj_6092), 
          .C0(n147_adj_6497), .D0(integrator5_adj_6562[48]), .A1(integrator4_adj_6561[49]), 
          .B1(cout_adj_6092), .C1(n144_adj_6496), .D1(integrator5_adj_6562[49]), 
          .CIN(n16334), .COUT(n16335), .S0(integrator5_71__N_1248_adj_6577[48]), 
          .S1(integrator5_71__N_1248_adj_6577[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_13 (.A0(integrator4_adj_6561[46]), .B0(cout_adj_6092), 
          .C0(n153_adj_6499), .D0(integrator5_adj_6562[46]), .A1(integrator4_adj_6561[47]), 
          .B1(cout_adj_6092), .C1(n150_adj_6498), .D1(integrator5_adj_6562[47]), 
          .CIN(n16333), .COUT(n16334), .S0(integrator5_71__N_1248_adj_6577[46]), 
          .S1(integrator5_71__N_1248_adj_6577[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_11 (.A0(integrator4_adj_6561[44]), .B0(cout_adj_6092), 
          .C0(n159_adj_6501), .D0(integrator5_adj_6562[44]), .A1(integrator4_adj_6561[45]), 
          .B1(cout_adj_6092), .C1(n156_adj_6500), .D1(integrator5_adj_6562[45]), 
          .CIN(n16332), .COUT(n16333), .S0(integrator5_71__N_1248_adj_6577[44]), 
          .S1(integrator5_71__N_1248_adj_6577[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_9 (.A0(integrator4_adj_6561[42]), .B0(cout_adj_6092), 
          .C0(n165_adj_6503), .D0(integrator5_adj_6562[42]), .A1(integrator4_adj_6561[43]), 
          .B1(cout_adj_6092), .C1(n162_adj_6502), .D1(integrator5_adj_6562[43]), 
          .CIN(n16331), .COUT(n16332), .S0(integrator5_71__N_1248_adj_6577[42]), 
          .S1(integrator5_71__N_1248_adj_6577[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_7 (.A0(integrator4_adj_6561[40]), .B0(cout_adj_6092), 
          .C0(n171_adj_6505), .D0(integrator5_adj_6562[40]), .A1(integrator4_adj_6561[41]), 
          .B1(cout_adj_6092), .C1(n168_adj_6504), .D1(integrator5_adj_6562[41]), 
          .CIN(n16330), .COUT(n16331), .S0(integrator5_71__N_1248_adj_6577[40]), 
          .S1(integrator5_71__N_1248_adj_6577[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_5 (.A0(integrator4_adj_6561[38]), .B0(cout_adj_6092), 
          .C0(n177_adj_6507), .D0(integrator5_adj_6562[38]), .A1(integrator4_adj_6561[39]), 
          .B1(cout_adj_6092), .C1(n174_adj_6506), .D1(integrator5_adj_6562[39]), 
          .CIN(n16329), .COUT(n16330), .S0(integrator5_71__N_1248_adj_6577[38]), 
          .S1(integrator5_71__N_1248_adj_6577[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_3 (.A0(integrator4_adj_6561[36]), .B0(cout_adj_6092), 
          .C0(n183_adj_6509), .D0(integrator5_adj_6562[36]), .A1(integrator4_adj_6561[37]), 
          .B1(cout_adj_6092), .C1(n180_adj_6508), .D1(integrator5_adj_6562[37]), 
          .CIN(n16328), .COUT(n16329), .S0(integrator5_71__N_1248_adj_6577[36]), 
          .S1(integrator5_71__N_1248_adj_6577[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3660_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3660_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_20 (.A0(comb_d9_adj_6570[17]), .B0(comb9_adj_6569[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[18]), .B1(comb9_adj_6569[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17706), .COUT(n17707));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_18 (.A0(comb_d9_adj_6570[15]), .B0(comb9_adj_6569[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[16]), .B1(comb9_adj_6569[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17705), .COUT(n17706));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_9 (.A0(comb6_adj_6563[42]), .B0(cout_adj_5627), 
          .C0(n165_adj_5754), .D0(n31_adj_5521), .A1(comb6_adj_6563[43]), 
          .B1(cout_adj_5627), .C1(n162_adj_5753), .D1(n30_adj_5520), .CIN(n17215), 
          .COUT(n17216), .S0(comb7_71__N_2065_adj_6590[42]), .S1(comb7_71__N_2065_adj_6590[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_16 (.A0(comb_d9_adj_6570[13]), .B0(comb9_adj_6569[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[14]), .B1(comb9_adj_6569[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17704), .COUT(n17705));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_14 (.A0(comb_d9_adj_6570[11]), .B0(comb9_adj_6569[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[12]), .B1(comb9_adj_6569[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17703), .COUT(n17704));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_12 (.A0(comb_d9_adj_6570[9]), .B0(comb9_adj_6569[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[10]), .B1(comb9_adj_6569[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17702), .COUT(n17703));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_7 (.A0(comb6_adj_6563[40]), .B0(cout_adj_5627), 
          .C0(n171_adj_5756), .D0(n33_adj_5523), .A1(comb6_adj_6563[41]), 
          .B1(cout_adj_5627), .C1(n168_adj_5755), .D1(n32_adj_5522), .CIN(n17214), 
          .COUT(n17215), .S0(comb7_71__N_2065_adj_6590[40]), .S1(comb7_71__N_2065_adj_6590[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_5 (.A0(comb6_adj_6563[38]), .B0(cout_adj_5627), 
          .C0(n177_adj_5758), .D0(n35_adj_5525), .A1(comb6_adj_6563[39]), 
          .B1(cout_adj_5627), .C1(n174_adj_5757), .D1(n34_adj_5524), .CIN(n17213), 
          .COUT(n17214), .S0(comb7_71__N_2065_adj_6590[38]), .S1(comb7_71__N_2065_adj_6590[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_10 (.A0(comb_d9_adj_6570[7]), .B0(comb9_adj_6569[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[8]), .B1(comb9_adj_6569[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17701), .COUT(n17702));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3660_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_6092), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16328));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3660_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3660_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3660_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3660_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_38 (.A0(comb_d6_adj_6564[35]), .B0(comb6_adj_6563[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16324), .S0(comb7_71__N_2065_adj_6590[35]), 
          .S1(cout_adj_5627));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3675_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_36 (.A0(comb_d6_adj_6564[33]), .B0(comb6_adj_6563[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[34]), .B1(comb6_adj_6563[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16323), .COUT(n16324), .S0(comb7_71__N_2065_adj_6590[33]), 
          .S1(comb7_71__N_2065_adj_6590[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_34 (.A0(comb_d6_adj_6564[31]), .B0(comb6_adj_6563[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[32]), .B1(comb6_adj_6563[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16322), .COUT(n16323), .S0(comb7_71__N_2065_adj_6590[31]), 
          .S1(comb7_71__N_2065_adj_6590[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_32 (.A0(comb_d6_adj_6564[29]), .B0(comb6_adj_6563[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[30]), .B1(comb6_adj_6563[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16321), .COUT(n16322), .S0(comb7_71__N_2065_adj_6590[29]), 
          .S1(comb7_71__N_2065_adj_6590[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_30 (.A0(comb_d6_adj_6564[27]), .B0(comb6_adj_6563[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[28]), .B1(comb6_adj_6563[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16320), .COUT(n16321), .S0(comb7_71__N_2065_adj_6590[27]), 
          .S1(comb7_71__N_2065_adj_6590[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_28 (.A0(comb_d6_adj_6564[25]), .B0(comb6_adj_6563[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[26]), .B1(comb6_adj_6563[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16319), .COUT(n16320), .S0(comb7_71__N_2065_adj_6590[25]), 
          .S1(comb7_71__N_2065_adj_6590[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_26 (.A0(comb_d6_adj_6564[23]), .B0(comb6_adj_6563[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[24]), .B1(comb6_adj_6563[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16318), .COUT(n16319), .S0(comb7_71__N_2065_adj_6590[23]), 
          .S1(comb7_71__N_2065_adj_6590[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_24 (.A0(comb_d6_adj_6564[21]), .B0(comb6_adj_6563[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[22]), .B1(comb6_adj_6563[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16317), .COUT(n16318), .S0(comb7_71__N_2065_adj_6590[21]), 
          .S1(comb7_71__N_2065_adj_6590[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_22 (.A0(comb_d6_adj_6564[19]), .B0(comb6_adj_6563[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[20]), .B1(comb6_adj_6563[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16316), .COUT(n16317), .S0(comb7_71__N_2065_adj_6590[19]), 
          .S1(comb7_71__N_2065_adj_6590[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_20 (.A0(comb_d6_adj_6564[17]), .B0(comb6_adj_6563[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[18]), .B1(comb6_adj_6563[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16315), .COUT(n16316), .S0(comb7_71__N_2065_adj_6590[17]), 
          .S1(comb7_71__N_2065_adj_6590[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_18 (.A0(comb_d6_adj_6564[15]), .B0(comb6_adj_6563[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[16]), .B1(comb6_adj_6563[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16314), .COUT(n16315), .S0(comb7_71__N_2065_adj_6590[15]), 
          .S1(comb7_71__N_2065_adj_6590[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_16 (.A0(comb_d6_adj_6564[13]), .B0(comb6_adj_6563[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[14]), .B1(comb6_adj_6563[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16313), .COUT(n16314), .S0(comb7_71__N_2065_adj_6590[13]), 
          .S1(comb7_71__N_2065_adj_6590[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_14 (.A0(comb_d6_adj_6564[11]), .B0(comb6_adj_6563[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[12]), .B1(comb6_adj_6563[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16312), .COUT(n16313), .S0(comb7_71__N_2065_adj_6590[11]), 
          .S1(comb7_71__N_2065_adj_6590[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_12 (.A0(comb_d6_adj_6564[9]), .B0(comb6_adj_6563[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[10]), .B1(comb6_adj_6563[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16311), .COUT(n16312), .S0(comb7_71__N_2065_adj_6590[9]), 
          .S1(comb7_71__N_2065_adj_6590[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_10 (.A0(comb_d6_adj_6564[7]), .B0(comb6_adj_6563[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[8]), .B1(comb6_adj_6563[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16310), .COUT(n16311), .S0(comb7_71__N_2065_adj_6590[7]), 
          .S1(comb7_71__N_2065_adj_6590[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_8 (.A0(comb_d6_adj_6564[5]), .B0(comb6_adj_6563[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[6]), .B1(comb6_adj_6563[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16309), .COUT(n16310), .S0(comb7_71__N_2065_adj_6590[5]), 
          .S1(comb7_71__N_2065_adj_6590[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_6 (.A0(comb_d6_adj_6564[3]), .B0(comb6_adj_6563[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[4]), .B1(comb6_adj_6563[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16308), .COUT(n16309), .S0(comb7_71__N_2065_adj_6590[3]), 
          .S1(comb7_71__N_2065_adj_6590[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_4 (.A0(comb_d6_adj_6564[1]), .B0(comb6_adj_6563[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[2]), .B1(comb6_adj_6563[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16307), .COUT(n16308), .S0(comb7_71__N_2065_adj_6590[1]), 
          .S1(comb7_71__N_2065_adj_6590[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3675_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3675_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6_adj_6564[0]), .B1(comb6_adj_6563[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16307), .S1(comb7_71__N_2065_adj_6590[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3675_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3675_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3675_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3675_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_37 (.A0(integrator1[70]), .B0(cout_adj_6289), 
          .C0(n81_adj_6202), .D0(mix_sinewave[11]), .A1(integrator1[71]), 
          .B1(cout_adj_6289), .C1(n78_adj_6201), .D1(mix_sinewave[11]), 
          .CIN(n16305), .S0(integrator1_71__N_960[70]), .S1(integrator1_71__N_960[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_35 (.A0(integrator1[68]), .B0(cout_adj_6289), 
          .C0(n87_adj_6204), .D0(mix_sinewave[11]), .A1(integrator1[69]), 
          .B1(cout_adj_6289), .C1(n84_adj_6203), .D1(mix_sinewave[11]), 
          .CIN(n16304), .COUT(n16305), .S0(integrator1_71__N_960[68]), 
          .S1(integrator1_71__N_960[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_33 (.A0(integrator1[66]), .B0(cout_adj_6289), 
          .C0(n93_adj_6206), .D0(mix_sinewave[11]), .A1(integrator1[67]), 
          .B1(cout_adj_6289), .C1(n90_adj_6205), .D1(mix_sinewave[11]), 
          .CIN(n16303), .COUT(n16304), .S0(integrator1_71__N_960[66]), 
          .S1(integrator1_71__N_960[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_31 (.A0(integrator1[64]), .B0(cout_adj_6289), 
          .C0(n99_adj_6208), .D0(mix_sinewave[11]), .A1(integrator1[65]), 
          .B1(cout_adj_6289), .C1(n96_adj_6207), .D1(mix_sinewave[11]), 
          .CIN(n16302), .COUT(n16303), .S0(integrator1_71__N_960[64]), 
          .S1(integrator1_71__N_960[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_29 (.A0(integrator1[62]), .B0(cout_adj_6289), 
          .C0(n105_adj_6210), .D0(mix_sinewave[11]), .A1(integrator1[63]), 
          .B1(cout_adj_6289), .C1(n102_adj_6209), .D1(mix_sinewave[11]), 
          .CIN(n16301), .COUT(n16302), .S0(integrator1_71__N_960[62]), 
          .S1(integrator1_71__N_960[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_27 (.A0(integrator1[60]), .B0(cout_adj_6289), 
          .C0(n111_adj_6212), .D0(mix_sinewave[11]), .A1(integrator1[61]), 
          .B1(cout_adj_6289), .C1(n108_adj_6211), .D1(mix_sinewave[11]), 
          .CIN(n16300), .COUT(n16301), .S0(integrator1_71__N_960[60]), 
          .S1(integrator1_71__N_960[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_25 (.A0(integrator1[58]), .B0(cout_adj_6289), 
          .C0(n117_adj_6214), .D0(mix_sinewave[11]), .A1(integrator1[59]), 
          .B1(cout_adj_6289), .C1(n114_adj_6213), .D1(mix_sinewave[11]), 
          .CIN(n16299), .COUT(n16300), .S0(integrator1_71__N_960[58]), 
          .S1(integrator1_71__N_960[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_23 (.A0(integrator1[56]), .B0(cout_adj_6289), 
          .C0(n123_adj_6216), .D0(mix_sinewave[11]), .A1(integrator1[57]), 
          .B1(cout_adj_6289), .C1(n120_adj_6215), .D1(mix_sinewave[11]), 
          .CIN(n16298), .COUT(n16299), .S0(integrator1_71__N_960[56]), 
          .S1(integrator1_71__N_960[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_21 (.A0(integrator1[54]), .B0(cout_adj_6289), 
          .C0(n129_adj_6218), .D0(mix_sinewave[11]), .A1(integrator1[55]), 
          .B1(cout_adj_6289), .C1(n126_adj_6217), .D1(mix_sinewave[11]), 
          .CIN(n16297), .COUT(n16298), .S0(integrator1_71__N_960[54]), 
          .S1(integrator1_71__N_960[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_19 (.A0(integrator1[52]), .B0(cout_adj_6289), 
          .C0(n135_adj_6220), .D0(mix_sinewave[11]), .A1(integrator1[53]), 
          .B1(cout_adj_6289), .C1(n132_adj_6219), .D1(mix_sinewave[11]), 
          .CIN(n16296), .COUT(n16297), .S0(integrator1_71__N_960[52]), 
          .S1(integrator1_71__N_960[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_17 (.A0(integrator1[50]), .B0(cout_adj_6289), 
          .C0(n141_adj_6222), .D0(mix_sinewave[11]), .A1(integrator1[51]), 
          .B1(cout_adj_6289), .C1(n138_adj_6221), .D1(mix_sinewave[11]), 
          .CIN(n16295), .COUT(n16296), .S0(integrator1_71__N_960[50]), 
          .S1(integrator1_71__N_960[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_15 (.A0(integrator1[48]), .B0(cout_adj_6289), 
          .C0(n147_adj_6224), .D0(mix_sinewave[11]), .A1(integrator1[49]), 
          .B1(cout_adj_6289), .C1(n144_adj_6223), .D1(mix_sinewave[11]), 
          .CIN(n16294), .COUT(n16295), .S0(integrator1_71__N_960[48]), 
          .S1(integrator1_71__N_960[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_13 (.A0(integrator1[46]), .B0(cout_adj_6289), 
          .C0(n153_adj_6226), .D0(mix_sinewave[11]), .A1(integrator1[47]), 
          .B1(cout_adj_6289), .C1(n150_adj_6225), .D1(mix_sinewave[11]), 
          .CIN(n16293), .COUT(n16294), .S0(integrator1_71__N_960[46]), 
          .S1(integrator1_71__N_960[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_13.INJECT1_1 = "NO";
    LUT4 i5021_2_lut (.A(phase_increment_1__63__N_17[6]), .B(led_0_6), .Z(n4097)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i5021_2_lut.init = 16'heeee;
    LUT4 i5022_2_lut (.A(phase_increment_1__63__N_21[6]), .B(rx_byte[0]), 
         .Z(n4112)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i5022_2_lut.init = 16'heeee;
    FD1S3AX square_sum_e3__i2 (.D(n123_adj_5601), .CK(cic_sine_clk), .Q(square_sum[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i2.GSR = "ENABLED";
    CCU2C _add_1_3648_add_4_3 (.A0(comb6_adj_6563[36]), .B0(cout_adj_5627), 
          .C0(n183_adj_5760), .D0(n37_adj_5527), .A1(comb6_adj_6563[37]), 
          .B1(cout_adj_5627), .C1(n180_adj_5759), .D1(n36_adj_5526), .CIN(n17212), 
          .COUT(n17213), .S0(comb7_71__N_2065_adj_6590[36]), .S1(comb7_71__N_2065_adj_6590[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3648_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3648_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3648_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5627), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17212));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3648_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3648_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3648_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3648_add_4_1.INJECT1_1 = "NO";
    PFUMX mux_1393_i1 (.BLUT(n2613), .ALUT(n2619), .C0(n19302), .Z(n2622));
    CCU2C _add_1_3651_add_4_37 (.A0(comb7_adj_6565[70]), .B0(cout_adj_5840), 
          .C0(n81_adj_5676), .D0(n3_adj_5529), .A1(comb7_adj_6565[71]), 
          .B1(cout_adj_5840), .C1(n78_adj_5675), .D1(n2_adj_5528), .CIN(n17207), 
          .S0(comb8_71__N_2137_adj_6591[70]), .S1(comb8_71__N_2137_adj_6591[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_35 (.A0(comb7_adj_6565[68]), .B0(cout_adj_5840), 
          .C0(n87_adj_5678), .D0(n5_adj_5531), .A1(comb7_adj_6565[69]), 
          .B1(cout_adj_5840), .C1(n84_adj_5677), .D1(n4_adj_5530), .CIN(n17206), 
          .COUT(n17207), .S0(comb8_71__N_2137_adj_6591[68]), .S1(comb8_71__N_2137_adj_6591[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_33 (.A0(comb7_adj_6565[66]), .B0(cout_adj_5840), 
          .C0(n93_adj_5680), .D0(n7_adj_5533), .A1(comb7_adj_6565[67]), 
          .B1(cout_adj_5840), .C1(n90_adj_5679), .D1(n6_adj_5532), .CIN(n17205), 
          .COUT(n17206), .S0(comb8_71__N_2137_adj_6591[66]), .S1(comb8_71__N_2137_adj_6591[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_31 (.A0(comb7_adj_6565[64]), .B0(cout_adj_5840), 
          .C0(n99_adj_5682), .D0(n9_adj_5535), .A1(comb7_adj_6565[65]), 
          .B1(cout_adj_5840), .C1(n96_adj_5681), .D1(n8_adj_5534), .CIN(n17204), 
          .COUT(n17205), .S0(comb8_71__N_2137_adj_6591[64]), .S1(comb8_71__N_2137_adj_6591[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_29 (.A0(comb7_adj_6565[62]), .B0(cout_adj_5840), 
          .C0(n105_adj_5684), .D0(n11_adj_5537), .A1(comb7_adj_6565[63]), 
          .B1(cout_adj_5840), .C1(n102_adj_5683), .D1(n10_adj_5536), .CIN(n17203), 
          .COUT(n17204), .S0(comb8_71__N_2137_adj_6591[62]), .S1(comb8_71__N_2137_adj_6591[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_27 (.A0(comb7_adj_6565[60]), .B0(cout_adj_5840), 
          .C0(n111_adj_5686), .D0(n13_adj_5539), .A1(comb7_adj_6565[61]), 
          .B1(cout_adj_5840), .C1(n108_adj_5685), .D1(n12_adj_5538), .CIN(n17202), 
          .COUT(n17203), .S0(comb8_71__N_2137_adj_6591[60]), .S1(comb8_71__N_2137_adj_6591[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_25 (.A0(comb7_adj_6565[58]), .B0(cout_adj_5840), 
          .C0(n117_adj_5688), .D0(n15_adj_5541), .A1(comb7_adj_6565[59]), 
          .B1(cout_adj_5840), .C1(n114_adj_5687), .D1(n14_adj_5540), .CIN(n17201), 
          .COUT(n17202), .S0(comb8_71__N_2137_adj_6591[58]), .S1(comb8_71__N_2137_adj_6591[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_23 (.A0(comb7_adj_6565[56]), .B0(cout_adj_5840), 
          .C0(n123_adj_5690), .D0(n17_adj_5543), .A1(comb7_adj_6565[57]), 
          .B1(cout_adj_5840), .C1(n120_adj_5689), .D1(n16_adj_5542), .CIN(n17200), 
          .COUT(n17201), .S0(comb8_71__N_2137_adj_6591[56]), .S1(comb8_71__N_2137_adj_6591[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_21 (.A0(comb7_adj_6565[54]), .B0(cout_adj_5840), 
          .C0(n129_adj_5692), .D0(n19_adj_5545), .A1(comb7_adj_6565[55]), 
          .B1(cout_adj_5840), .C1(n126_adj_5691), .D1(n18_adj_5544), .CIN(n17199), 
          .COUT(n17200), .S0(comb8_71__N_2137_adj_6591[54]), .S1(comb8_71__N_2137_adj_6591[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_19 (.A0(comb7_adj_6565[52]), .B0(cout_adj_5840), 
          .C0(n135_adj_5694), .D0(n21_adj_5547), .A1(comb7_adj_6565[53]), 
          .B1(cout_adj_5840), .C1(n132_adj_5693), .D1(n20_adj_5546), .CIN(n17198), 
          .COUT(n17199), .S0(comb8_71__N_2137_adj_6591[52]), .S1(comb8_71__N_2137_adj_6591[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_17 (.A0(comb7_adj_6565[50]), .B0(cout_adj_5840), 
          .C0(n141_adj_5696), .D0(n23_adj_5549), .A1(comb7_adj_6565[51]), 
          .B1(cout_adj_5840), .C1(n138_adj_5695), .D1(n22_adj_5548), .CIN(n17197), 
          .COUT(n17198), .S0(comb8_71__N_2137_adj_6591[50]), .S1(comb8_71__N_2137_adj_6591[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_11 (.A0(integrator1[44]), .B0(cout_adj_6289), 
          .C0(n159_adj_6228), .D0(mix_sinewave[11]), .A1(integrator1[45]), 
          .B1(cout_adj_6289), .C1(n156_adj_6227), .D1(mix_sinewave[11]), 
          .CIN(n16292), .COUT(n16293), .S0(integrator1_71__N_960[44]), 
          .S1(integrator1_71__N_960[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_9 (.A0(integrator1[42]), .B0(cout_adj_6289), 
          .C0(n165_adj_6230), .D0(mix_sinewave[11]), .A1(integrator1[43]), 
          .B1(cout_adj_6289), .C1(n162_adj_6229), .D1(mix_sinewave[11]), 
          .CIN(n16291), .COUT(n16292), .S0(integrator1_71__N_960[42]), 
          .S1(integrator1_71__N_960[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_7 (.A0(integrator1[40]), .B0(cout_adj_6289), 
          .C0(n171_adj_6232), .D0(mix_sinewave[11]), .A1(integrator1[41]), 
          .B1(cout_adj_6289), .C1(n168_adj_6231), .D1(mix_sinewave[11]), 
          .CIN(n16290), .COUT(n16291), .S0(integrator1_71__N_960[40]), 
          .S1(integrator1_71__N_960[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_5 (.A0(integrator1[38]), .B0(cout_adj_6289), 
          .C0(n177_adj_6234), .D0(mix_sinewave[11]), .A1(integrator1[39]), 
          .B1(cout_adj_6289), .C1(n174_adj_6233), .D1(mix_sinewave[11]), 
          .CIN(n16289), .COUT(n16290), .S0(integrator1_71__N_960[38]), 
          .S1(integrator1_71__N_960[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_3 (.A0(integrator1[36]), .B0(cout_adj_6289), 
          .C0(n183_adj_6236), .D0(mix_sinewave[11]), .A1(integrator1[37]), 
          .B1(cout_adj_6289), .C1(n180_adj_6235), .D1(mix_sinewave[11]), 
          .CIN(n16288), .COUT(n16289), .S0(integrator1_71__N_960[36]), 
          .S1(integrator1_71__N_960[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3552_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3552_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3552_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_6289), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16288));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(73[20:41])
    defparam _add_1_3552_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3552_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3552_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3552_add_4_1.INJECT1_1 = "NO";
    LUT4 rx_byte_2__bdd_3_lut_8610 (.A(rx_byte[2]), .B(n19575), .C(rx_byte[3]), 
         .Z(n19576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam rx_byte_2__bdd_3_lut_8610.init = 16'hcaca;
    PFUMX mux_2163_i1 (.BLUT(n3647), .ALUT(n3653), .C0(n19301), .Z(n3656));
    CCU2C _add_1_3663_add_4_37 (.A0(integrator3_adj_6560[70]), .B0(cout_adj_6091), 
          .C0(n81_adj_6425), .D0(integrator4_adj_6561[70]), .A1(integrator3_adj_6560[71]), 
          .B1(cout_adj_6091), .C1(n78_adj_6424), .D1(integrator4_adj_6561[71]), 
          .CIN(n16283), .S0(integrator4_71__N_1176_adj_6576[70]), .S1(integrator4_71__N_1176_adj_6576[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_35 (.A0(integrator3_adj_6560[68]), .B0(cout_adj_6091), 
          .C0(n87_adj_6427), .D0(integrator4_adj_6561[68]), .A1(integrator3_adj_6560[69]), 
          .B1(cout_adj_6091), .C1(n84_adj_6426), .D1(integrator4_adj_6561[69]), 
          .CIN(n16282), .COUT(n16283), .S0(integrator4_71__N_1176_adj_6576[68]), 
          .S1(integrator4_71__N_1176_adj_6576[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_33 (.A0(integrator3_adj_6560[66]), .B0(cout_adj_6091), 
          .C0(n93_adj_6429), .D0(integrator4_adj_6561[66]), .A1(integrator3_adj_6560[67]), 
          .B1(cout_adj_6091), .C1(n90_adj_6428), .D1(integrator4_adj_6561[67]), 
          .CIN(n16281), .COUT(n16282), .S0(integrator4_71__N_1176_adj_6576[66]), 
          .S1(integrator4_71__N_1176_adj_6576[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_31 (.A0(integrator3_adj_6560[64]), .B0(cout_adj_6091), 
          .C0(n99_adj_6431), .D0(integrator4_adj_6561[64]), .A1(integrator3_adj_6560[65]), 
          .B1(cout_adj_6091), .C1(n96_adj_6430), .D1(integrator4_adj_6561[65]), 
          .CIN(n16280), .COUT(n16281), .S0(integrator4_71__N_1176_adj_6576[64]), 
          .S1(integrator4_71__N_1176_adj_6576[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_29 (.A0(integrator3_adj_6560[62]), .B0(cout_adj_6091), 
          .C0(n105_adj_6433), .D0(integrator4_adj_6561[62]), .A1(integrator3_adj_6560[63]), 
          .B1(cout_adj_6091), .C1(n102_adj_6432), .D1(integrator4_adj_6561[63]), 
          .CIN(n16279), .COUT(n16280), .S0(integrator4_71__N_1176_adj_6576[62]), 
          .S1(integrator4_71__N_1176_adj_6576[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_27 (.A0(integrator3_adj_6560[60]), .B0(cout_adj_6091), 
          .C0(n111_adj_6435), .D0(integrator4_adj_6561[60]), .A1(integrator3_adj_6560[61]), 
          .B1(cout_adj_6091), .C1(n108_adj_6434), .D1(integrator4_adj_6561[61]), 
          .CIN(n16278), .COUT(n16279), .S0(integrator4_71__N_1176_adj_6576[60]), 
          .S1(integrator4_71__N_1176_adj_6576[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_25 (.A0(integrator3_adj_6560[58]), .B0(cout_adj_6091), 
          .C0(n117_adj_6437), .D0(integrator4_adj_6561[58]), .A1(integrator3_adj_6560[59]), 
          .B1(cout_adj_6091), .C1(n114_adj_6436), .D1(integrator4_adj_6561[59]), 
          .CIN(n16277), .COUT(n16278), .S0(integrator4_71__N_1176_adj_6576[58]), 
          .S1(integrator4_71__N_1176_adj_6576[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_23 (.A0(integrator3_adj_6560[56]), .B0(cout_adj_6091), 
          .C0(n123_adj_6439), .D0(integrator4_adj_6561[56]), .A1(integrator3_adj_6560[57]), 
          .B1(cout_adj_6091), .C1(n120_adj_6438), .D1(integrator4_adj_6561[57]), 
          .CIN(n16276), .COUT(n16277), .S0(integrator4_71__N_1176_adj_6576[56]), 
          .S1(integrator4_71__N_1176_adj_6576[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_21 (.A0(integrator3_adj_6560[54]), .B0(cout_adj_6091), 
          .C0(n129_adj_6441), .D0(integrator4_adj_6561[54]), .A1(integrator3_adj_6560[55]), 
          .B1(cout_adj_6091), .C1(n126_adj_6440), .D1(integrator4_adj_6561[55]), 
          .CIN(n16275), .COUT(n16276), .S0(integrator4_71__N_1176_adj_6576[54]), 
          .S1(integrator4_71__N_1176_adj_6576[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_19 (.A0(integrator3_adj_6560[52]), .B0(cout_adj_6091), 
          .C0(n135_adj_6443), .D0(integrator4_adj_6561[52]), .A1(integrator3_adj_6560[53]), 
          .B1(cout_adj_6091), .C1(n132_adj_6442), .D1(integrator4_adj_6561[53]), 
          .CIN(n16274), .COUT(n16275), .S0(integrator4_71__N_1176_adj_6576[52]), 
          .S1(integrator4_71__N_1176_adj_6576[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_17 (.A0(integrator3_adj_6560[50]), .B0(cout_adj_6091), 
          .C0(n141_adj_6445), .D0(integrator4_adj_6561[50]), .A1(integrator3_adj_6560[51]), 
          .B1(cout_adj_6091), .C1(n138_adj_6444), .D1(integrator4_adj_6561[51]), 
          .CIN(n16273), .COUT(n16274), .S0(integrator4_71__N_1176_adj_6576[50]), 
          .S1(integrator4_71__N_1176_adj_6576[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_15 (.A0(integrator3_adj_6560[48]), .B0(cout_adj_6091), 
          .C0(n147_adj_6447), .D0(integrator4_adj_6561[48]), .A1(integrator3_adj_6560[49]), 
          .B1(cout_adj_6091), .C1(n144_adj_6446), .D1(integrator4_adj_6561[49]), 
          .CIN(n16272), .COUT(n16273), .S0(integrator4_71__N_1176_adj_6576[48]), 
          .S1(integrator4_71__N_1176_adj_6576[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_13 (.A0(integrator3_adj_6560[46]), .B0(cout_adj_6091), 
          .C0(n153_adj_6449), .D0(integrator4_adj_6561[46]), .A1(integrator3_adj_6560[47]), 
          .B1(cout_adj_6091), .C1(n150_adj_6448), .D1(integrator4_adj_6561[47]), 
          .CIN(n16271), .COUT(n16272), .S0(integrator4_71__N_1176_adj_6576[46]), 
          .S1(integrator4_71__N_1176_adj_6576[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_11 (.A0(integrator3_adj_6560[44]), .B0(cout_adj_6091), 
          .C0(n159_adj_6451), .D0(integrator4_adj_6561[44]), .A1(integrator3_adj_6560[45]), 
          .B1(cout_adj_6091), .C1(n156_adj_6450), .D1(integrator4_adj_6561[45]), 
          .CIN(n16270), .COUT(n16271), .S0(integrator4_71__N_1176_adj_6576[44]), 
          .S1(integrator4_71__N_1176_adj_6576[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_9 (.A0(integrator3_adj_6560[42]), .B0(cout_adj_6091), 
          .C0(n165_adj_6453), .D0(integrator4_adj_6561[42]), .A1(integrator3_adj_6560[43]), 
          .B1(cout_adj_6091), .C1(n162_adj_6452), .D1(integrator4_adj_6561[43]), 
          .CIN(n16269), .COUT(n16270), .S0(integrator4_71__N_1176_adj_6576[42]), 
          .S1(integrator4_71__N_1176_adj_6576[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_7 (.A0(integrator3_adj_6560[40]), .B0(cout_adj_6091), 
          .C0(n171_adj_6455), .D0(integrator4_adj_6561[40]), .A1(integrator3_adj_6560[41]), 
          .B1(cout_adj_6091), .C1(n168_adj_6454), .D1(integrator4_adj_6561[41]), 
          .CIN(n16268), .COUT(n16269), .S0(integrator4_71__N_1176_adj_6576[40]), 
          .S1(integrator4_71__N_1176_adj_6576[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_5 (.A0(integrator3_adj_6560[38]), .B0(cout_adj_6091), 
          .C0(n177_adj_6457), .D0(integrator4_adj_6561[38]), .A1(integrator3_adj_6560[39]), 
          .B1(cout_adj_6091), .C1(n174_adj_6456), .D1(integrator4_adj_6561[39]), 
          .CIN(n16267), .COUT(n16268), .S0(integrator4_71__N_1176_adj_6576[38]), 
          .S1(integrator4_71__N_1176_adj_6576[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_3 (.A0(integrator3_adj_6560[36]), .B0(cout_adj_6091), 
          .C0(n183_adj_6459), .D0(integrator4_adj_6561[36]), .A1(integrator3_adj_6560[37]), 
          .B1(cout_adj_6091), .C1(n180_adj_6458), .D1(integrator4_adj_6561[37]), 
          .CIN(n16266), .COUT(n16267), .S0(integrator4_71__N_1176_adj_6576[36]), 
          .S1(integrator4_71__N_1176_adj_6576[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3663_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3663_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3663_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_6091), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16266));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3663_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3663_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3663_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3663_add_4_1.INJECT1_1 = "NO";
    LUT4 n3998_bdd_3_lut_8464 (.A(n3998), .B(rx_byte[2]), .C(rx_byte[3]), 
         .Z(n19443)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n3998_bdd_3_lut_8464.init = 16'hacac;
    LUT4 n3998_bdd_3_lut (.A(phase_increment_1__63__N_19[8]), .B(phase_increment_1__63__N_20[8]), 
         .C(rx_byte[0]), .Z(n19444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3998_bdd_3_lut.init = 16'hcaca;
    CCU2C _add_1_3666_add_4_37 (.A0(integrator2_adj_6559[70]), .B0(cout), 
          .C0(n81_adj_6389), .D0(integrator3_adj_6560[70]), .A1(integrator2_adj_6559[71]), 
          .B1(cout), .C1(n78_adj_6388), .D1(integrator3_adj_6560[71]), 
          .CIN(n16261), .S0(integrator3_71__N_1104_adj_6575[70]), .S1(integrator3_71__N_1104_adj_6575[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_35 (.A0(integrator2_adj_6559[68]), .B0(cout), 
          .C0(n87_adj_6391), .D0(integrator3_adj_6560[68]), .A1(integrator2_adj_6559[69]), 
          .B1(cout), .C1(n84_adj_6390), .D1(integrator3_adj_6560[69]), 
          .CIN(n16260), .COUT(n16261), .S0(integrator3_71__N_1104_adj_6575[68]), 
          .S1(integrator3_71__N_1104_adj_6575[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_33 (.A0(integrator2_adj_6559[66]), .B0(cout), 
          .C0(n93_adj_6393), .D0(integrator3_adj_6560[66]), .A1(integrator2_adj_6559[67]), 
          .B1(cout), .C1(n90_adj_6392), .D1(integrator3_adj_6560[67]), 
          .CIN(n16259), .COUT(n16260), .S0(integrator3_71__N_1104_adj_6575[66]), 
          .S1(integrator3_71__N_1104_adj_6575[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_31 (.A0(integrator2_adj_6559[64]), .B0(cout), 
          .C0(n99_adj_6395), .D0(integrator3_adj_6560[64]), .A1(integrator2_adj_6559[65]), 
          .B1(cout), .C1(n96_adj_6394), .D1(integrator3_adj_6560[65]), 
          .CIN(n16258), .COUT(n16259), .S0(integrator3_71__N_1104_adj_6575[64]), 
          .S1(integrator3_71__N_1104_adj_6575[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_29 (.A0(integrator2_adj_6559[62]), .B0(cout), 
          .C0(n105_adj_6397), .D0(integrator3_adj_6560[62]), .A1(integrator2_adj_6559[63]), 
          .B1(cout), .C1(n102_adj_6396), .D1(integrator3_adj_6560[63]), 
          .CIN(n16257), .COUT(n16258), .S0(integrator3_71__N_1104_adj_6575[62]), 
          .S1(integrator3_71__N_1104_adj_6575[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_27 (.A0(integrator2_adj_6559[60]), .B0(cout), 
          .C0(n111_adj_6399), .D0(integrator3_adj_6560[60]), .A1(integrator2_adj_6559[61]), 
          .B1(cout), .C1(n108_adj_6398), .D1(integrator3_adj_6560[61]), 
          .CIN(n16256), .COUT(n16257), .S0(integrator3_71__N_1104_adj_6575[60]), 
          .S1(integrator3_71__N_1104_adj_6575[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_8 (.A0(comb_d9_adj_6570[5]), .B0(comb9_adj_6569[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[6]), .B1(comb9_adj_6569[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17700), .COUT(n17701));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_8.INJECT1_1 = "NO";
    LUT4 phase_increment_1__63__N_21_23__bdd_2_lut_9021 (.A(phase_increment_1__63__N_21[23]), 
         .B(rx_byte[0]), .Z(n19581)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_23__bdd_2_lut_9021.init = 16'heeee;
    CCU2C _add_1_3651_add_4_15 (.A0(comb7_adj_6565[48]), .B0(cout_adj_5840), 
          .C0(n147_adj_5698), .D0(n25_adj_5551), .A1(comb7_adj_6565[49]), 
          .B1(cout_adj_5840), .C1(n144_adj_5697), .D1(n24_adj_5550), .CIN(n17196), 
          .COUT(n17197), .S0(comb8_71__N_2137_adj_6591[48]), .S1(comb8_71__N_2137_adj_6591[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_13 (.A0(comb7_adj_6565[46]), .B0(cout_adj_5840), 
          .C0(n153_adj_5700), .D0(n27_adj_5553), .A1(comb7_adj_6565[47]), 
          .B1(cout_adj_5840), .C1(n150_adj_5699), .D1(n26_adj_5552), .CIN(n17195), 
          .COUT(n17196), .S0(comb8_71__N_2137_adj_6591[46]), .S1(comb8_71__N_2137_adj_6591[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_6 (.A0(comb_d9_adj_6570[3]), .B0(comb9_adj_6569[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[4]), .B1(comb9_adj_6569[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17699), .COUT(n17700));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_11 (.A0(comb7_adj_6565[44]), .B0(cout_adj_5840), 
          .C0(n159_adj_5702), .D0(n29_adj_5555), .A1(comb7_adj_6565[45]), 
          .B1(cout_adj_5840), .C1(n156_adj_5701), .D1(n28_adj_5554), .CIN(n17194), 
          .COUT(n17195), .S0(comb8_71__N_2137_adj_6591[44]), .S1(comb8_71__N_2137_adj_6591[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3597_add_4_13 (.A0(cosine_table_value[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17503), .S0(n28_adj_6338));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[48:67])
    defparam _add_1_3597_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_3597_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_3597_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3597_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_9 (.A0(comb7_adj_6565[42]), .B0(cout_adj_5840), 
          .C0(n165_adj_5704), .D0(n31_adj_5557), .A1(comb7_adj_6565[43]), 
          .B1(cout_adj_5840), .C1(n162_adj_5703), .D1(n30_adj_5556), .CIN(n17193), 
          .COUT(n17194), .S0(comb8_71__N_2137_adj_6591[42]), .S1(comb8_71__N_2137_adj_6591[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_25 (.A0(integrator2_adj_6559[58]), .B0(cout), 
          .C0(n117_adj_6401), .D0(integrator3_adj_6560[58]), .A1(integrator2_adj_6559[59]), 
          .B1(cout), .C1(n114_adj_6400), .D1(integrator3_adj_6560[59]), 
          .CIN(n16255), .COUT(n16256), .S0(integrator3_71__N_1104_adj_6575[58]), 
          .S1(integrator3_71__N_1104_adj_6575[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_23 (.A0(integrator2_adj_6559[56]), .B0(cout), 
          .C0(n123_adj_6403), .D0(integrator3_adj_6560[56]), .A1(integrator2_adj_6559[57]), 
          .B1(cout), .C1(n120_adj_6402), .D1(integrator3_adj_6560[57]), 
          .CIN(n16254), .COUT(n16255), .S0(integrator3_71__N_1104_adj_6575[56]), 
          .S1(integrator3_71__N_1104_adj_6575[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_21 (.A0(integrator2_adj_6559[54]), .B0(cout), 
          .C0(n129_adj_6405), .D0(integrator3_adj_6560[54]), .A1(integrator2_adj_6559[55]), 
          .B1(cout), .C1(n126_adj_6404), .D1(integrator3_adj_6560[55]), 
          .CIN(n16253), .COUT(n16254), .S0(integrator3_71__N_1104_adj_6575[54]), 
          .S1(integrator3_71__N_1104_adj_6575[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_19 (.A0(integrator2_adj_6559[52]), .B0(cout), 
          .C0(n135_adj_6407), .D0(integrator3_adj_6560[52]), .A1(integrator2_adj_6559[53]), 
          .B1(cout), .C1(n132_adj_6406), .D1(integrator3_adj_6560[53]), 
          .CIN(n16252), .COUT(n16253), .S0(integrator3_71__N_1104_adj_6575[52]), 
          .S1(integrator3_71__N_1104_adj_6575[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_17 (.A0(integrator2_adj_6559[50]), .B0(cout), 
          .C0(n141_adj_6409), .D0(integrator3_adj_6560[50]), .A1(integrator2_adj_6559[51]), 
          .B1(cout), .C1(n138_adj_6408), .D1(integrator3_adj_6560[51]), 
          .CIN(n16251), .COUT(n16252), .S0(integrator3_71__N_1104_adj_6575[50]), 
          .S1(integrator3_71__N_1104_adj_6575[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_15 (.A0(integrator2_adj_6559[48]), .B0(cout), 
          .C0(n147_adj_6411), .D0(integrator3_adj_6560[48]), .A1(integrator2_adj_6559[49]), 
          .B1(cout), .C1(n144_adj_6410), .D1(integrator3_adj_6560[49]), 
          .CIN(n16250), .COUT(n16251), .S0(integrator3_71__N_1104_adj_6575[48]), 
          .S1(integrator3_71__N_1104_adj_6575[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_13 (.A0(integrator2_adj_6559[46]), .B0(cout), 
          .C0(n153_adj_6413), .D0(integrator3_adj_6560[46]), .A1(integrator2_adj_6559[47]), 
          .B1(cout), .C1(n150_adj_6412), .D1(integrator3_adj_6560[47]), 
          .CIN(n16249), .COUT(n16250), .S0(integrator3_71__N_1104_adj_6575[46]), 
          .S1(integrator3_71__N_1104_adj_6575[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_11 (.A0(integrator2_adj_6559[44]), .B0(cout), 
          .C0(n159_adj_6415), .D0(integrator3_adj_6560[44]), .A1(integrator2_adj_6559[45]), 
          .B1(cout), .C1(n156_adj_6414), .D1(integrator3_adj_6560[45]), 
          .CIN(n16248), .COUT(n16249), .S0(integrator3_71__N_1104_adj_6575[44]), 
          .S1(integrator3_71__N_1104_adj_6575[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_9 (.A0(integrator2_adj_6559[42]), .B0(cout), 
          .C0(n165_adj_6417), .D0(integrator3_adj_6560[42]), .A1(integrator2_adj_6559[43]), 
          .B1(cout), .C1(n162_adj_6416), .D1(integrator3_adj_6560[43]), 
          .CIN(n16247), .COUT(n16248), .S0(integrator3_71__N_1104_adj_6575[42]), 
          .S1(integrator3_71__N_1104_adj_6575[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_7 (.A0(integrator2_adj_6559[40]), .B0(cout), 
          .C0(n171_adj_6419), .D0(integrator3_adj_6560[40]), .A1(integrator2_adj_6559[41]), 
          .B1(cout), .C1(n168_adj_6418), .D1(integrator3_adj_6560[41]), 
          .CIN(n16246), .COUT(n16247), .S0(integrator3_71__N_1104_adj_6575[40]), 
          .S1(integrator3_71__N_1104_adj_6575[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_5 (.A0(integrator2_adj_6559[38]), .B0(cout), 
          .C0(n177_adj_6421), .D0(integrator3_adj_6560[38]), .A1(integrator2_adj_6559[39]), 
          .B1(cout), .C1(n174_adj_6420), .D1(integrator3_adj_6560[39]), 
          .CIN(n16245), .COUT(n16246), .S0(integrator3_71__N_1104_adj_6575[38]), 
          .S1(integrator3_71__N_1104_adj_6575[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_3 (.A0(integrator2_adj_6559[36]), .B0(cout), 
          .C0(n183_adj_6423), .D0(integrator3_adj_6560[36]), .A1(integrator2_adj_6559[37]), 
          .B1(cout), .C1(n180_adj_6422), .D1(integrator3_adj_6560[37]), 
          .CIN(n16244), .COUT(n16245), .S0(integrator3_71__N_1104_adj_6575[36]), 
          .S1(integrator3_71__N_1104_adj_6575[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3666_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3666_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3666_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16244));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3666_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3666_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3666_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3666_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_37 (.A0(integrator1_adj_6558[70]), .B0(cout_adj_5269), 
          .C0(n81_adj_6291), .D0(integrator2_adj_6559[70]), .A1(integrator1_adj_6558[71]), 
          .B1(cout_adj_5269), .C1(n78_adj_6290), .D1(integrator2_adj_6559[71]), 
          .CIN(n16239), .S0(integrator2_71__N_1032_adj_6574[70]), .S1(integrator2_71__N_1032_adj_6574[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_35 (.A0(integrator1_adj_6558[68]), .B0(cout_adj_5269), 
          .C0(n87_adj_6293), .D0(integrator2_adj_6559[68]), .A1(integrator1_adj_6558[69]), 
          .B1(cout_adj_5269), .C1(n84_adj_6292), .D1(integrator2_adj_6559[69]), 
          .CIN(n16238), .COUT(n16239), .S0(integrator2_71__N_1032_adj_6574[68]), 
          .S1(integrator2_71__N_1032_adj_6574[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_33 (.A0(integrator1_adj_6558[66]), .B0(cout_adj_5269), 
          .C0(n93_adj_6295), .D0(integrator2_adj_6559[66]), .A1(integrator1_adj_6558[67]), 
          .B1(cout_adj_5269), .C1(n90_adj_6294), .D1(integrator2_adj_6559[67]), 
          .CIN(n16237), .COUT(n16238), .S0(integrator2_71__N_1032_adj_6574[66]), 
          .S1(integrator2_71__N_1032_adj_6574[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_31 (.A0(integrator1_adj_6558[64]), .B0(cout_adj_5269), 
          .C0(n99_adj_6297), .D0(integrator2_adj_6559[64]), .A1(integrator1_adj_6558[65]), 
          .B1(cout_adj_5269), .C1(n96_adj_6296), .D1(integrator2_adj_6559[65]), 
          .CIN(n16236), .COUT(n16237), .S0(integrator2_71__N_1032_adj_6574[64]), 
          .S1(integrator2_71__N_1032_adj_6574[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_29 (.A0(integrator1_adj_6558[62]), .B0(cout_adj_5269), 
          .C0(n105_adj_6299), .D0(integrator2_adj_6559[62]), .A1(integrator1_adj_6558[63]), 
          .B1(cout_adj_5269), .C1(n102_adj_6298), .D1(integrator2_adj_6559[63]), 
          .CIN(n16235), .COUT(n16236), .S0(integrator2_71__N_1032_adj_6574[62]), 
          .S1(integrator2_71__N_1032_adj_6574[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_27 (.A0(integrator1_adj_6558[60]), .B0(cout_adj_5269), 
          .C0(n111_adj_6301), .D0(integrator2_adj_6559[60]), .A1(integrator1_adj_6558[61]), 
          .B1(cout_adj_5269), .C1(n108_adj_6300), .D1(integrator2_adj_6559[61]), 
          .CIN(n16234), .COUT(n16235), .S0(integrator2_71__N_1032_adj_6574[60]), 
          .S1(integrator2_71__N_1032_adj_6574[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_25 (.A0(integrator1_adj_6558[58]), .B0(cout_adj_5269), 
          .C0(n117_adj_6303), .D0(integrator2_adj_6559[58]), .A1(integrator1_adj_6558[59]), 
          .B1(cout_adj_5269), .C1(n114_adj_6302), .D1(integrator2_adj_6559[59]), 
          .CIN(n16233), .COUT(n16234), .S0(integrator2_71__N_1032_adj_6574[58]), 
          .S1(integrator2_71__N_1032_adj_6574[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_23 (.A0(integrator1_adj_6558[56]), .B0(cout_adj_5269), 
          .C0(n123_adj_6305), .D0(integrator2_adj_6559[56]), .A1(integrator1_adj_6558[57]), 
          .B1(cout_adj_5269), .C1(n120_adj_6304), .D1(integrator2_adj_6559[57]), 
          .CIN(n16232), .COUT(n16233), .S0(integrator2_71__N_1032_adj_6574[56]), 
          .S1(integrator2_71__N_1032_adj_6574[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_21 (.A0(integrator1_adj_6558[54]), .B0(cout_adj_5269), 
          .C0(n129_adj_6307), .D0(integrator2_adj_6559[54]), .A1(integrator1_adj_6558[55]), 
          .B1(cout_adj_5269), .C1(n126_adj_6306), .D1(integrator2_adj_6559[55]), 
          .CIN(n16231), .COUT(n16232), .S0(integrator2_71__N_1032_adj_6574[54]), 
          .S1(integrator2_71__N_1032_adj_6574[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_19 (.A0(integrator1_adj_6558[52]), .B0(cout_adj_5269), 
          .C0(n135_adj_6309), .D0(integrator2_adj_6559[52]), .A1(integrator1_adj_6558[53]), 
          .B1(cout_adj_5269), .C1(n132_adj_6308), .D1(integrator2_adj_6559[53]), 
          .CIN(n16230), .COUT(n16231), .S0(integrator2_71__N_1032_adj_6574[52]), 
          .S1(integrator2_71__N_1032_adj_6574[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_17 (.A0(integrator1_adj_6558[50]), .B0(cout_adj_5269), 
          .C0(n141_adj_6311), .D0(integrator2_adj_6559[50]), .A1(integrator1_adj_6558[51]), 
          .B1(cout_adj_5269), .C1(n138_adj_6310), .D1(integrator2_adj_6559[51]), 
          .CIN(n16229), .COUT(n16230), .S0(integrator2_71__N_1032_adj_6574[50]), 
          .S1(integrator2_71__N_1032_adj_6574[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_15 (.A0(integrator1_adj_6558[48]), .B0(cout_adj_5269), 
          .C0(n147_adj_6313), .D0(integrator2_adj_6559[48]), .A1(integrator1_adj_6558[49]), 
          .B1(cout_adj_5269), .C1(n144_adj_6312), .D1(integrator2_adj_6559[49]), 
          .CIN(n16228), .COUT(n16229), .S0(integrator2_71__N_1032_adj_6574[48]), 
          .S1(integrator2_71__N_1032_adj_6574[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_13 (.A0(integrator1_adj_6558[46]), .B0(cout_adj_5269), 
          .C0(n153_adj_6315), .D0(integrator2_adj_6559[46]), .A1(integrator1_adj_6558[47]), 
          .B1(cout_adj_5269), .C1(n150_adj_6314), .D1(integrator2_adj_6559[47]), 
          .CIN(n16227), .COUT(n16228), .S0(integrator2_71__N_1032_adj_6574[46]), 
          .S1(integrator2_71__N_1032_adj_6574[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_11 (.A0(integrator1_adj_6558[44]), .B0(cout_adj_5269), 
          .C0(n159_adj_6317), .D0(integrator2_adj_6559[44]), .A1(integrator1_adj_6558[45]), 
          .B1(cout_adj_5269), .C1(n156_adj_6316), .D1(integrator2_adj_6559[45]), 
          .CIN(n16226), .COUT(n16227), .S0(integrator2_71__N_1032_adj_6574[44]), 
          .S1(integrator2_71__N_1032_adj_6574[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_9 (.A0(integrator1_adj_6558[42]), .B0(cout_adj_5269), 
          .C0(n165_adj_6319), .D0(integrator2_adj_6559[42]), .A1(integrator1_adj_6558[43]), 
          .B1(cout_adj_5269), .C1(n162_adj_6318), .D1(integrator2_adj_6559[43]), 
          .CIN(n16225), .COUT(n16226), .S0(integrator2_71__N_1032_adj_6574[42]), 
          .S1(integrator2_71__N_1032_adj_6574[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_7 (.A0(integrator1_adj_6558[40]), .B0(cout_adj_5269), 
          .C0(n171_adj_6321), .D0(integrator2_adj_6559[40]), .A1(integrator1_adj_6558[41]), 
          .B1(cout_adj_5269), .C1(n168_adj_6320), .D1(integrator2_adj_6559[41]), 
          .CIN(n16224), .COUT(n16225), .S0(integrator2_71__N_1032_adj_6574[40]), 
          .S1(integrator2_71__N_1032_adj_6574[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_5 (.A0(integrator1_adj_6558[38]), .B0(cout_adj_5269), 
          .C0(n177_adj_6323), .D0(integrator2_adj_6559[38]), .A1(integrator1_adj_6558[39]), 
          .B1(cout_adj_5269), .C1(n174_adj_6322), .D1(integrator2_adj_6559[39]), 
          .CIN(n16223), .COUT(n16224), .S0(integrator2_71__N_1032_adj_6574[38]), 
          .S1(integrator2_71__N_1032_adj_6574[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_3 (.A0(integrator1_adj_6558[36]), .B0(cout_adj_5269), 
          .C0(n183_adj_6325), .D0(integrator2_adj_6559[36]), .A1(integrator1_adj_6558[37]), 
          .B1(cout_adj_5269), .C1(n180_adj_6324), .D1(integrator2_adj_6559[37]), 
          .CIN(n16222), .COUT(n16223), .S0(integrator2_71__N_1032_adj_6574[36]), 
          .S1(integrator2_71__N_1032_adj_6574[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3669_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3669_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3669_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5269), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16222));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3669_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3669_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3669_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3669_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3597_add_4_11 (.A0(cosine_table_value[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cosine_table_value[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17502), .COUT(n17503), .S0(n34_adj_6340), 
          .S1(n31_adj_6339));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[48:67])
    defparam _add_1_3597_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_3597_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_3597_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3597_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3597_add_4_9 (.A0(cosine_table_value[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cosine_table_value[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17501), .COUT(n17502), .S0(n40_adj_6342), 
          .S1(n37_adj_6341));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[48:67])
    defparam _add_1_3597_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_3597_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_3597_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3597_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3597_add_4_7 (.A0(cosine_table_value[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cosine_table_value[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17500), .COUT(n17501), .S0(n46_adj_6344), 
          .S1(n43_adj_6343));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[48:67])
    defparam _add_1_3597_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_3597_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_3597_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3597_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3597_add_4_5 (.A0(cosine_table_value[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cosine_table_value[4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17499), .COUT(n17500), .S0(n52_adj_6346), 
          .S1(n49_adj_6345));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[48:67])
    defparam _add_1_3597_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_3597_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_3597_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3597_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3597_add_4_3 (.A0(cosine_table_value[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cosine_table_value[2]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17498), .COUT(n17499), .S0(n58_adj_6348), 
          .S1(n55_adj_6347));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[48:67])
    defparam _add_1_3597_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_3597_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_3597_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3597_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3597_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cosine_table_value[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17498), .S1(n61_adj_6349));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[48:67])
    defparam _add_1_3597_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3597_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_3597_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3597_add_4_1.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_26 (.A0(q_squared[23]), .B0(i_squared[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17497), .S0(n54));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_26.INIT0 = 16'h666a;
    defparam square_sum_add_4_26.INIT1 = 16'h0000;
    defparam square_sum_add_4_26.INJECT1_0 = "NO";
    defparam square_sum_add_4_26.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_24 (.A0(q_squared[22]), .B0(i_squared[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(q_squared[23]), .B1(i_squared[23]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17496), .COUT(n17497), .S0(n60), .S1(n57));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_24.INIT0 = 16'h666a;
    defparam square_sum_add_4_24.INIT1 = 16'h666a;
    defparam square_sum_add_4_24.INJECT1_0 = "NO";
    defparam square_sum_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_4 (.A0(comb_d9_adj_6570[1]), .B0(comb9_adj_6569[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6570[2]), .B1(comb9_adj_6569[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17698), .COUT(n17699));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3801_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3801_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9_adj_6570[0]), .B1(comb9_adj_6569[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n17698));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3801_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3801_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3801_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3801_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_61 (.A0(\phase_increment[0] [63]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17697), .S0(phase_increment_1__63__N_16[63]));
    defparam _add_1_3804_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_61.INIT1 = 16'h0000;
    defparam _add_1_3804_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_61.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_14 (.A0(integrator5_adj_6562[47]), .B0(integrator4_adj_6561[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[48]), .B1(integrator4_adj_6561[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17408), .COUT(n17409), .S0(n150_adj_6498), 
          .S1(n147_adj_6497));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_59 (.A0(\phase_increment[0] [61]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [62]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17696), .COUT(n17697), .S0(phase_increment_1__63__N_16[61]), 
          .S1(phase_increment_1__63__N_16[62]));
    defparam _add_1_3804_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_57 (.A0(\phase_increment[0] [59]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [60]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17695), .COUT(n17696), .S0(phase_increment_1__63__N_16[59]), 
          .S1(phase_increment_1__63__N_16[60]));
    defparam _add_1_3804_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_55 (.A0(\phase_increment[0] [57]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [58]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17694), .COUT(n17695), .S0(phase_increment_1__63__N_16[57]), 
          .S1(phase_increment_1__63__N_16[58]));
    defparam _add_1_3804_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_53 (.A0(\phase_increment[0] [55]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [56]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17693), .COUT(n17694), .S0(phase_increment_1__63__N_16[55]), 
          .S1(phase_increment_1__63__N_16[56]));
    defparam _add_1_3804_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_51 (.A0(\phase_increment[0] [53]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [54]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17692), .COUT(n17693), .S0(phase_increment_1__63__N_16[53]), 
          .S1(phase_increment_1__63__N_16[54]));
    defparam _add_1_3804_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_49 (.A0(\phase_increment[0] [51]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [52]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17691), .COUT(n17692), .S0(phase_increment_1__63__N_16[51]), 
          .S1(phase_increment_1__63__N_16[52]));
    defparam _add_1_3804_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_47 (.A0(\phase_increment[0] [49]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [50]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17690), .COUT(n17691), .S0(phase_increment_1__63__N_16[49]), 
          .S1(phase_increment_1__63__N_16[50]));
    defparam _add_1_3804_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_3804_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_45 (.A0(\phase_increment[0] [47]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [48]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17689), .COUT(n17690), .S0(phase_increment_1__63__N_16[47]), 
          .S1(phase_increment_1__63__N_16[48]));
    defparam _add_1_3804_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_45.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_43 (.A0(\phase_increment[0] [45]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [46]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17688), .COUT(n17689), .S0(phase_increment_1__63__N_16[45]), 
          .S1(phase_increment_1__63__N_16[46]));
    defparam _add_1_3804_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_43.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_43.INJECT1_1 = "NO";
    FD1S3AX square_sum_e3__i3 (.D(n120_adj_5602), .CK(cic_sine_clk), .Q(square_sum[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i3.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i4 (.D(n117_adj_5603), .CK(cic_sine_clk), .Q(square_sum[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i4.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i5 (.D(n114_adj_5604), .CK(cic_sine_clk), .Q(square_sum[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i5.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i6 (.D(n111_adj_5605), .CK(cic_sine_clk), .Q(square_sum[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i6.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i7 (.D(n108_adj_5606), .CK(cic_sine_clk), .Q(square_sum[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i7.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i8 (.D(n105_adj_5607), .CK(cic_sine_clk), .Q(square_sum[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i8.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i9 (.D(n102_adj_5608), .CK(cic_sine_clk), .Q(square_sum[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i9.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i10 (.D(n99_adj_5609), .CK(cic_sine_clk), .Q(square_sum[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i10.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i11 (.D(n96_adj_5610), .CK(cic_sine_clk), .Q(square_sum[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i11.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i12 (.D(n93_adj_5611), .CK(cic_sine_clk), .Q(square_sum[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i12.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i13 (.D(n90), .CK(cic_sine_clk), .Q(square_sum[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i13.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i14 (.D(n87), .CK(cic_sine_clk), .Q(square_sum[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i14.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i15 (.D(n84), .CK(cic_sine_clk), .Q(square_sum[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i15.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i16 (.D(n81), .CK(cic_sine_clk), .Q(square_sum[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i16.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i17 (.D(n78), .CK(cic_sine_clk), .Q(square_sum[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i17.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i18 (.D(n75), .CK(cic_sine_clk), .Q(square_sum[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i18.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i19 (.D(n72), .CK(cic_sine_clk), .Q(square_sum[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i19.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i20 (.D(n69), .CK(cic_sine_clk), .Q(square_sum[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i20.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i21 (.D(n66), .CK(cic_sine_clk), .Q(square_sum[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i21.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i22 (.D(n63), .CK(cic_sine_clk), .Q(square_sum[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i22.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i23 (.D(n60), .CK(cic_sine_clk), .Q(square_sum[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i23.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i24 (.D(n57), .CK(cic_sine_clk), .Q(square_sum[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i24.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i25 (.D(n54), .CK(cic_sine_clk), .Q(square_sum[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_e3__i25.GSR = "ENABLED";
    CCU2C _add_1_3804_add_4_41 (.A0(\phase_increment[0] [43]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [44]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17687), .COUT(n17688), .S0(phase_increment_1__63__N_16[43]), 
          .S1(phase_increment_1__63__N_16[44]));
    defparam _add_1_3804_add_4_41.INIT0 = 16'haaa0;
    defparam _add_1_3804_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_39 (.A0(\phase_increment[0] [41]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [42]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17686), .COUT(n17687), .S0(phase_increment_1__63__N_16[41]), 
          .S1(phase_increment_1__63__N_16[42]));
    defparam _add_1_3804_add_4_39.INIT0 = 16'haaa0;
    defparam _add_1_3804_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_37 (.A0(\phase_increment[0] [39]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [40]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17685), .COUT(n17686), .S0(phase_increment_1__63__N_16[39]), 
          .S1(phase_increment_1__63__N_16[40]));
    defparam _add_1_3804_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_37.INJECT1_1 = "NO";
    FD1P3AX cic_gain__i2 (.D(cic_gain_7__N_544[1]), .SP(rx_data_valid), 
            .CK(clk_80mhz), .Q(cic_gain[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam cic_gain__i2.GSR = "ENABLED";
    CCU2C square_sum_add_4_22 (.A0(q_squared[20]), .B0(i_squared[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(q_squared[21]), .B1(i_squared[21]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17495), .COUT(n17496), .S0(n66), .S1(n63));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_22.INIT0 = 16'h666a;
    defparam square_sum_add_4_22.INIT1 = 16'h666a;
    defparam square_sum_add_4_22.INJECT1_0 = "NO";
    defparam square_sum_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_35 (.A0(\phase_increment[0] [37]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [38]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17684), .COUT(n17685), .S0(phase_increment_1__63__N_16[37]), 
          .S1(phase_increment_1__63__N_16[38]));
    defparam _add_1_3804_add_4_35.INIT0 = 16'haaa0;
    defparam _add_1_3804_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_33 (.A0(\phase_increment[0] [35]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [36]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17683), .COUT(n17684), .S0(phase_increment_1__63__N_16[35]), 
          .S1(phase_increment_1__63__N_16[36]));
    defparam _add_1_3804_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_31 (.A0(\phase_increment[0] [33]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [34]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17682), .COUT(n17683), .S0(phase_increment_1__63__N_16[33]), 
          .S1(phase_increment_1__63__N_16[34]));
    defparam _add_1_3804_add_4_31.INIT0 = 16'haaa0;
    defparam _add_1_3804_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_29 (.A0(\phase_increment[0] [31]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [32]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17681), .COUT(n17682), .S0(phase_increment_1__63__N_16[31]), 
          .S1(phase_increment_1__63__N_16[32]));
    defparam _add_1_3804_add_4_29.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_29.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_12 (.A0(integrator5_adj_6562[45]), .B0(integrator4_adj_6561[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[46]), .B1(integrator4_adj_6561[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17407), .COUT(n17408), .S0(n156_adj_6500), 
          .S1(n153_adj_6499));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_27 (.A0(\phase_increment[0] [29]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [30]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17680), .COUT(n17681), .S0(phase_increment_1__63__N_16[29]), 
          .S1(phase_increment_1__63__N_16[30]));
    defparam _add_1_3804_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_25 (.A0(\phase_increment[0] [27]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [28]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17679), .COUT(n17680), .S0(phase_increment_1__63__N_16[27]), 
          .S1(phase_increment_1__63__N_16[28]));
    defparam _add_1_3804_add_4_25.INIT0 = 16'haaa0;
    defparam _add_1_3804_add_4_25.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_23 (.A0(\phase_increment[0] [25]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [26]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17678), .COUT(n17679), .S0(phase_increment_1__63__N_16[25]), 
          .S1(phase_increment_1__63__N_16[26]));
    defparam _add_1_3804_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_21 (.A0(\phase_increment[0] [23]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [24]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17677), .COUT(n17678), .S0(phase_increment_1__63__N_16[23]), 
          .S1(phase_increment_1__63__N_16[24]));
    defparam _add_1_3804_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_21.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_20 (.A0(q_squared[18]), .B0(i_squared[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(q_squared[19]), .B1(i_squared[19]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17494), .COUT(n17495), .S0(n72), .S1(n69));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_20.INIT0 = 16'h666a;
    defparam square_sum_add_4_20.INIT1 = 16'h666a;
    defparam square_sum_add_4_20.INJECT1_0 = "NO";
    defparam square_sum_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_19 (.A0(\phase_increment[0] [21]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [22]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17676), .COUT(n17677), .S0(phase_increment_1__63__N_16[21]), 
          .S1(phase_increment_1__63__N_16[22]));
    defparam _add_1_3804_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_3804_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_17 (.A0(\phase_increment[0] [19]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [20]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17675), .COUT(n17676), .S0(phase_increment_1__63__N_16[19]), 
          .S1(phase_increment_1__63__N_16[20]));
    defparam _add_1_3804_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_3804_add_4_17.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_15 (.A0(\phase_increment[0] [17]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [18]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17674), .COUT(n17675), .S0(phase_increment_1__63__N_16[17]), 
          .S1(phase_increment_1__63__N_16[18]));
    defparam _add_1_3804_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_15.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_30 (.A0(integrator4_adj_6561[63]), .B0(integrator3_adj_6560[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[64]), .B1(integrator3_adj_6560[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17442), .COUT(n17443), .S0(n102_adj_6432), 
          .S1(n99_adj_6431));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_13 (.A0(\phase_increment[0] [15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [16]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17673), .COUT(n17674), .S0(phase_increment_1__63__N_16[15]), 
          .S1(phase_increment_1__63__N_16[16]));
    defparam _add_1_3804_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3804_add_4_13.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_11 (.A0(\phase_increment[0] [13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17672), .COUT(n17673), .S0(phase_increment_1__63__N_16[13]), 
          .S1(phase_increment_1__63__N_16[14]));
    defparam _add_1_3804_add_4_11.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_9 (.A0(\phase_increment[0] [11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17671), .COUT(n17672), .S0(phase_increment_1__63__N_16[11]), 
          .S1(phase_increment_1__63__N_16[12]));
    defparam _add_1_3804_add_4_9.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_7 (.A0(\phase_increment[0] [9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17670), .COUT(n17671), .S0(phase_increment_1__63__N_16[9]), 
          .S1(phase_increment_1__63__N_16[10]));
    defparam _add_1_3804_add_4_7.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_7.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_18 (.A0(q_squared[16]), .B0(i_squared[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(q_squared[17]), .B1(i_squared[17]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17493), .COUT(n17494), .S0(n78), .S1(n75));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_18.INIT0 = 16'h666a;
    defparam square_sum_add_4_18.INIT1 = 16'h666a;
    defparam square_sum_add_4_18.INJECT1_0 = "NO";
    defparam square_sum_add_4_18.INJECT1_1 = "NO";
    LUT4 mux_2557_i1_3_lut (.A(phase_increment_1__63__N_16[4]), .B(phase_increment_1__63__N_18[4]), 
         .C(rx_byte[0]), .Z(n4186)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2557_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3804_add_4_5 (.A0(\phase_increment[0] [7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17669), .COUT(n17670), .S0(phase_increment_1__63__N_16[7]), 
          .S1(phase_increment_1__63__N_16[8]));
    defparam _add_1_3804_add_4_5.INIT0 = 16'h555f;
    defparam _add_1_3804_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_3 (.A0(\phase_increment[0] [5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17668), .COUT(n17669), .S0(phase_increment_1__63__N_16[5]), 
          .S1(phase_increment_1__63__N_16[6]));
    defparam _add_1_3804_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_3804_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_3804_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3804_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\phase_increment[0] [4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17668), .S1(phase_increment_1__63__N_16[4]));
    defparam _add_1_3804_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3804_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3804_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3804_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_10 (.A0(integrator5_adj_6562[43]), .B0(integrator4_adj_6561[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[44]), .B1(integrator4_adj_6561[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17406), .COUT(n17407), .S0(n162_adj_6502), 
          .S1(n159_adj_6501));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_7 (.A0(comb7_adj_6565[40]), .B0(cout_adj_5840), 
          .C0(n171_adj_5706), .D0(n33_adj_5559), .A1(comb7_adj_6565[41]), 
          .B1(cout_adj_5840), .C1(n168_adj_5705), .D1(n32_adj_5558), .CIN(n17192), 
          .COUT(n17193), .S0(comb8_71__N_2137_adj_6591[40]), .S1(comb8_71__N_2137_adj_6591[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_65 (.A0(\phase_increment[0] [63]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17662), .S0(phase_increment_1__63__N_18[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_65.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_65.INIT1 = 16'h0000;
    defparam _add_1_3807_add_4_65.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_65.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_63 (.A0(\phase_increment[0] [61]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [62]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17661), .COUT(n17662), .S0(phase_increment_1__63__N_18[61]), 
          .S1(phase_increment_1__63__N_18[62]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_63.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_63.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_63.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_63.INJECT1_1 = "NO";
    CCU2C _add_1_3651_add_4_5 (.A0(comb7_adj_6565[38]), .B0(cout_adj_5840), 
          .C0(n177_adj_5708), .D0(n35_adj_5561), .A1(comb7_adj_6565[39]), 
          .B1(cout_adj_5840), .C1(n174_adj_5707), .D1(n34_adj_5560), .CIN(n17191), 
          .COUT(n17192), .S0(comb8_71__N_2137_adj_6591[38]), .S1(comb8_71__N_2137_adj_6591[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_5.INJECT1_1 = "NO";
    LUT4 i4981_4_lut (.A(phase_increment_1__63__N_16[21]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[21]), .D(rx_byte[0]), .Z(n3412)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4981_4_lut.init = 16'hc088;
    CCU2C _add_1_3651_add_4_3 (.A0(comb7_adj_6565[36]), .B0(cout_adj_5840), 
          .C0(n183_adj_5710), .D0(n37_adj_5563), .A1(comb7_adj_6565[37]), 
          .B1(cout_adj_5840), .C1(n180_adj_5709), .D1(n36_adj_5562), .CIN(n17190), 
          .COUT(n17191), .S0(comb8_71__N_2137_adj_6591[36]), .S1(comb8_71__N_2137_adj_6591[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3651_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3651_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_61 (.A0(\phase_increment[0] [59]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [60]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17660), .COUT(n17661), .S0(phase_increment_1__63__N_18[59]), 
          .S1(phase_increment_1__63__N_18[60]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_61.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_61.INJECT1_1 = "NO";
    PFUMX mux_1358_i1 (.BLUT(n2566), .ALUT(n2572), .C0(n19300), .Z(n2575));
    LUT4 phase_increment_1__63__N_21_39__bdd_2_lut_8895 (.A(phase_increment_1__63__N_21[39]), 
         .B(rx_byte[0]), .Z(n19648)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_39__bdd_2_lut_8895.init = 16'heeee;
    PLL pll_inst (.clk_25mhz_c(clk_25mhz_c), .clk_80mhz(clk_80mhz), .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(96[8] 99[5])
    CCU2C _add_1_3651_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5840), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17190));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3651_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3651_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3651_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3651_add_4_1.INJECT1_1 = "NO";
    PFUMX mux_1321_i1 (.BLUT(n2509), .ALUT(n2519), .C0(led_0_6), .Z(n2525));
    CCU2C _add_1_3576_add_4_15 (.A0(amdemod_out_d_11__N_2567), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2564), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17185), .S1(amdemod_out_d_11__N_2380[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3576_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3576_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3576_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3576_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3576_add_4_13 (.A0(amdemod_out_d_11__N_2573), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2570), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17184), .COUT(n17185), .S0(amdemod_out_d_11__N_2380[11]), 
          .S1(amdemod_out_d_11__N_2380[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3576_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3576_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3576_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3576_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3576_add_4_11 (.A0(amdemod_out_d_11__N_2579), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2576), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17183), .COUT(n17184), .S0(amdemod_out_d_11__N_2380[9]), 
          .S1(amdemod_out_d_11__N_2380[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3576_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3576_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3576_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3576_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3576_add_4_9 (.A0(amdemod_out_d_11__N_2585), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2582), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17182), .COUT(n17183), .S0(amdemod_out_d_11__N_2380[7]), 
          .S1(amdemod_out_d_11__N_2380[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3576_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_3576_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_3576_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3576_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3576_add_4_7 (.A0(square_sum[25]), .B0(n19824), .C0(amdemod_out_d_11__N_2591), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(amdemod_out_d_11__N_2588), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17181), .COUT(n17182), .S0(amdemod_out_d_11__N_2380[5]), 
          .S1(amdemod_out_d_11__N_2380[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3576_add_4_7.INIT0 = 16'h1e1e;
    defparam _add_1_3576_add_4_7.INIT1 = 16'h666a;
    defparam _add_1_3576_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3576_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3576_add_4_5 (.A0(n19816), .B0(amdemod_out_d_11__N_2597), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2363), .B1(amdemod_out_d_11__N_2594), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17180), .COUT(n17181), .S0(amdemod_out_d_11__N_2380[3]), 
          .S1(amdemod_out_d_11__N_2380[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3576_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3576_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_3576_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3576_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3576_add_4_3 (.A0(n19815), .B0(square_sum[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19815), .B1(amdemod_out_d_11__N_2600), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17179), .COUT(n17180), .S0(amdemod_out_d_11__N_2380[1]), 
          .S1(amdemod_out_d_11__N_2380[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3576_add_4_3.INIT0 = 16'h666a;
    defparam _add_1_3576_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3576_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3576_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3576_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17179), .S1(amdemod_out_d_11__N_2380[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3576_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3576_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3576_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3576_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3579_add_4_15 (.A0(amdemod_out_d_11__N_2645), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2642), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17177), .S1(amdemod_out_d_11__N_2390[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3579_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3579_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3579_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3579_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3579_add_4_13 (.A0(amdemod_out_d_11__N_2651), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2648), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17176), .COUT(n17177), .S0(amdemod_out_d_11__N_2390[11]), 
          .S1(amdemod_out_d_11__N_2390[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3579_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3579_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3579_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3579_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3579_add_4_11 (.A0(amdemod_out_d_11__N_2657), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2654), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17175), .COUT(n17176), .S0(amdemod_out_d_11__N_2390[9]), 
          .S1(amdemod_out_d_11__N_2390[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3579_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3579_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3579_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3579_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3579_add_4_9 (.A0(square_sum[25]), .B0(n19824), .C0(amdemod_out_d_11__N_2663), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(amdemod_out_d_11__N_2660), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17174), .COUT(n17175), .S0(amdemod_out_d_11__N_2390[7]), 
          .S1(amdemod_out_d_11__N_2390[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3579_add_4_9.INIT0 = 16'h1e1e;
    defparam _add_1_3579_add_4_9.INIT1 = 16'h666a;
    defparam _add_1_3579_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3579_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3579_add_4_7 (.A0(n19816), .B0(amdemod_out_d_11__N_2669), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2363), .B1(amdemod_out_d_11__N_2666), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17173), .COUT(n17174), .S0(amdemod_out_d_11__N_2390[5]), 
          .S1(amdemod_out_d_11__N_2390[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3579_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_3579_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_3579_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3579_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3579_add_4_5 (.A0(n19814), .B0(amdemod_out_d_11__N_2675), 
          .C0(GND_net), .D0(VCC_net), .A1(n19815), .B1(amdemod_out_d_11__N_2672), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17172), .COUT(n17173), .S0(amdemod_out_d_11__N_2390[3]), 
          .S1(amdemod_out_d_11__N_2390[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3579_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3579_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_3579_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3579_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3579_add_4_3 (.A0(n19813), .B0(square_sum[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19813), .B1(amdemod_out_d_11__N_2678), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17171), .COUT(n17172), .S0(amdemod_out_d_11__N_2390[1]), 
          .S1(amdemod_out_d_11__N_2390[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3579_add_4_3.INIT0 = 16'h666a;
    defparam _add_1_3579_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3579_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3579_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3579_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17171), .S1(amdemod_out_d_11__N_2390[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3579_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3579_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3579_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3579_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3582_add_4_15 (.A0(amdemod_out_d_11__N_2723), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2720), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17169), .S1(amdemod_out_d_11__N_2400[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3582_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3582_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3582_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3582_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3582_add_4_13 (.A0(amdemod_out_d_11__N_2729), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2726), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17168), .COUT(n17169), .S0(amdemod_out_d_11__N_2400[11]), 
          .S1(amdemod_out_d_11__N_2400[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3582_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3582_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3582_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3582_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3582_add_4_11 (.A0(square_sum[25]), .B0(n19824), .C0(amdemod_out_d_11__N_2735), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(amdemod_out_d_11__N_2732), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17167), .COUT(n17168), .S0(amdemod_out_d_11__N_2400[9]), 
          .S1(amdemod_out_d_11__N_2400[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3582_add_4_11.INIT0 = 16'h1e1e;
    defparam _add_1_3582_add_4_11.INIT1 = 16'h666a;
    defparam _add_1_3582_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3582_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3582_add_4_9 (.A0(n19816), .B0(amdemod_out_d_11__N_2741), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2363), .B1(amdemod_out_d_11__N_2738), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17166), .COUT(n17167), .S0(amdemod_out_d_11__N_2400[7]), 
          .S1(amdemod_out_d_11__N_2400[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3582_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_3582_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_3582_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3582_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3582_add_4_7 (.A0(n19814), .B0(amdemod_out_d_11__N_2747), 
          .C0(GND_net), .D0(VCC_net), .A1(n19815), .B1(amdemod_out_d_11__N_2744), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17165), .COUT(n17166), .S0(amdemod_out_d_11__N_2400[5]), 
          .S1(amdemod_out_d_11__N_2400[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3582_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_3582_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_3582_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3582_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3582_add_4_5 (.A0(n19812), .B0(amdemod_out_d_11__N_2753), 
          .C0(GND_net), .D0(VCC_net), .A1(n19813), .B1(amdemod_out_d_11__N_2750), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17164), .COUT(n17165), .S0(amdemod_out_d_11__N_2400[3]), 
          .S1(amdemod_out_d_11__N_2400[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3582_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3582_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_3582_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3582_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3582_add_4_3 (.A0(n19811), .B0(square_sum[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19811), .B1(amdemod_out_d_11__N_2756), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17163), .COUT(n17164), .S0(amdemod_out_d_11__N_2400[1]), 
          .S1(amdemod_out_d_11__N_2400[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3582_add_4_3.INIT0 = 16'h666a;
    defparam _add_1_3582_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3582_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3582_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3582_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17163), .S1(amdemod_out_d_11__N_2400[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3582_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3582_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3582_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3582_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3585_add_4_15 (.A0(amdemod_out_d_11__N_2801), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2798), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17161), .S1(amdemod_out_d_11__N_2410[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3585_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3585_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3585_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3585_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3585_add_4_13 (.A0(square_sum[25]), .B0(n19824), .C0(amdemod_out_d_11__N_2807), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(amdemod_out_d_11__N_2804), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17160), .COUT(n17161), .S0(amdemod_out_d_11__N_2410[11]), 
          .S1(amdemod_out_d_11__N_2410[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3585_add_4_13.INIT0 = 16'h1e1e;
    defparam _add_1_3585_add_4_13.INIT1 = 16'h666a;
    defparam _add_1_3585_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3585_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3585_add_4_11 (.A0(n19816), .B0(amdemod_out_d_11__N_2813), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2363), .B1(amdemod_out_d_11__N_2810), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17159), .COUT(n17160), .S0(amdemod_out_d_11__N_2410[9]), 
          .S1(amdemod_out_d_11__N_2410[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3585_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_3585_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_3585_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3585_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3585_add_4_9 (.A0(n19814), .B0(amdemod_out_d_11__N_2819), 
          .C0(GND_net), .D0(VCC_net), .A1(n19815), .B1(amdemod_out_d_11__N_2816), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17158), .COUT(n17159), .S0(amdemod_out_d_11__N_2410[7]), 
          .S1(amdemod_out_d_11__N_2410[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3585_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_3585_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_3585_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3585_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3585_add_4_7 (.A0(n19812), .B0(amdemod_out_d_11__N_2825), 
          .C0(GND_net), .D0(VCC_net), .A1(n19813), .B1(amdemod_out_d_11__N_2822), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17157), .COUT(n17158), .S0(amdemod_out_d_11__N_2410[5]), 
          .S1(amdemod_out_d_11__N_2410[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3585_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_3585_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_3585_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3585_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3585_add_4_5 (.A0(n19810), .B0(amdemod_out_d_11__N_2831), 
          .C0(GND_net), .D0(VCC_net), .A1(n19811), .B1(amdemod_out_d_11__N_2828), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17156), .COUT(n17157), .S0(amdemod_out_d_11__N_2410[3]), 
          .S1(amdemod_out_d_11__N_2410[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3585_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3585_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_3585_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3585_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3585_add_4_3 (.A0(n19809), .B0(square_sum[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19809), .B1(amdemod_out_d_11__N_2834), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17155), .COUT(n17156), .S0(amdemod_out_d_11__N_2410[1]), 
          .S1(amdemod_out_d_11__N_2410[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3585_add_4_3.INIT0 = 16'h666a;
    defparam _add_1_3585_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3585_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3585_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3585_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17155), .S1(amdemod_out_d_11__N_2410[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3585_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3585_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3585_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3585_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_38 (.A0(comb_d7[35]), .B0(comb7[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17154), .S0(comb8_71__N_2137[35]), .S1(cout_adj_6543));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3561_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_36 (.A0(comb_d7[33]), .B0(comb7[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[34]), .B1(comb7[34]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17153), .COUT(n17154), .S0(comb8_71__N_2137[33]), 
          .S1(comb8_71__N_2137[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_34 (.A0(comb_d7[31]), .B0(comb7[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[32]), .B1(comb7[32]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17152), .COUT(n17153), .S0(comb8_71__N_2137[31]), 
          .S1(comb8_71__N_2137[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_32 (.A0(comb_d7[29]), .B0(comb7[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[30]), .B1(comb7[30]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17151), .COUT(n17152), .S0(comb8_71__N_2137[29]), 
          .S1(comb8_71__N_2137[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_30 (.A0(comb_d7[27]), .B0(comb7[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[28]), .B1(comb7[28]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17150), .COUT(n17151), .S0(comb8_71__N_2137[27]), 
          .S1(comb8_71__N_2137[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_28 (.A0(comb_d7[25]), .B0(comb7[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[26]), .B1(comb7[26]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17149), .COUT(n17150), .S0(comb8_71__N_2137[25]), 
          .S1(comb8_71__N_2137[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_26 (.A0(comb_d7[23]), .B0(comb7[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[24]), .B1(comb7[24]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17148), .COUT(n17149), .S0(comb8_71__N_2137[23]), 
          .S1(comb8_71__N_2137[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_24 (.A0(comb_d7[21]), .B0(comb7[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[22]), .B1(comb7[22]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17147), .COUT(n17148), .S0(comb8_71__N_2137[21]), 
          .S1(comb8_71__N_2137[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_22 (.A0(comb_d7[19]), .B0(comb7[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[20]), .B1(comb7[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17146), .COUT(n17147), .S0(comb8_71__N_2137[19]), 
          .S1(comb8_71__N_2137[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_20 (.A0(comb_d7[17]), .B0(comb7[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[18]), .B1(comb7[18]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17145), .COUT(n17146), .S0(comb8_71__N_2137[17]), 
          .S1(comb8_71__N_2137[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_18 (.A0(comb_d7[15]), .B0(comb7[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[16]), .B1(comb7[16]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17144), .COUT(n17145), .S0(comb8_71__N_2137[15]), 
          .S1(comb8_71__N_2137[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_16 (.A0(comb_d7[13]), .B0(comb7[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[14]), .B1(comb7[14]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17143), .COUT(n17144), .S0(comb8_71__N_2137[13]), 
          .S1(comb8_71__N_2137[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_14 (.A0(comb_d7[11]), .B0(comb7[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[12]), .B1(comb7[12]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17142), .COUT(n17143), .S0(comb8_71__N_2137[11]), 
          .S1(comb8_71__N_2137[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_12 (.A0(comb_d7[9]), .B0(comb7[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[10]), .B1(comb7[10]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17141), .COUT(n17142), .S0(comb8_71__N_2137[9]), 
          .S1(comb8_71__N_2137[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_10 (.A0(comb_d7[7]), .B0(comb7[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[8]), .B1(comb7[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17140), .COUT(n17141), .S0(comb8_71__N_2137[7]), 
          .S1(comb8_71__N_2137[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_8 (.A0(comb_d7[5]), .B0(comb7[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[6]), .B1(comb7[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17139), .COUT(n17140), .S0(comb8_71__N_2137[5]), 
          .S1(comb8_71__N_2137[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_6 (.A0(comb_d7[3]), .B0(comb7[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[4]), .B1(comb7[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17138), .COUT(n17139), .S0(comb8_71__N_2137[3]), 
          .S1(comb8_71__N_2137[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_4 (.A0(comb_d7[1]), .B0(comb7[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[2]), .B1(comb7[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17137), .COUT(n17138), .S0(comb8_71__N_2137[1]), 
          .S1(comb8_71__N_2137[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3561_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3561_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[0]), .B1(comb7[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17137), .S1(comb8_71__N_2137[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3561_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3561_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3561_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3561_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_38 (.A0(comb_d8[35]), .B0(comb8[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17136), .S0(comb9_71__N_2209[35]), .S1(cout_adj_6544));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3564_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_36 (.A0(comb_d8[33]), .B0(comb8[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[34]), .B1(comb8[34]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17135), .COUT(n17136), .S0(comb9_71__N_2209[33]), 
          .S1(comb9_71__N_2209[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_34 (.A0(comb_d8[31]), .B0(comb8[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[32]), .B1(comb8[32]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17134), .COUT(n17135), .S0(comb9_71__N_2209[31]), 
          .S1(comb9_71__N_2209[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_32 (.A0(comb_d8[29]), .B0(comb8[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[30]), .B1(comb8[30]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17133), .COUT(n17134), .S0(comb9_71__N_2209[29]), 
          .S1(comb9_71__N_2209[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_30 (.A0(comb_d8[27]), .B0(comb8[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[28]), .B1(comb8[28]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17132), .COUT(n17133), .S0(comb9_71__N_2209[27]), 
          .S1(comb9_71__N_2209[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_28 (.A0(comb_d8[25]), .B0(comb8[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[26]), .B1(comb8[26]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17131), .COUT(n17132), .S0(comb9_71__N_2209[25]), 
          .S1(comb9_71__N_2209[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_26 (.A0(comb_d8[23]), .B0(comb8[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[24]), .B1(comb8[24]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17130), .COUT(n17131), .S0(comb9_71__N_2209[23]), 
          .S1(comb9_71__N_2209[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_24 (.A0(comb_d8[21]), .B0(comb8[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[22]), .B1(comb8[22]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17129), .COUT(n17130), .S0(comb9_71__N_2209[21]), 
          .S1(comb9_71__N_2209[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_22 (.A0(comb_d8[19]), .B0(comb8[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[20]), .B1(comb8[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17128), .COUT(n17129), .S0(comb9_71__N_2209[19]), 
          .S1(comb9_71__N_2209[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_20 (.A0(comb_d8[17]), .B0(comb8[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[18]), .B1(comb8[18]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17127), .COUT(n17128), .S0(comb9_71__N_2209[17]), 
          .S1(comb9_71__N_2209[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_18 (.A0(comb_d8[15]), .B0(comb8[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[16]), .B1(comb8[16]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17126), .COUT(n17127), .S0(comb9_71__N_2209[15]), 
          .S1(comb9_71__N_2209[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_16 (.A0(comb_d8[13]), .B0(comb8[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[14]), .B1(comb8[14]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17125), .COUT(n17126), .S0(comb9_71__N_2209[13]), 
          .S1(comb9_71__N_2209[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_14 (.A0(comb_d8[11]), .B0(comb8[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[12]), .B1(comb8[12]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17124), .COUT(n17125), .S0(comb9_71__N_2209[11]), 
          .S1(comb9_71__N_2209[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_12 (.A0(comb_d8[9]), .B0(comb8[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[10]), .B1(comb8[10]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17123), .COUT(n17124), .S0(comb9_71__N_2209[9]), 
          .S1(comb9_71__N_2209[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_10 (.A0(comb_d8[7]), .B0(comb8[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[8]), .B1(comb8[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17122), .COUT(n17123), .S0(comb9_71__N_2209[7]), 
          .S1(comb9_71__N_2209[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_8 (.A0(comb_d8[5]), .B0(comb8[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[6]), .B1(comb8[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17121), .COUT(n17122), .S0(comb9_71__N_2209[5]), 
          .S1(comb9_71__N_2209[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_6 (.A0(comb_d8[3]), .B0(comb8[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[4]), .B1(comb8[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17120), .COUT(n17121), .S0(comb9_71__N_2209[3]), 
          .S1(comb9_71__N_2209[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_4 (.A0(comb_d8[1]), .B0(comb8[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[2]), .B1(comb8[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17119), .COUT(n17120), .S0(comb9_71__N_2209[1]), 
          .S1(comb9_71__N_2209[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3564_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3564_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[0]), .B1(comb8[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17119), .S1(comb9_71__N_2209[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3564_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3564_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3564_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3564_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_37 (.A0(comb8_adj_6567[70]), .B0(cout_adj_5891), 
          .C0(n81_adj_5629), .D0(n3_adj_5565), .A1(comb8_adj_6567[71]), 
          .B1(cout_adj_5891), .C1(n78_adj_5628), .D1(n2_adj_5564), .CIN(n17117), 
          .S0(comb9_71__N_2209_adj_6592[70]), .S1(comb9_71__N_2209_adj_6592[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_35 (.A0(comb8_adj_6567[68]), .B0(cout_adj_5891), 
          .C0(n87_adj_5631), .D0(n5_adj_5567), .A1(comb8_adj_6567[69]), 
          .B1(cout_adj_5891), .C1(n84_adj_5630), .D1(n4_adj_5566), .CIN(n17116), 
          .COUT(n17117), .S0(comb9_71__N_2209_adj_6592[68]), .S1(comb9_71__N_2209_adj_6592[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_33 (.A0(comb8_adj_6567[66]), .B0(cout_adj_5891), 
          .C0(n93_adj_5633), .D0(n7_adj_5569), .A1(comb8_adj_6567[67]), 
          .B1(cout_adj_5891), .C1(n90_adj_5632), .D1(n6_adj_5568), .CIN(n17115), 
          .COUT(n17116), .S0(comb9_71__N_2209_adj_6592[66]), .S1(comb9_71__N_2209_adj_6592[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_31 (.A0(comb8_adj_6567[64]), .B0(cout_adj_5891), 
          .C0(n99_adj_5635), .D0(n9_adj_5571), .A1(comb8_adj_6567[65]), 
          .B1(cout_adj_5891), .C1(n96_adj_5634), .D1(n8_adj_5570), .CIN(n17114), 
          .COUT(n17115), .S0(comb9_71__N_2209_adj_6592[64]), .S1(comb9_71__N_2209_adj_6592[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_29 (.A0(comb8_adj_6567[62]), .B0(cout_adj_5891), 
          .C0(n105_adj_5637), .D0(n11_adj_5573), .A1(comb8_adj_6567[63]), 
          .B1(cout_adj_5891), .C1(n102_adj_5636), .D1(n10_adj_5572), .CIN(n17113), 
          .COUT(n17114), .S0(comb9_71__N_2209_adj_6592[62]), .S1(comb9_71__N_2209_adj_6592[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_27 (.A0(comb8_adj_6567[60]), .B0(cout_adj_5891), 
          .C0(n111_adj_5639), .D0(n13_adj_5575), .A1(comb8_adj_6567[61]), 
          .B1(cout_adj_5891), .C1(n108_adj_5638), .D1(n12_adj_5574), .CIN(n17112), 
          .COUT(n17113), .S0(comb9_71__N_2209_adj_6592[60]), .S1(comb9_71__N_2209_adj_6592[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_25 (.A0(comb8_adj_6567[58]), .B0(cout_adj_5891), 
          .C0(n117_adj_5641), .D0(n15_adj_5577), .A1(comb8_adj_6567[59]), 
          .B1(cout_adj_5891), .C1(n114_adj_5640), .D1(n14_adj_5576), .CIN(n17111), 
          .COUT(n17112), .S0(comb9_71__N_2209_adj_6592[58]), .S1(comb9_71__N_2209_adj_6592[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_23 (.A0(comb8_adj_6567[56]), .B0(cout_adj_5891), 
          .C0(n123_adj_5643), .D0(n17_adj_5579), .A1(comb8_adj_6567[57]), 
          .B1(cout_adj_5891), .C1(n120_adj_5642), .D1(n16_adj_5578), .CIN(n17110), 
          .COUT(n17111), .S0(comb9_71__N_2209_adj_6592[56]), .S1(comb9_71__N_2209_adj_6592[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_21 (.A0(comb8_adj_6567[54]), .B0(cout_adj_5891), 
          .C0(n129_adj_5645), .D0(n19_adj_5581), .A1(comb8_adj_6567[55]), 
          .B1(cout_adj_5891), .C1(n126_adj_5644), .D1(n18_adj_5580), .CIN(n17109), 
          .COUT(n17110), .S0(comb9_71__N_2209_adj_6592[54]), .S1(comb9_71__N_2209_adj_6592[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_19 (.A0(comb8_adj_6567[52]), .B0(cout_adj_5891), 
          .C0(n135_adj_5647), .D0(n21_adj_5583), .A1(comb8_adj_6567[53]), 
          .B1(cout_adj_5891), .C1(n132_adj_5646), .D1(n20_adj_5582), .CIN(n17108), 
          .COUT(n17109), .S0(comb9_71__N_2209_adj_6592[52]), .S1(comb9_71__N_2209_adj_6592[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_17 (.A0(comb8_adj_6567[50]), .B0(cout_adj_5891), 
          .C0(n141_adj_5649), .D0(n23_adj_5585), .A1(comb8_adj_6567[51]), 
          .B1(cout_adj_5891), .C1(n138_adj_5648), .D1(n22_adj_5584), .CIN(n17107), 
          .COUT(n17108), .S0(comb9_71__N_2209_adj_6592[50]), .S1(comb9_71__N_2209_adj_6592[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_15 (.A0(comb8_adj_6567[48]), .B0(cout_adj_5891), 
          .C0(n147_adj_5651), .D0(n25_adj_5587), .A1(comb8_adj_6567[49]), 
          .B1(cout_adj_5891), .C1(n144_adj_5650), .D1(n24_adj_5586), .CIN(n17106), 
          .COUT(n17107), .S0(comb9_71__N_2209_adj_6592[48]), .S1(comb9_71__N_2209_adj_6592[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_13 (.A0(comb8_adj_6567[46]), .B0(cout_adj_5891), 
          .C0(n153_adj_5653), .D0(n27_adj_5589), .A1(comb8_adj_6567[47]), 
          .B1(cout_adj_5891), .C1(n150_adj_5652), .D1(n26_adj_5588), .CIN(n17105), 
          .COUT(n17106), .S0(comb9_71__N_2209_adj_6592[46]), .S1(comb9_71__N_2209_adj_6592[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_11 (.A0(comb8_adj_6567[44]), .B0(cout_adj_5891), 
          .C0(n159_adj_5655), .D0(n29_adj_5591), .A1(comb8_adj_6567[45]), 
          .B1(cout_adj_5891), .C1(n156_adj_5654), .D1(n28_adj_5590), .CIN(n17104), 
          .COUT(n17105), .S0(comb9_71__N_2209_adj_6592[44]), .S1(comb9_71__N_2209_adj_6592[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_9 (.A0(comb8_adj_6567[42]), .B0(cout_adj_5891), 
          .C0(n165_adj_5657), .D0(n31_adj_5593), .A1(comb8_adj_6567[43]), 
          .B1(cout_adj_5891), .C1(n162_adj_5656), .D1(n30_adj_5592), .CIN(n17103), 
          .COUT(n17104), .S0(comb9_71__N_2209_adj_6592[42]), .S1(comb9_71__N_2209_adj_6592[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_7 (.A0(comb8_adj_6567[40]), .B0(cout_adj_5891), 
          .C0(n171_adj_5659), .D0(n33_adj_5595), .A1(comb8_adj_6567[41]), 
          .B1(cout_adj_5891), .C1(n168_adj_5658), .D1(n32_adj_5594), .CIN(n17102), 
          .COUT(n17103), .S0(comb9_71__N_2209_adj_6592[40]), .S1(comb9_71__N_2209_adj_6592[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_5 (.A0(comb8_adj_6567[38]), .B0(cout_adj_5891), 
          .C0(n177_adj_5661), .D0(n35_adj_5597), .A1(comb8_adj_6567[39]), 
          .B1(cout_adj_5891), .C1(n174_adj_5660), .D1(n34_adj_5596), .CIN(n17101), 
          .COUT(n17102), .S0(comb9_71__N_2209_adj_6592[38]), .S1(comb9_71__N_2209_adj_6592[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_3 (.A0(comb8_adj_6567[36]), .B0(cout_adj_5891), 
          .C0(n183_adj_5663), .D0(n37_adj_5599), .A1(comb8_adj_6567[37]), 
          .B1(cout_adj_5891), .C1(n180_adj_5662), .D1(n36_adj_5598), .CIN(n17100), 
          .COUT(n17101), .S0(comb9_71__N_2209_adj_6592[36]), .S1(comb9_71__N_2209_adj_6592[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3654_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3654_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3654_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5891), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17100));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3654_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3654_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3654_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3654_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_63 (.A0(\phase_increment[0] [62]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [63]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17095), .S0(phase_increment_1__63__N_21[62]), 
          .S1(phase_increment_1__63__N_21[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_63.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_63.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_63.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_63.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_61 (.A0(\phase_increment[0] [60]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [61]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17094), .COUT(n17095), .S0(phase_increment_1__63__N_21[60]), 
          .S1(phase_increment_1__63__N_21[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_61.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_61.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_61.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_59 (.A0(\phase_increment[0] [58]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [59]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17093), .COUT(n17094), .S0(phase_increment_1__63__N_21[58]), 
          .S1(phase_increment_1__63__N_21[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_59.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_59.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_57 (.A0(\phase_increment[0] [56]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [57]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17092), .COUT(n17093), .S0(phase_increment_1__63__N_21[56]), 
          .S1(phase_increment_1__63__N_21[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_57.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_57.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_55 (.A0(\phase_increment[0] [54]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [55]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17091), .COUT(n17092), .S0(phase_increment_1__63__N_21[54]), 
          .S1(phase_increment_1__63__N_21[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_55.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_55.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_53 (.A0(\phase_increment[0] [52]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [53]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17090), .COUT(n17091), .S0(phase_increment_1__63__N_21[52]), 
          .S1(phase_increment_1__63__N_21[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_53.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_53.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_51 (.A0(\phase_increment[0] [50]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [51]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17089), .COUT(n17090), .S0(phase_increment_1__63__N_21[50]), 
          .S1(phase_increment_1__63__N_21[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_51.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_51.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_49 (.A0(\phase_increment[0] [48]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [49]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17088), .COUT(n17089), .S0(phase_increment_1__63__N_21[48]), 
          .S1(phase_increment_1__63__N_21[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_49.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_49.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_47 (.A0(\phase_increment[0] [46]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [47]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17087), .COUT(n17088), .S0(phase_increment_1__63__N_21[46]), 
          .S1(phase_increment_1__63__N_21[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_47.INIT0 = 16'h555f;
    defparam _add_1_3492_add_4_47.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_45 (.A0(\phase_increment[0] [44]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [45]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17086), .COUT(n17087), .S0(phase_increment_1__63__N_21[44]), 
          .S1(phase_increment_1__63__N_21[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_45.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_45.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_43 (.A0(\phase_increment[0] [42]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [43]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17085), .COUT(n17086), .S0(phase_increment_1__63__N_21[42]), 
          .S1(phase_increment_1__63__N_21[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_43.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_43.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_41 (.A0(\phase_increment[0] [40]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [41]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17084), .COUT(n17085), .S0(phase_increment_1__63__N_21[40]), 
          .S1(phase_increment_1__63__N_21[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_41.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_41.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_39 (.A0(\phase_increment[0] [38]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [39]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17083), .COUT(n17084), .S0(phase_increment_1__63__N_21[38]), 
          .S1(phase_increment_1__63__N_21[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_39.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_39.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_37 (.A0(\phase_increment[0] [36]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [37]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17082), .COUT(n17083), .S0(phase_increment_1__63__N_21[36]), 
          .S1(phase_increment_1__63__N_21[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_37.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_37.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_35 (.A0(\phase_increment[0] [34]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [35]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17081), .COUT(n17082), .S0(phase_increment_1__63__N_21[34]), 
          .S1(phase_increment_1__63__N_21[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_35.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_35.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_33 (.A0(\phase_increment[0] [32]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [33]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17080), .COUT(n17081), .S0(phase_increment_1__63__N_21[32]), 
          .S1(phase_increment_1__63__N_21[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_33.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_33.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_31 (.A0(\phase_increment[0] [30]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [31]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17079), .COUT(n17080), .S0(phase_increment_1__63__N_21[30]), 
          .S1(phase_increment_1__63__N_21[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_31.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_31.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_29 (.A0(\phase_increment[0] [28]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [29]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17078), .COUT(n17079), .S0(phase_increment_1__63__N_21[28]), 
          .S1(phase_increment_1__63__N_21[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_29.INIT0 = 16'h555f;
    defparam _add_1_3492_add_4_29.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_27 (.A0(\phase_increment[0] [26]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [27]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17077), .COUT(n17078), .S0(phase_increment_1__63__N_21[26]), 
          .S1(phase_increment_1__63__N_21[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_27.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_27.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_25 (.A0(\phase_increment[0] [24]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [25]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17076), .COUT(n17077), .S0(phase_increment_1__63__N_21[24]), 
          .S1(phase_increment_1__63__N_21[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_25.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_25.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_23 (.A0(\phase_increment[0] [22]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [23]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17075), .COUT(n17076), .S0(phase_increment_1__63__N_21[22]), 
          .S1(phase_increment_1__63__N_21[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_23.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_23.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_21 (.A0(\phase_increment[0] [20]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [21]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17074), .COUT(n17075), .S0(phase_increment_1__63__N_21[20]), 
          .S1(phase_increment_1__63__N_21[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_21.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_21.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_19 (.A0(\phase_increment[0] [18]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [19]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17073), .COUT(n17074), .S0(phase_increment_1__63__N_21[18]), 
          .S1(phase_increment_1__63__N_21[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_19.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_17 (.A0(\phase_increment[0] [16]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [17]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17072), .COUT(n17073), .S0(phase_increment_1__63__N_21[16]), 
          .S1(phase_increment_1__63__N_21[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_17.INIT0 = 16'h555f;
    defparam _add_1_3492_add_4_17.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_15 (.A0(\phase_increment[0] [14]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [15]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17071), .COUT(n17072), .S0(phase_increment_1__63__N_21[14]), 
          .S1(phase_increment_1__63__N_21[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_15.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_13 (.A0(\phase_increment[0] [12]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [13]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17070), .COUT(n17071), .S0(phase_increment_1__63__N_21[12]), 
          .S1(phase_increment_1__63__N_21[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3492_add_4_13.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_11 (.A0(\phase_increment[0] [10]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [11]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17069), .COUT(n17070), .S0(phase_increment_1__63__N_21[10]), 
          .S1(phase_increment_1__63__N_21[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_11.INIT0 = 16'h555f;
    defparam _add_1_3492_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_9 (.A0(\phase_increment[0] [8]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [9]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17068), .COUT(n17069), .S0(phase_increment_1__63__N_21[8]), 
          .S1(phase_increment_1__63__N_21[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_9.INIT0 = 16'h555f;
    defparam _add_1_3492_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_7 (.A0(\phase_increment[0] [6]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [7]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17067), .COUT(n17068), .S0(phase_increment_1__63__N_21[6]), 
          .S1(phase_increment_1__63__N_21[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_7.INIT0 = 16'h555f;
    defparam _add_1_3492_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_3492_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_5 (.A0(\phase_increment[0] [4]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [5]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17066), .COUT(n17067), .S0(phase_increment_1__63__N_21[4]), 
          .S1(phase_increment_1__63__N_21[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_5.INIT0 = 16'h555f;
    defparam _add_1_3492_add_4_5.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_3 (.A0(phase_increment_1__63__N_17[2]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_increment_1__63__N_17[3]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17065), .COUT(n17066), 
          .S0(phase_increment_1__63__N_21[2]), .S1(phase_increment_1__63__N_21[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_3.INIT0 = 16'h555f;
    defparam _add_1_3492_add_4_3.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3492_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_increment_1__63__N_17[1]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .COUT(n17065), .S1(phase_increment_1__63__N_21[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(287[40:78])
    defparam _add_1_3492_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3492_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3492_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3492_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3789_add_4_14 (.A0(amdemod_out_d_11__N_2363), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17056), .S0(amdemod_out_d_11__N_2369[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3789_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_3789_add_4_14.INIT1 = 16'h0000;
    defparam _add_1_3789_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3789_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3789_add_4_12 (.A0(amdemod_out_d_11__N_2501), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2363), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17055), .COUT(n17056), .S0(amdemod_out_d_11__N_2369[9]), 
          .S1(amdemod_out_d_11__N_2369[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3789_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_3789_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_3789_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3789_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3789_add_4_10 (.A0(amdemod_out_d_11__N_2507), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2504), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17054), .COUT(n17055), .S0(amdemod_out_d_11__N_2369[7]), 
          .S1(amdemod_out_d_11__N_2369[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3789_add_4_10.INIT0 = 16'h555f;
    defparam _add_1_3789_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_3789_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3789_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3789_add_4_8 (.A0(amdemod_out_d_11__N_2513), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2510), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17053), .COUT(n17054), .S0(amdemod_out_d_11__N_2369[5]), 
          .S1(amdemod_out_d_11__N_2369[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3789_add_4_8.INIT0 = 16'h555f;
    defparam _add_1_3789_add_4_8.INIT1 = 16'h555f;
    defparam _add_1_3789_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3789_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3789_add_4_6 (.A0(square_sum[25]), .B0(n19824), .C0(n45_adj_6287), 
          .D0(n13876), .A1(amdemod_out_d_11__N_2358[5]), .B1(square_sum[25]), 
          .C1(n42_adj_6286), .D1(n13878), .CIN(n17052), .COUT(n17053), 
          .S0(amdemod_out_d_11__N_2369[3]), .S1(amdemod_out_d_11__N_2369[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3789_add_4_6.INIT0 = 16'he4b1;
    defparam _add_1_3789_add_4_6.INIT1 = 16'h596a;
    defparam _add_1_3789_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3789_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3789_add_4_4 (.A0(amdemod_out_d_11__N_2363), .B0(square_sum[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2363), .B1(square_sum[25]), 
          .C1(n48_adj_6288), .D1(n13815), .CIN(n17051), .COUT(n17052), 
          .S0(amdemod_out_d_11__N_2369[1]), .S1(amdemod_out_d_11__N_2369[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3789_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3789_add_4_4.INIT1 = 16'h596a;
    defparam _add_1_3789_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3789_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3789_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[18]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17051), .S1(amdemod_out_d_11__N_2369[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3789_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3789_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3789_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3789_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_65 (.A0(\phase_increment[0] [63]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17050), .S0(phase_increment_1__63__N_19[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_65.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_65.INIT1 = 16'h0000;
    defparam _add_1_3498_add_4_65.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_65.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_63 (.A0(\phase_increment[0] [61]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [62]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17049), .COUT(n17050), .S0(phase_increment_1__63__N_19[61]), 
          .S1(phase_increment_1__63__N_19[62]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_63.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_63.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_63.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_63.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_61 (.A0(\phase_increment[0] [59]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [60]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17048), .COUT(n17049), .S0(phase_increment_1__63__N_19[59]), 
          .S1(phase_increment_1__63__N_19[60]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_61.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_61.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_61.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_59 (.A0(\phase_increment[0] [57]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [58]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17047), .COUT(n17048), .S0(phase_increment_1__63__N_19[57]), 
          .S1(phase_increment_1__63__N_19[58]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_59.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_59.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_57 (.A0(\phase_increment[0] [55]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [56]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17046), .COUT(n17047), .S0(phase_increment_1__63__N_19[55]), 
          .S1(phase_increment_1__63__N_19[56]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_57.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_57.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_55 (.A0(\phase_increment[0] [53]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [54]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17045), .COUT(n17046), .S0(phase_increment_1__63__N_19[53]), 
          .S1(phase_increment_1__63__N_19[54]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_55.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_55.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_53 (.A0(\phase_increment[0] [51]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [52]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17044), .COUT(n17045), .S0(phase_increment_1__63__N_19[51]), 
          .S1(phase_increment_1__63__N_19[52]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_53.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_53.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_51 (.A0(\phase_increment[0] [49]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [50]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17043), .COUT(n17044), .S0(phase_increment_1__63__N_19[49]), 
          .S1(phase_increment_1__63__N_19[50]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_51.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_51.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_49 (.A0(\phase_increment[0] [47]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [48]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17042), .COUT(n17043), .S0(phase_increment_1__63__N_19[47]), 
          .S1(phase_increment_1__63__N_19[48]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_49.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_49.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_47 (.A0(\phase_increment[0] [45]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [46]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17041), .COUT(n17042), .S0(phase_increment_1__63__N_19[45]), 
          .S1(phase_increment_1__63__N_19[46]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_45 (.A0(\phase_increment[0] [43]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [44]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17040), .COUT(n17041), .S0(phase_increment_1__63__N_19[43]), 
          .S1(phase_increment_1__63__N_19[44]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_45.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_45.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_43 (.A0(\phase_increment[0] [41]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [42]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17039), .COUT(n17040), .S0(phase_increment_1__63__N_19[41]), 
          .S1(phase_increment_1__63__N_19[42]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_43.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_43.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_41 (.A0(\phase_increment[0] [39]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [40]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17038), .COUT(n17039), .S0(phase_increment_1__63__N_19[39]), 
          .S1(phase_increment_1__63__N_19[40]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_41.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_39 (.A0(\phase_increment[0] [37]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [38]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17037), .COUT(n17038), .S0(phase_increment_1__63__N_19[37]), 
          .S1(phase_increment_1__63__N_19[38]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_39.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_39.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_37 (.A0(\phase_increment[0] [35]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [36]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17036), .COUT(n17037), .S0(phase_increment_1__63__N_19[35]), 
          .S1(phase_increment_1__63__N_19[36]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_37.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_37.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_35 (.A0(\phase_increment[0] [33]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [34]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17035), .COUT(n17036), .S0(phase_increment_1__63__N_19[33]), 
          .S1(phase_increment_1__63__N_19[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_35.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_33 (.A0(\phase_increment[0] [31]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [32]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17034), .COUT(n17035), .S0(phase_increment_1__63__N_19[31]), 
          .S1(phase_increment_1__63__N_19[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_31 (.A0(\phase_increment[0] [29]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [30]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17033), .COUT(n17034), .S0(phase_increment_1__63__N_19[29]), 
          .S1(phase_increment_1__63__N_19[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_31.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_29 (.A0(\phase_increment[0] [27]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [28]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17032), .COUT(n17033), .S0(phase_increment_1__63__N_19[27]), 
          .S1(phase_increment_1__63__N_19[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_29.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_29.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_27 (.A0(\phase_increment[0] [25]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [26]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17031), .COUT(n17032), .S0(phase_increment_1__63__N_19[25]), 
          .S1(phase_increment_1__63__N_19[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_27.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_25 (.A0(\phase_increment[0] [23]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [24]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17030), .COUT(n17031), .S0(phase_increment_1__63__N_19[23]), 
          .S1(phase_increment_1__63__N_19[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_25.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_25.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_23 (.A0(\phase_increment[0] [21]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [22]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17029), .COUT(n17030), .S0(phase_increment_1__63__N_19[21]), 
          .S1(phase_increment_1__63__N_19[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_23.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_21 (.A0(\phase_increment[0] [19]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [20]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17028), .COUT(n17029), .S0(phase_increment_1__63__N_19[19]), 
          .S1(phase_increment_1__63__N_19[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_21.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_19 (.A0(\phase_increment[0] [17]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [18]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17027), .COUT(n17028), .S0(phase_increment_1__63__N_19[17]), 
          .S1(phase_increment_1__63__N_19[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_19.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_17 (.A0(\phase_increment[0] [15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [16]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17026), .COUT(n17027), .S0(phase_increment_1__63__N_19[15]), 
          .S1(phase_increment_1__63__N_19[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_17.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_17.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_15 (.A0(\phase_increment[0] [13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17025), .COUT(n17026), .S0(phase_increment_1__63__N_19[13]), 
          .S1(phase_increment_1__63__N_19[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_15.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_13 (.A0(\phase_increment[0] [11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17024), .COUT(n17025), .S0(phase_increment_1__63__N_19[11]), 
          .S1(phase_increment_1__63__N_19[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_13.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_11 (.A0(\phase_increment[0] [9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17023), .COUT(n17024), .S0(phase_increment_1__63__N_19[9]), 
          .S1(phase_increment_1__63__N_19[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_11.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_11.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_9 (.A0(\phase_increment[0] [7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17022), .COUT(n17023), .S0(phase_increment_1__63__N_19[7]), 
          .S1(phase_increment_1__63__N_19[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_9.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_7 (.A0(\phase_increment[0] [5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17021), .COUT(n17022), .S0(phase_increment_1__63__N_19[5]), 
          .S1(phase_increment_1__63__N_19[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_7.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_5 (.A0(phase_increment_1__63__N_17[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17020), .COUT(n17021), .S0(phase_increment_1__63__N_19[3]), 
          .S1(phase_increment_1__63__N_19[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_3498_add_4_5.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_3 (.A0(phase_increment_1__63__N_17[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_increment_1__63__N_17[2]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17019), .COUT(n17020), 
          .S0(phase_increment_1__63__N_19[1]), .S1(phase_increment_1__63__N_19[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_3.INIT0 = 16'h555f;
    defparam _add_1_3498_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_3498_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3498_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_increment_1__63__N_21[0]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .COUT(n17019), .S1(phase_increment_1__63__N_19[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(285[40:78])
    defparam _add_1_3498_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3498_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3498_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3498_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_38 (.A0(integrator_d_tmp[35]), .B0(integrator_tmp[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17018), .S0(comb6_71__N_1993[35]), .S1(cout_adj_5271));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3528_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_36 (.A0(integrator_d_tmp[33]), .B0(integrator_tmp[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[34]), .B1(integrator_tmp[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17017), .COUT(n17018), .S0(comb6_71__N_1993[33]), 
          .S1(comb6_71__N_1993[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_34 (.A0(integrator_d_tmp[31]), .B0(integrator_tmp[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[32]), .B1(integrator_tmp[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17016), .COUT(n17017), .S0(comb6_71__N_1993[31]), 
          .S1(comb6_71__N_1993[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_32 (.A0(integrator_d_tmp[29]), .B0(integrator_tmp[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[30]), .B1(integrator_tmp[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17015), .COUT(n17016), .S0(comb6_71__N_1993[29]), 
          .S1(comb6_71__N_1993[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_30 (.A0(integrator_d_tmp[27]), .B0(integrator_tmp[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[28]), .B1(integrator_tmp[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17014), .COUT(n17015), .S0(comb6_71__N_1993[27]), 
          .S1(comb6_71__N_1993[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_28 (.A0(integrator_d_tmp[25]), .B0(integrator_tmp[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[26]), .B1(integrator_tmp[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17013), .COUT(n17014), .S0(comb6_71__N_1993[25]), 
          .S1(comb6_71__N_1993[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_26 (.A0(integrator_d_tmp[23]), .B0(integrator_tmp[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[24]), .B1(integrator_tmp[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17012), .COUT(n17013), .S0(comb6_71__N_1993[23]), 
          .S1(comb6_71__N_1993[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_24 (.A0(integrator_d_tmp[21]), .B0(integrator_tmp[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[22]), .B1(integrator_tmp[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17011), .COUT(n17012), .S0(comb6_71__N_1993[21]), 
          .S1(comb6_71__N_1993[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_22 (.A0(integrator_d_tmp[19]), .B0(integrator_tmp[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[20]), .B1(integrator_tmp[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17010), .COUT(n17011), .S0(comb6_71__N_1993[19]), 
          .S1(comb6_71__N_1993[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_20 (.A0(integrator_d_tmp[17]), .B0(integrator_tmp[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[18]), .B1(integrator_tmp[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17009), .COUT(n17010), .S0(comb6_71__N_1993[17]), 
          .S1(comb6_71__N_1993[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_18 (.A0(integrator_d_tmp[15]), .B0(integrator_tmp[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[16]), .B1(integrator_tmp[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17008), .COUT(n17009), .S0(comb6_71__N_1993[15]), 
          .S1(comb6_71__N_1993[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_16 (.A0(integrator_d_tmp[13]), .B0(integrator_tmp[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[14]), .B1(integrator_tmp[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17007), .COUT(n17008), .S0(comb6_71__N_1993[13]), 
          .S1(comb6_71__N_1993[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_14 (.A0(integrator_d_tmp[11]), .B0(integrator_tmp[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[12]), .B1(integrator_tmp[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17006), .COUT(n17007), .S0(comb6_71__N_1993[11]), 
          .S1(comb6_71__N_1993[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_12 (.A0(integrator_d_tmp[9]), .B0(integrator_tmp[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[10]), .B1(integrator_tmp[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17005), .COUT(n17006), .S0(comb6_71__N_1993[9]), 
          .S1(comb6_71__N_1993[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_10 (.A0(integrator_d_tmp[7]), .B0(integrator_tmp[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[8]), .B1(integrator_tmp[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17004), .COUT(n17005), .S0(comb6_71__N_1993[7]), 
          .S1(comb6_71__N_1993[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_8 (.A0(integrator_d_tmp[5]), .B0(integrator_tmp[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[6]), .B1(integrator_tmp[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17003), .COUT(n17004), .S0(comb6_71__N_1993[5]), 
          .S1(comb6_71__N_1993[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_6 (.A0(integrator_d_tmp[3]), .B0(integrator_tmp[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[4]), .B1(integrator_tmp[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17002), .COUT(n17003), .S0(comb6_71__N_1993[3]), 
          .S1(comb6_71__N_1993[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_4 (.A0(integrator_d_tmp[1]), .B0(integrator_tmp[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[2]), .B1(integrator_tmp[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17001), .COUT(n17002), .S0(comb6_71__N_1993[1]), 
          .S1(comb6_71__N_1993[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3528_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3528_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator_d_tmp[0]), .B1(integrator_tmp[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n17001), .S1(comb6_71__N_1993[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3528_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3528_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3528_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3528_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_38 (.A0(integrator4[71]), .B0(integrator3[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17000), .S0(n78_adj_6093));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3546_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_36 (.A0(integrator4[69]), .B0(integrator3[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[70]), .B1(integrator3[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16999), .COUT(n17000), .S0(n84_adj_6095), 
          .S1(n81_adj_6094));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_34 (.A0(integrator4[67]), .B0(integrator3[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[68]), .B1(integrator3[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16998), .COUT(n16999), .S0(n90_adj_6097), 
          .S1(n87_adj_6096));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_32 (.A0(integrator4[65]), .B0(integrator3[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[66]), .B1(integrator3[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16997), .COUT(n16998), .S0(n96_adj_6099), 
          .S1(n93_adj_6098));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_30 (.A0(integrator4[63]), .B0(integrator3[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[64]), .B1(integrator3[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16996), .COUT(n16997), .S0(n102_adj_6101), 
          .S1(n99_adj_6100));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_28 (.A0(integrator4[61]), .B0(integrator3[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[62]), .B1(integrator3[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16995), .COUT(n16996), .S0(n108_adj_6103), 
          .S1(n105_adj_6102));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_26 (.A0(integrator4[59]), .B0(integrator3[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[60]), .B1(integrator3[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16994), .COUT(n16995), .S0(n114_adj_6105), 
          .S1(n111_adj_6104));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_24 (.A0(integrator4[57]), .B0(integrator3[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[58]), .B1(integrator3[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16993), .COUT(n16994), .S0(n120_adj_6107), 
          .S1(n117_adj_6106));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_22 (.A0(integrator4[55]), .B0(integrator3[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[56]), .B1(integrator3[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16992), .COUT(n16993), .S0(n126_adj_6109), 
          .S1(n123_adj_6108));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_20 (.A0(integrator4[53]), .B0(integrator3[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[54]), .B1(integrator3[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16991), .COUT(n16992), .S0(n132_adj_6111), 
          .S1(n129_adj_6110));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_18 (.A0(integrator4[51]), .B0(integrator3[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[52]), .B1(integrator3[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16990), .COUT(n16991), .S0(n138_adj_6113), 
          .S1(n135_adj_6112));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_16 (.A0(integrator4[49]), .B0(integrator3[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[50]), .B1(integrator3[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16989), .COUT(n16990), .S0(n144_adj_6115), 
          .S1(n141_adj_6114));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_14 (.A0(integrator4[47]), .B0(integrator3[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[48]), .B1(integrator3[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16988), .COUT(n16989), .S0(n150_adj_6117), 
          .S1(n147_adj_6116));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_12 (.A0(integrator4[45]), .B0(integrator3[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[46]), .B1(integrator3[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16987), .COUT(n16988), .S0(n156_adj_6119), 
          .S1(n153_adj_6118));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_10 (.A0(integrator4[43]), .B0(integrator3[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[44]), .B1(integrator3[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16986), .COUT(n16987), .S0(n162_adj_6121), 
          .S1(n159_adj_6120));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_8 (.A0(integrator4[41]), .B0(integrator3[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[42]), .B1(integrator3[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16985), .COUT(n16986), .S0(n168_adj_6123), 
          .S1(n165_adj_6122));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_6 (.A0(integrator4[39]), .B0(integrator3[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[40]), .B1(integrator3[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16984), .COUT(n16985), .S0(n174_adj_6125), 
          .S1(n171_adj_6124));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_4 (.A0(integrator4[37]), .B0(integrator3[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[38]), .B1(integrator3[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16983), .COUT(n16984), .S0(n180_adj_6127), 
          .S1(n177_adj_6126));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3546_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3546_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator4[36]), .B1(integrator3[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16983), .S1(n183_adj_6128));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3546_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3546_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3546_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3546_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3531_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16982), .S0(n28));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3531_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3531_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_3531_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3531_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3531_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16981), .COUT(n16982), .S0(n34), .S1(n31));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3531_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3531_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3531_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3531_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3531_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16980), .COUT(n16981), .S0(n40), .S1(n37_adj_5270));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3531_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_3531_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_3531_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3531_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3531_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16979), .COUT(n16980), .S0(n46), .S1(n43));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3531_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_3531_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_3531_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3531_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3531_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16978), .COUT(n16979), .S0(n52), .S1(n49));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3531_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_3531_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_3531_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3531_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3531_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16977), .COUT(n16978), .S0(n58), .S1(n55));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3531_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_3531_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_3531_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3531_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3531_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16977), .S1(n61));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3531_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3531_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3531_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3531_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_38 (.A0(comb_d8_adj_6568[71]), .B0(comb8_adj_6567[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16976), .S0(n78_adj_5628));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3678_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_36 (.A0(comb_d8_adj_6568[69]), .B0(comb8_adj_6567[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[70]), .B1(comb8_adj_6567[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16975), .COUT(n16976), .S0(n84_adj_5630), 
          .S1(n81_adj_5629));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_34 (.A0(comb_d8_adj_6568[67]), .B0(comb8_adj_6567[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[68]), .B1(comb8_adj_6567[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16974), .COUT(n16975), .S0(n90_adj_5632), 
          .S1(n87_adj_5631));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_32 (.A0(comb_d8_adj_6568[65]), .B0(comb8_adj_6567[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[66]), .B1(comb8_adj_6567[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16973), .COUT(n16974), .S0(n96_adj_5634), 
          .S1(n93_adj_5633));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_30 (.A0(comb_d8_adj_6568[63]), .B0(comb8_adj_6567[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[64]), .B1(comb8_adj_6567[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16972), .COUT(n16973), .S0(n102_adj_5636), 
          .S1(n99_adj_5635));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_28 (.A0(comb_d8_adj_6568[61]), .B0(comb8_adj_6567[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[62]), .B1(comb8_adj_6567[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16971), .COUT(n16972), .S0(n108_adj_5638), 
          .S1(n105_adj_5637));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_26 (.A0(comb_d8_adj_6568[59]), .B0(comb8_adj_6567[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[60]), .B1(comb8_adj_6567[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16970), .COUT(n16971), .S0(n114_adj_5640), 
          .S1(n111_adj_5639));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_24 (.A0(comb_d8_adj_6568[57]), .B0(comb8_adj_6567[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[58]), .B1(comb8_adj_6567[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16969), .COUT(n16970), .S0(n120_adj_5642), 
          .S1(n117_adj_5641));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_22 (.A0(comb_d8_adj_6568[55]), .B0(comb8_adj_6567[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[56]), .B1(comb8_adj_6567[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16968), .COUT(n16969), .S0(n126_adj_5644), 
          .S1(n123_adj_5643));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_20 (.A0(comb_d8_adj_6568[53]), .B0(comb8_adj_6567[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[54]), .B1(comb8_adj_6567[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16967), .COUT(n16968), .S0(n132_adj_5646), 
          .S1(n129_adj_5645));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_18 (.A0(comb_d8_adj_6568[51]), .B0(comb8_adj_6567[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[52]), .B1(comb8_adj_6567[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16966), .COUT(n16967), .S0(n138_adj_5648), 
          .S1(n135_adj_5647));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_16 (.A0(comb_d8_adj_6568[49]), .B0(comb8_adj_6567[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[50]), .B1(comb8_adj_6567[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16965), .COUT(n16966), .S0(n144_adj_5650), 
          .S1(n141_adj_5649));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_14 (.A0(comb_d8_adj_6568[47]), .B0(comb8_adj_6567[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[48]), .B1(comb8_adj_6567[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16964), .COUT(n16965), .S0(n150_adj_5652), 
          .S1(n147_adj_5651));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_12 (.A0(comb_d8_adj_6568[45]), .B0(comb8_adj_6567[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[46]), .B1(comb8_adj_6567[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16963), .COUT(n16964), .S0(n156_adj_5654), 
          .S1(n153_adj_5653));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_10 (.A0(comb_d8_adj_6568[43]), .B0(comb8_adj_6567[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[44]), .B1(comb8_adj_6567[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16962), .COUT(n16963), .S0(n162_adj_5656), 
          .S1(n159_adj_5655));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_8 (.A0(comb_d8_adj_6568[41]), .B0(comb8_adj_6567[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[42]), .B1(comb8_adj_6567[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16961), .COUT(n16962), .S0(n168_adj_5658), 
          .S1(n165_adj_5657));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_6 (.A0(comb_d8_adj_6568[39]), .B0(comb8_adj_6567[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[40]), .B1(comb8_adj_6567[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16960), .COUT(n16961), .S0(n174_adj_5660), 
          .S1(n171_adj_5659));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_4 (.A0(comb_d8_adj_6568[37]), .B0(comb8_adj_6567[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6568[38]), .B1(comb8_adj_6567[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16959), .COUT(n16960), .S0(n180_adj_5662), 
          .S1(n177_adj_5661));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3678_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3678_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8_adj_6568[36]), .B1(comb8_adj_6567[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16959), .S1(n183_adj_5663));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3678_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3678_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3678_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3678_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_38 (.A0(comb_d6[35]), .B0(comb6[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16958), .S0(comb7_71__N_2065[35]), .S1(cout_adj_6129));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3549_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_36 (.A0(comb_d6[33]), .B0(comb6[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[34]), .B1(comb6[34]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16957), .COUT(n16958), .S0(comb7_71__N_2065[33]), 
          .S1(comb7_71__N_2065[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_34 (.A0(comb_d6[31]), .B0(comb6[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[32]), .B1(comb6[32]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16956), .COUT(n16957), .S0(comb7_71__N_2065[31]), 
          .S1(comb7_71__N_2065[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_32 (.A0(comb_d6[29]), .B0(comb6[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[30]), .B1(comb6[30]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16955), .COUT(n16956), .S0(comb7_71__N_2065[29]), 
          .S1(comb7_71__N_2065[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_30 (.A0(comb_d6[27]), .B0(comb6[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[28]), .B1(comb6[28]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16954), .COUT(n16955), .S0(comb7_71__N_2065[27]), 
          .S1(comb7_71__N_2065[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_28 (.A0(comb_d6[25]), .B0(comb6[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[26]), .B1(comb6[26]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16953), .COUT(n16954), .S0(comb7_71__N_2065[25]), 
          .S1(comb7_71__N_2065[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_26 (.A0(comb_d6[23]), .B0(comb6[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[24]), .B1(comb6[24]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16952), .COUT(n16953), .S0(comb7_71__N_2065[23]), 
          .S1(comb7_71__N_2065[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_24 (.A0(comb_d6[21]), .B0(comb6[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[22]), .B1(comb6[22]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16951), .COUT(n16952), .S0(comb7_71__N_2065[21]), 
          .S1(comb7_71__N_2065[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_22 (.A0(comb_d6[19]), .B0(comb6[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[20]), .B1(comb6[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16950), .COUT(n16951), .S0(comb7_71__N_2065[19]), 
          .S1(comb7_71__N_2065[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_20 (.A0(comb_d6[17]), .B0(comb6[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[18]), .B1(comb6[18]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16949), .COUT(n16950), .S0(comb7_71__N_2065[17]), 
          .S1(comb7_71__N_2065[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_18 (.A0(comb_d6[15]), .B0(comb6[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[16]), .B1(comb6[16]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16948), .COUT(n16949), .S0(comb7_71__N_2065[15]), 
          .S1(comb7_71__N_2065[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_16 (.A0(comb_d6[13]), .B0(comb6[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[14]), .B1(comb6[14]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16947), .COUT(n16948), .S0(comb7_71__N_2065[13]), 
          .S1(comb7_71__N_2065[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_14 (.A0(comb_d6[11]), .B0(comb6[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[12]), .B1(comb6[12]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16946), .COUT(n16947), .S0(comb7_71__N_2065[11]), 
          .S1(comb7_71__N_2065[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_12 (.A0(comb_d6[9]), .B0(comb6[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[10]), .B1(comb6[10]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16945), .COUT(n16946), .S0(comb7_71__N_2065[9]), 
          .S1(comb7_71__N_2065[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_10 (.A0(comb_d6[7]), .B0(comb6[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[8]), .B1(comb6[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16944), .COUT(n16945), .S0(comb7_71__N_2065[7]), 
          .S1(comb7_71__N_2065[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_8 (.A0(comb_d6[5]), .B0(comb6[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[6]), .B1(comb6[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16943), .COUT(n16944), .S0(comb7_71__N_2065[5]), 
          .S1(comb7_71__N_2065[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_6 (.A0(comb_d6[3]), .B0(comb6[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[4]), .B1(comb6[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16942), .COUT(n16943), .S0(comb7_71__N_2065[3]), 
          .S1(comb7_71__N_2065[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_4 (.A0(comb_d6[1]), .B0(comb6[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[2]), .B1(comb6[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16941), .COUT(n16942), .S0(comb7_71__N_2065[1]), 
          .S1(comb7_71__N_2065[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3549_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3549_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[0]), .B1(comb6[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16941), .S1(comb7_71__N_2065[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3549_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3549_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3549_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3549_add_4_2.INJECT1_1 = "NO";
    CCU2C add_5423_15 (.A0(amdemod_out_d_11__N_2409[12]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16940), .S0(n34_adj_6542));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5423_15.INIT0 = 16'haaa0;
    defparam add_5423_15.INIT1 = 16'h0000;
    defparam add_5423_15.INJECT1_0 = "NO";
    defparam add_5423_15.INJECT1_1 = "NO";
    CCU2C add_5423_13 (.A0(square_sum[25]), .B0(n19824), .C0(amdemod_out_d_11__N_2409[10]), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(amdemod_out_d_11__N_2409[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16939), .COUT(n16940));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5423_13.INIT0 = 16'h1e1e;
    defparam add_5423_13.INIT1 = 16'h666a;
    defparam add_5423_13.INJECT1_0 = "NO";
    defparam add_5423_13.INJECT1_1 = "NO";
    CCU2C add_5423_11 (.A0(n19816), .B0(amdemod_out_d_11__N_2409[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_out_d_11__N_2363), .B1(amdemod_out_d_11__N_2409[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16938), .COUT(n16939));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5423_11.INIT0 = 16'h9995;
    defparam add_5423_11.INIT1 = 16'h9995;
    defparam add_5423_11.INJECT1_0 = "NO";
    defparam add_5423_11.INJECT1_1 = "NO";
    CCU2C add_5423_9 (.A0(n19814), .B0(amdemod_out_d_11__N_2409[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19815), .B1(amdemod_out_d_11__N_2409[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16937), .COUT(n16938));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5423_9.INIT0 = 16'h9995;
    defparam add_5423_9.INIT1 = 16'h9995;
    defparam add_5423_9.INJECT1_0 = "NO";
    defparam add_5423_9.INJECT1_1 = "NO";
    CCU2C add_5423_7 (.A0(n19812), .B0(amdemod_out_d_11__N_2409[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19813), .B1(amdemod_out_d_11__N_2409[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16936), .COUT(n16937));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5423_7.INIT0 = 16'h9995;
    defparam add_5423_7.INIT1 = 16'h9995;
    defparam add_5423_7.INJECT1_0 = "NO";
    defparam add_5423_7.INJECT1_1 = "NO";
    CCU2C add_5423_5 (.A0(n19810), .B0(amdemod_out_d_11__N_2409[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19811), .B1(amdemod_out_d_11__N_2409[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16935), .COUT(n16936));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5423_5.INIT0 = 16'h9995;
    defparam add_5423_5.INIT1 = 16'h9995;
    defparam add_5423_5.INJECT1_0 = "NO";
    defparam add_5423_5.INJECT1_1 = "NO";
    CCU2C add_5423_3 (.A0(n19808), .B0(amdemod_out_d_11__N_2409[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19809), .B1(amdemod_out_d_11__N_2409[1]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16934), .COUT(n16935));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5423_3.INIT0 = 16'h9995;
    defparam add_5423_3.INIT1 = 16'h9995;
    defparam add_5423_3.INJECT1_0 = "NO";
    defparam add_5423_3.INJECT1_1 = "NO";
    CCU2C add_5423_1 (.A0(square_sum[0]), .B0(GND_net), .C0(GND_net), 
          .D0(square_sum[0]), .A1(square_sum[1]), .B1(amdemod_out_d_11__N_2410[14]), 
          .C1(n19809), .D1(amdemod_out_d_11__N_2409[14]), .COUT(n16934));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5423_1.INIT0 = 16'h000A;
    defparam add_5423_1.INIT1 = 16'h656a;
    defparam add_5423_1.INJECT1_0 = "NO";
    defparam add_5423_1.INJECT1_1 = "NO";
    CCU2C _add_1_3681_add_4_16 (.A0(amdemod_out_d_11__N_2389[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2389[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16932), .S1(n36_adj_5664));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3681_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_3681_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3681_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3681_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3681_add_4_14 (.A0(amdemod_out_d_11__N_2389[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2389[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16931), .COUT(n16932), 
          .S0(n45_adj_5665), .S1(n42));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3681_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_3681_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_3681_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3681_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3681_add_4_12 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2389[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2389[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16930), .COUT(n16931), 
          .S0(n51), .S1(n48));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3681_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3681_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_3681_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3681_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3681_add_4_10 (.A0(amdemod_out_d_11__N_2389[5]), .B0(square_sum[25]), 
          .C0(n30_adj_6282), .D0(n13890), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2389[6]), .D1(VCC_net), .CIN(n16929), 
          .COUT(n16930), .S0(n57_adj_5667), .S1(n54_adj_5666));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3681_add_4_10.INIT0 = 16'h596a;
    defparam _add_1_3681_add_4_10.INIT1 = 16'he1e1;
    defparam _add_1_3681_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3681_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3681_add_4_8 (.A0(n19815), .B0(amdemod_out_d_11__N_2389[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2389[4]), 
          .B1(amdemod_out_d_11__N_2370[11]), .C1(amdemod_out_d_11__N_2363), 
          .D1(amdemod_out_d_11__N_2369[11]), .CIN(n16928), .COUT(n16929), 
          .S0(n63_adj_5669), .S1(n60_adj_5668));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3681_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3681_add_4_8.INIT1 = 16'h656a;
    defparam _add_1_3681_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3681_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3681_add_4_6 (.A0(n19813), .B0(amdemod_out_d_11__N_2389[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2389[2]), 
          .B1(amdemod_out_d_11__N_2380[14]), .C1(n19815), .D1(amdemod_out_d_11__N_2379[14]), 
          .CIN(n16927), .COUT(n16928), .S0(n69_adj_5671), .S1(n66_adj_5670));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3681_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3681_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_3681_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3681_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3681_add_4_4 (.A0(n19812), .B0(square_sum[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_out_d_11__N_2389[0]), .B1(amdemod_out_d_11__N_2390[14]), 
          .C1(n19813), .D1(amdemod_out_d_11__N_2389[14]), .CIN(n16926), 
          .COUT(n16927), .S0(n75_adj_5673), .S1(n72_adj_5672));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3681_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3681_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_3681_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3681_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3681_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16926), .S1(n78_adj_5674));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3681_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3681_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3681_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3681_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_38 (.A0(comb_d7_adj_6566[71]), .B0(comb7_adj_6565[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16925), .S0(n78_adj_5675));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3684_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_36 (.A0(comb_d7_adj_6566[69]), .B0(comb7_adj_6565[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[70]), .B1(comb7_adj_6565[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16924), .COUT(n16925), .S0(n84_adj_5677), 
          .S1(n81_adj_5676));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_34 (.A0(comb_d7_adj_6566[67]), .B0(comb7_adj_6565[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[68]), .B1(comb7_adj_6565[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16923), .COUT(n16924), .S0(n90_adj_5679), 
          .S1(n87_adj_5678));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_32 (.A0(comb_d7_adj_6566[65]), .B0(comb7_adj_6565[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[66]), .B1(comb7_adj_6565[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16922), .COUT(n16923), .S0(n96_adj_5681), 
          .S1(n93_adj_5680));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_30 (.A0(comb_d7_adj_6566[63]), .B0(comb7_adj_6565[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[64]), .B1(comb7_adj_6565[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16921), .COUT(n16922), .S0(n102_adj_5683), 
          .S1(n99_adj_5682));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_28 (.A0(comb_d7_adj_6566[61]), .B0(comb7_adj_6565[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[62]), .B1(comb7_adj_6565[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16920), .COUT(n16921), .S0(n108_adj_5685), 
          .S1(n105_adj_5684));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_26 (.A0(comb_d7_adj_6566[59]), .B0(comb7_adj_6565[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[60]), .B1(comb7_adj_6565[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16919), .COUT(n16920), .S0(n114_adj_5687), 
          .S1(n111_adj_5686));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_24 (.A0(comb_d7_adj_6566[57]), .B0(comb7_adj_6565[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[58]), .B1(comb7_adj_6565[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16918), .COUT(n16919), .S0(n120_adj_5689), 
          .S1(n117_adj_5688));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_22 (.A0(comb_d7_adj_6566[55]), .B0(comb7_adj_6565[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[56]), .B1(comb7_adj_6565[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16917), .COUT(n16918), .S0(n126_adj_5691), 
          .S1(n123_adj_5690));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_20 (.A0(comb_d7_adj_6566[53]), .B0(comb7_adj_6565[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[54]), .B1(comb7_adj_6565[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16916), .COUT(n16917), .S0(n132_adj_5693), 
          .S1(n129_adj_5692));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_18 (.A0(comb_d7_adj_6566[51]), .B0(comb7_adj_6565[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[52]), .B1(comb7_adj_6565[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16915), .COUT(n16916), .S0(n138_adj_5695), 
          .S1(n135_adj_5694));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_16 (.A0(comb_d7_adj_6566[49]), .B0(comb7_adj_6565[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[50]), .B1(comb7_adj_6565[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16914), .COUT(n16915), .S0(n144_adj_5697), 
          .S1(n141_adj_5696));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_14 (.A0(comb_d7_adj_6566[47]), .B0(comb7_adj_6565[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[48]), .B1(comb7_adj_6565[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16913), .COUT(n16914), .S0(n150_adj_5699), 
          .S1(n147_adj_5698));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_12 (.A0(comb_d7_adj_6566[45]), .B0(comb7_adj_6565[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[46]), .B1(comb7_adj_6565[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16912), .COUT(n16913), .S0(n156_adj_5701), 
          .S1(n153_adj_5700));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_10 (.A0(comb_d7_adj_6566[43]), .B0(comb7_adj_6565[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[44]), .B1(comb7_adj_6565[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16911), .COUT(n16912), .S0(n162_adj_5703), 
          .S1(n159_adj_5702));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_8 (.A0(comb_d7_adj_6566[41]), .B0(comb7_adj_6565[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[42]), .B1(comb7_adj_6565[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16910), .COUT(n16911), .S0(n168_adj_5705), 
          .S1(n165_adj_5704));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_6 (.A0(comb_d7_adj_6566[39]), .B0(comb7_adj_6565[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[40]), .B1(comb7_adj_6565[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16909), .COUT(n16910), .S0(n174_adj_5707), 
          .S1(n171_adj_5706));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_4 (.A0(comb_d7_adj_6566[37]), .B0(comb7_adj_6565[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6566[38]), .B1(comb7_adj_6565[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16908), .COUT(n16909), .S0(n180_adj_5709), 
          .S1(n177_adj_5708));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3684_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3684_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7_adj_6566[36]), .B1(comb7_adj_6565[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16908), .S1(n183_adj_5710));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3684_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3684_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3684_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3684_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3687_add_4_16 (.A0(amdemod_out_d_11__N_2380[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2380[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16906), .S1(n36_adj_5711));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3687_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_3687_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3687_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3687_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3687_add_4_14 (.A0(amdemod_out_d_11__N_2380[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2380[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16905), .COUT(n16906), 
          .S0(n45_adj_5713), .S1(n42_adj_5712));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3687_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_3687_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_3687_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3687_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3687_add_4_12 (.A0(amdemod_out_d_11__N_2380[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2380[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16904), .COUT(n16905), 
          .S0(n51_adj_5715), .S1(n48_adj_5714));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3687_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_3687_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_3687_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3687_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3687_add_4_10 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2380[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2380[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16903), .COUT(n16904), 
          .S0(n57_adj_5717), .S1(n54_adj_5716));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3687_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3687_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_3687_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3687_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3687_add_4_8 (.A0(amdemod_out_d_11__N_2380[3]), .B0(square_sum[25]), 
          .C0(n30_adj_6282), .D0(n13890), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2380[4]), .D1(VCC_net), .CIN(n16902), 
          .COUT(n16903), .S0(n63_adj_5719), .S1(n60_adj_5718));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3687_add_4_8.INIT0 = 16'h596a;
    defparam _add_1_3687_add_4_8.INIT1 = 16'he1e1;
    defparam _add_1_3687_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3687_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3687_add_4_6 (.A0(n19815), .B0(amdemod_out_d_11__N_2380[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2380[2]), 
          .B1(amdemod_out_d_11__N_2370[11]), .C1(amdemod_out_d_11__N_2363), 
          .D1(amdemod_out_d_11__N_2369[11]), .CIN(n16901), .COUT(n16902), 
          .S0(n69_adj_5721), .S1(n66_adj_5720));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3687_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3687_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_3687_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3687_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3687_add_4_4 (.A0(n19814), .B0(square_sum[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_out_d_11__N_2380[0]), .B1(amdemod_out_d_11__N_2380[14]), 
          .C1(n19815), .D1(amdemod_out_d_11__N_2379[14]), .CIN(n16900), 
          .COUT(n16901), .S0(n75_adj_5723), .S1(n72_adj_5722));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3687_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3687_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_3687_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3687_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3687_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16900), .S1(n78_adj_5724));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3687_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3687_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3687_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3687_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_38 (.A0(comb_d6_adj_6564[71]), .B0(comb6_adj_6563[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16899), .S0(n78_adj_5725));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3690_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_36 (.A0(comb_d6_adj_6564[69]), .B0(comb6_adj_6563[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[70]), .B1(comb6_adj_6563[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16898), .COUT(n16899), .S0(n84_adj_5727), 
          .S1(n81_adj_5726));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_34 (.A0(comb_d6_adj_6564[67]), .B0(comb6_adj_6563[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[68]), .B1(comb6_adj_6563[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16897), .COUT(n16898), .S0(n90_adj_5729), 
          .S1(n87_adj_5728));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_32 (.A0(comb_d6_adj_6564[65]), .B0(comb6_adj_6563[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[66]), .B1(comb6_adj_6563[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16896), .COUT(n16897), .S0(n96_adj_5731), 
          .S1(n93_adj_5730));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_30 (.A0(comb_d6_adj_6564[63]), .B0(comb6_adj_6563[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[64]), .B1(comb6_adj_6563[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16895), .COUT(n16896), .S0(n102_adj_5733), 
          .S1(n99_adj_5732));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_28 (.A0(comb_d6_adj_6564[61]), .B0(comb6_adj_6563[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[62]), .B1(comb6_adj_6563[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16894), .COUT(n16895), .S0(n108_adj_5735), 
          .S1(n105_adj_5734));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_26 (.A0(comb_d6_adj_6564[59]), .B0(comb6_adj_6563[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[60]), .B1(comb6_adj_6563[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16893), .COUT(n16894), .S0(n114_adj_5737), 
          .S1(n111_adj_5736));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_24 (.A0(comb_d6_adj_6564[57]), .B0(comb6_adj_6563[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[58]), .B1(comb6_adj_6563[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16892), .COUT(n16893), .S0(n120_adj_5739), 
          .S1(n117_adj_5738));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_22 (.A0(comb_d6_adj_6564[55]), .B0(comb6_adj_6563[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[56]), .B1(comb6_adj_6563[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16891), .COUT(n16892), .S0(n126_adj_5741), 
          .S1(n123_adj_5740));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_20 (.A0(comb_d6_adj_6564[53]), .B0(comb6_adj_6563[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[54]), .B1(comb6_adj_6563[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16890), .COUT(n16891), .S0(n132_adj_5743), 
          .S1(n129_adj_5742));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_18 (.A0(comb_d6_adj_6564[51]), .B0(comb6_adj_6563[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[52]), .B1(comb6_adj_6563[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16889), .COUT(n16890), .S0(n138_adj_5745), 
          .S1(n135_adj_5744));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_16 (.A0(comb_d6_adj_6564[49]), .B0(comb6_adj_6563[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[50]), .B1(comb6_adj_6563[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16888), .COUT(n16889), .S0(n144_adj_5747), 
          .S1(n141_adj_5746));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_14 (.A0(comb_d6_adj_6564[47]), .B0(comb6_adj_6563[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[48]), .B1(comb6_adj_6563[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16887), .COUT(n16888), .S0(n150_adj_5749), 
          .S1(n147_adj_5748));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_12 (.A0(comb_d6_adj_6564[45]), .B0(comb6_adj_6563[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[46]), .B1(comb6_adj_6563[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16886), .COUT(n16887), .S0(n156_adj_5751), 
          .S1(n153_adj_5750));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_10 (.A0(comb_d6_adj_6564[43]), .B0(comb6_adj_6563[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[44]), .B1(comb6_adj_6563[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16885), .COUT(n16886), .S0(n162_adj_5753), 
          .S1(n159_adj_5752));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_8 (.A0(comb_d6_adj_6564[41]), .B0(comb6_adj_6563[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[42]), .B1(comb6_adj_6563[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16884), .COUT(n16885), .S0(n168_adj_5755), 
          .S1(n165_adj_5754));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_6 (.A0(comb_d6_adj_6564[39]), .B0(comb6_adj_6563[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[40]), .B1(comb6_adj_6563[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16883), .COUT(n16884), .S0(n174_adj_5757), 
          .S1(n171_adj_5756));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_4 (.A0(comb_d6_adj_6564[37]), .B0(comb6_adj_6563[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6564[38]), .B1(comb6_adj_6563[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16882), .COUT(n16883), .S0(n180_adj_5759), 
          .S1(n177_adj_5758));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3690_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3690_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6_adj_6564[36]), .B1(comb6_adj_6563[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16882), .S1(n183_adj_5760));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam _add_1_3690_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3690_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3690_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3690_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_38 (.A0(integrator_d_tmp_adj_6557[71]), .B0(integrator_tmp_adj_6556[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16881), .S0(n78_adj_5761));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3693_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_36 (.A0(integrator_d_tmp_adj_6557[69]), .B0(integrator_tmp_adj_6556[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[70]), 
          .B1(integrator_tmp_adj_6556[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16880), .COUT(n16881), .S0(n84_adj_5763), .S1(n81_adj_5762));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_34 (.A0(integrator_d_tmp_adj_6557[67]), .B0(integrator_tmp_adj_6556[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[68]), 
          .B1(integrator_tmp_adj_6556[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16879), .COUT(n16880), .S0(n90_adj_5765), .S1(n87_adj_5764));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_32 (.A0(integrator_d_tmp_adj_6557[65]), .B0(integrator_tmp_adj_6556[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[66]), 
          .B1(integrator_tmp_adj_6556[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16878), .COUT(n16879), .S0(n96_adj_5767), .S1(n93_adj_5766));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_30 (.A0(integrator_d_tmp_adj_6557[63]), .B0(integrator_tmp_adj_6556[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[64]), 
          .B1(integrator_tmp_adj_6556[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16877), .COUT(n16878), .S0(n102_adj_5769), .S1(n99_adj_5768));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_28 (.A0(integrator_d_tmp_adj_6557[61]), .B0(integrator_tmp_adj_6556[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[62]), 
          .B1(integrator_tmp_adj_6556[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16876), .COUT(n16877), .S0(n108_adj_5771), .S1(n105_adj_5770));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_26 (.A0(integrator_d_tmp_adj_6557[59]), .B0(integrator_tmp_adj_6556[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[60]), 
          .B1(integrator_tmp_adj_6556[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16875), .COUT(n16876), .S0(n114_adj_5773), .S1(n111_adj_5772));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_24 (.A0(integrator_d_tmp_adj_6557[57]), .B0(integrator_tmp_adj_6556[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[58]), 
          .B1(integrator_tmp_adj_6556[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16874), .COUT(n16875), .S0(n120_adj_5775), .S1(n117_adj_5774));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_22 (.A0(integrator_d_tmp_adj_6557[55]), .B0(integrator_tmp_adj_6556[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[56]), 
          .B1(integrator_tmp_adj_6556[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16873), .COUT(n16874), .S0(n126_adj_5777), .S1(n123_adj_5776));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_20 (.A0(integrator_d_tmp_adj_6557[53]), .B0(integrator_tmp_adj_6556[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[54]), 
          .B1(integrator_tmp_adj_6556[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16872), .COUT(n16873), .S0(n132_adj_5779), .S1(n129_adj_5778));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_18 (.A0(integrator_d_tmp_adj_6557[51]), .B0(integrator_tmp_adj_6556[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[52]), 
          .B1(integrator_tmp_adj_6556[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16871), .COUT(n16872), .S0(n138_adj_5781), .S1(n135_adj_5780));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_16 (.A0(integrator_d_tmp_adj_6557[49]), .B0(integrator_tmp_adj_6556[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[50]), 
          .B1(integrator_tmp_adj_6556[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16870), .COUT(n16871), .S0(n144_adj_5783), .S1(n141_adj_5782));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_14 (.A0(integrator_d_tmp_adj_6557[47]), .B0(integrator_tmp_adj_6556[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[48]), 
          .B1(integrator_tmp_adj_6556[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16869), .COUT(n16870), .S0(n150_adj_5785), .S1(n147_adj_5784));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_12 (.A0(integrator_d_tmp_adj_6557[45]), .B0(integrator_tmp_adj_6556[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[46]), 
          .B1(integrator_tmp_adj_6556[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16868), .COUT(n16869), .S0(n156_adj_5787), .S1(n153_adj_5786));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_10 (.A0(integrator_d_tmp_adj_6557[43]), .B0(integrator_tmp_adj_6556[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[44]), 
          .B1(integrator_tmp_adj_6556[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16867), .COUT(n16868), .S0(n162_adj_5789), .S1(n159_adj_5788));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_8 (.A0(integrator_d_tmp_adj_6557[41]), .B0(integrator_tmp_adj_6556[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[42]), 
          .B1(integrator_tmp_adj_6556[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16866), .COUT(n16867), .S0(n168_adj_5791), .S1(n165_adj_5790));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_6 (.A0(integrator_d_tmp_adj_6557[39]), .B0(integrator_tmp_adj_6556[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[40]), 
          .B1(integrator_tmp_adj_6556[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16865), .COUT(n16866), .S0(n174_adj_5793), .S1(n171_adj_5792));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_4 (.A0(integrator_d_tmp_adj_6557[37]), .B0(integrator_tmp_adj_6556[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[38]), 
          .B1(integrator_tmp_adj_6556[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16864), .COUT(n16865), .S0(n180_adj_5795), .S1(n177_adj_5794));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3693_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3693_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator_d_tmp_adj_6557[36]), .B1(integrator_tmp_adj_6556[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16864), .S1(n183_adj_5796));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3693_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3693_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_3693_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3693_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3696_add_4_16 (.A0(amdemod_out_d_11__N_2379[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2379[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16862), .S1(n36_adj_5797));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3696_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_3696_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3696_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3696_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3696_add_4_14 (.A0(amdemod_out_d_11__N_2379[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2379[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16861), .COUT(n16862), 
          .S0(n45_adj_5799), .S1(n42_adj_5798));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3696_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_3696_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_3696_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3696_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3696_add_4_12 (.A0(amdemod_out_d_11__N_2379[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2379[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16860), .COUT(n16861), 
          .S0(n51_adj_5801), .S1(n48_adj_5800));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3696_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_3696_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_3696_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3696_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3696_add_4_10 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2379[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2379[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16859), .COUT(n16860), 
          .S0(n57_adj_5803), .S1(n54_adj_5802));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3696_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_3696_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_3696_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3696_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3696_add_4_8 (.A0(amdemod_out_d_11__N_2379[3]), .B0(square_sum[25]), 
          .C0(n30_adj_6282), .D0(n13890), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2379[4]), .D1(VCC_net), .CIN(n16858), 
          .COUT(n16859), .S0(n63_adj_5805), .S1(n60_adj_5804));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3696_add_4_8.INIT0 = 16'h596a;
    defparam _add_1_3696_add_4_8.INIT1 = 16'he1e1;
    defparam _add_1_3696_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3696_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3696_add_4_6 (.A0(n19815), .B0(amdemod_out_d_11__N_2379[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2379[2]), 
          .B1(amdemod_out_d_11__N_2370[11]), .C1(amdemod_out_d_11__N_2363), 
          .D1(amdemod_out_d_11__N_2369[11]), .CIN(n16857), .COUT(n16858), 
          .S0(n69_adj_5807), .S1(n66_adj_5806));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3696_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3696_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_3696_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3696_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3696_add_4_4 (.A0(n19814), .B0(square_sum[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_out_d_11__N_2379[0]), .B1(amdemod_out_d_11__N_2380[14]), 
          .C1(n19815), .D1(amdemod_out_d_11__N_2379[14]), .CIN(n16856), 
          .COUT(n16857), .S0(n75_adj_5809), .S1(n72_adj_5808));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3696_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3696_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_3696_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3696_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3696_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16856), .S1(n78_adj_5810));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3696_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3696_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3696_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3696_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3699_add_4_16 (.A0(amdemod_out_d_11__N_2370[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2370[11]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16854), .S1(n36_adj_5811));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3699_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_3699_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3699_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3699_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3699_add_4_14 (.A0(amdemod_out_d_11__N_2370[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2370[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16853), .COUT(n16854), 
          .S0(n45_adj_5813), .S1(n42_adj_5812));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3699_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_3699_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_3699_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3699_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3699_add_4_12 (.A0(amdemod_out_d_11__N_2370[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2370[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16852), .COUT(n16853), 
          .S0(n51_adj_5815), .S1(n48_adj_5814));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3699_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_3699_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_3699_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3699_add_4_12.INJECT1_1 = "NO";
    LUT4 mux_1437_i1_3_lut (.A(phase_increment_1__63__N_16[36]), .B(phase_increment_1__63__N_18[36]), 
         .C(rx_byte[0]), .Z(n2682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1437_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1402_i1_3_lut (.A(phase_increment_1__63__N_16[37]), .B(phase_increment_1__63__N_18[37]), 
         .C(rx_byte[0]), .Z(n2635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1402_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1507_i1_3_lut (.A(phase_increment_1__63__N_16[34]), .B(phase_increment_1__63__N_18[34]), 
         .C(rx_byte[0]), .Z(n2776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1507_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1472_i1_3_lut (.A(phase_increment_1__63__N_16[35]), .B(phase_increment_1__63__N_18[35]), 
         .C(rx_byte[0]), .Z(n2729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1472_i1_3_lut.init = 16'hcaca;
    LUT4 phase_increment_1__63__N_21_32__bdd_2_lut_8619 (.A(led_0_6), .B(phase_increment_1__63__N_17[32]), 
         .Z(n19662)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_32__bdd_2_lut_8619.init = 16'heeee;
    PFUMX mux_2618_i1 (.BLUT(n4248), .ALUT(n4264), .C0(n19134), .Z(n4267));
    LUT4 phase_increment_1__63__N_21_45__bdd_2_lut_8841 (.A(phase_increment_1__63__N_21[45]), 
         .B(rx_byte[0]), .Z(n19586)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_45__bdd_2_lut_8841.init = 16'heeee;
    LUT4 mux_2522_i1_3_lut (.A(phase_increment_1__63__N_16[5]), .B(phase_increment_1__63__N_18[5]), 
         .C(rx_byte[0]), .Z(n4139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2522_i1_3_lut.init = 16'hcaca;
    LUT4 phase_increment_1__63__N_21_59__bdd_2_lut_8469 (.A(phase_increment_1__63__N_17[59]), 
         .B(led_0_6), .Z(n19447)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_59__bdd_2_lut_8469.init = 16'heeee;
    LUT4 mux_784_i1_3_lut (.A(phase_increment_1__63__N_19[55]), .B(phase_increment_1__63__N_20[55]), 
         .C(rx_byte[0]), .Z(n1804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_784_i1_3_lut.init = 16'hcaca;
    PFUMX mux_2126_i1 (.BLUT(n3590), .ALUT(n3600), .C0(led_0_6), .Z(n3606));
    PFUMX mux_2583_i1 (.BLUT(n4211), .ALUT(n4217), .C0(n19300), .Z(n4220));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 mux_1974_i1_3_lut (.A(phase_increment_1__63__N_19[21]), .B(phase_increment_1__63__N_20[21]), 
         .C(rx_byte[0]), .Z(n3402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1974_i1_3_lut.init = 16'hcaca;
    LUT4 mux_2534_i1_3_lut (.A(phase_increment_1__63__N_19[5]), .B(phase_increment_1__63__N_20[5]), 
         .C(rx_byte[0]), .Z(n4154)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2534_i1_3_lut.init = 16'hcaca;
    PFUMX mux_1463_i1 (.BLUT(n2707), .ALUT(n2713), .C0(n19296), .Z(n2716));
    LUT4 n2870_bdd_3_lut_8622 (.A(n2870), .B(rx_byte[2]), .C(rx_byte[3]), 
         .Z(n19665)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n2870_bdd_3_lut_8622.init = 16'hacac;
    LUT4 n2870_bdd_3_lut (.A(phase_increment_1__63__N_19[32]), .B(phase_increment_1__63__N_20[32]), 
         .C(rx_byte[0]), .Z(n19666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n2870_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_1554_i1_3_lut (.A(phase_increment_1__63__N_19[33]), .B(phase_increment_1__63__N_20[33]), 
         .C(rx_byte[0]), .Z(n2838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1554_i1_3_lut.init = 16'hcaca;
    PFUMX mux_1428_i1 (.BLUT(n2660), .ALUT(n2666), .C0(n19295), .Z(n2669));
    LUT4 mux_1577_i1_3_lut (.A(phase_increment_1__63__N_16[32]), .B(phase_increment_1__63__N_18[32]), 
         .C(rx_byte[0]), .Z(n2870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1577_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1542_i1_3_lut (.A(phase_increment_1__63__N_16[33]), .B(phase_increment_1__63__N_18[33]), 
         .C(rx_byte[0]), .Z(n2823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1542_i1_3_lut.init = 16'hcaca;
    LUT4 mux_749_i1_3_lut (.A(phase_increment_1__63__N_19[56]), .B(phase_increment_1__63__N_20[56]), 
         .C(rx_byte[0]), .Z(n1757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_749_i1_3_lut.init = 16'hcaca;
    LUT4 phase_increment_1__63__N_21_26__bdd_2_lut_2_lut (.A(rx_byte[0]), 
         .B(phase_increment_1__63__N_21[26]), .Z(n19411)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam phase_increment_1__63__N_21_26__bdd_2_lut_2_lut.init = 16'h4444;
    PFUMX mux_1319_i1 (.BLUT(n2514), .ALUT(n2499), .C0(rx_byte[2]), .Z(n2522));
    LUT4 phase_increment_1__63__N_21_36__bdd_2_lut_8924 (.A(phase_increment_1__63__N_21[36]), 
         .B(rx_byte[0]), .Z(n19677)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_36__bdd_2_lut_8924.init = 16'heeee;
    PFUMX mux_1284_i1 (.BLUT(n2467), .ALUT(n2452), .C0(rx_byte[2]), .Z(n2475));
    LUT4 mux_2207_i1_3_lut (.A(phase_increment_1__63__N_16[14]), .B(phase_increment_1__63__N_18[14]), 
         .C(rx_byte[0]), .Z(n3716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2207_i1_3_lut.init = 16'hcaca;
    LUT4 i4889_2_lut_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[63]), 
         .Z(n1433)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i4889_2_lut_2_lut.init = 16'h4444;
    LUT4 i4876_2_lut_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[62]), 
         .Z(n1480)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i4876_2_lut_2_lut.init = 16'h4444;
    LUT4 mux_2569_i1_3_lut (.A(phase_increment_1__63__N_19[4]), .B(phase_increment_1__63__N_20[4]), 
         .C(rx_byte[0]), .Z(n4201)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2569_i1_3_lut.init = 16'hcaca;
    LUT4 i4961_2_lut (.A(phase_increment_1__63__N_17[29]), .B(led_0_6), 
         .Z(n3016)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4961_2_lut.init = 16'heeee;
    LUT4 mux_1787_i1_3_lut (.A(phase_increment_1__63__N_16[26]), .B(phase_increment_1__63__N_18[26]), 
         .C(rx_byte[0]), .Z(n3152)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1787_i1_3_lut.init = 16'hcaca;
    LUT4 phase_increment_1__63__N_21_37__bdd_2_lut_8635 (.A(phase_increment_1__63__N_17[37]), 
         .B(led_0_6), .Z(n19679)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_37__bdd_2_lut_8635.init = 16'heeee;
    LUT4 mux_1752_i1_3_lut (.A(phase_increment_1__63__N_16[27]), .B(phase_increment_1__63__N_18[27]), 
         .C(rx_byte[0]), .Z(n3105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1752_i1_3_lut.init = 16'hcaca;
    LUT4 i4866_2_lut_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[61]), 
         .Z(n1527)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i4866_2_lut_2_lut.init = 16'h4444;
    LUT4 i4115_2_lut_4_lut_rep_308 (.A(n26_adj_5299), .B(n19825), .C(n45), 
         .D(rx_data_valid), .Z(clk_80mhz_enable_223)) /* synthesis lut_function=(A (B (D))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(265[5] 289[6])
    defparam i4115_2_lut_4_lut_rep_308.init = 16'hc800;
    LUT4 mux_1647_i1_3_lut (.A(phase_increment_1__63__N_16[30]), .B(phase_increment_1__63__N_18[30]), 
         .C(rx_byte[0]), .Z(n2964)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1647_i1_3_lut.init = 16'hcaca;
    PFUMX mux_1498_i1 (.BLUT(n2754), .ALUT(n2760), .C0(n19294), .Z(n2763));
    LUT4 mux_1857_i1_3_lut (.A(phase_increment_1__63__N_16[24]), .B(phase_increment_1__63__N_18[24]), 
         .C(rx_byte[0]), .Z(n3246)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1857_i1_3_lut.init = 16'hcaca;
    LUT4 i47_4_lut_then_3_lut (.A(led_0_6), .B(rx_byte[2]), .C(rx_byte[3]), 
         .Z(n19857)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i47_4_lut_then_3_lut.init = 16'h0101;
    LUT4 mux_2612_i1_4_lut (.A(rx_byte[2]), .B(phase_increment_1__63__N_18[3]), 
         .C(rx_byte[3]), .D(rx_byte[0]), .Z(n4258)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2612_i1_4_lut.init = 16'hca0a;
    LUT4 mux_2347_i1_3_lut (.A(phase_increment_1__63__N_16[10]), .B(phase_increment_1__63__N_18[10]), 
         .C(rx_byte[0]), .Z(n3904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2347_i1_3_lut.init = 16'hcaca;
    LUT4 i47_4_lut_else_3_lut (.A(led_0_6), .B(rx_byte[2]), .C(rx_byte[3]), 
         .D(rx_byte[0]), .Z(n19856)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))) */ ;
    defparam i47_4_lut_else_3_lut.init = 16'h808a;
    LUT4 phase_increment_1__63__N_21_14__bdd_2_lut_8692 (.A(phase_increment_1__63__N_21[14]), 
         .B(rx_byte[0]), .Z(n19683)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_14__bdd_2_lut_8692.init = 16'heeee;
    LUT4 mux_1822_i1_3_lut (.A(phase_increment_1__63__N_16[25]), .B(phase_increment_1__63__N_18[25]), 
         .C(rx_byte[0]), .Z(n3199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1822_i1_3_lut.init = 16'hcaca;
    LUT4 i4904_2_lut_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[56]), 
         .Z(n1762)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i4904_2_lut_2_lut.init = 16'h4444;
    LUT4 i8017_3_lut (.A(n4295), .B(n4305), .C(led_0_6), .Z(n4311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i8017_3_lut.init = 16'hcaca;
    PFUMX i8502 (.BLUT(n19492), .ALUT(n19491), .C0(rx_byte[2]), .Z(n19493));
    PFUMX mux_2548_i1 (.BLUT(n4164), .ALUT(n4170), .C0(n19302), .Z(n4173));
    LUT4 i4908_2_lut_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[52]), 
         .Z(n1950)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i4908_2_lut_2_lut.init = 16'h4444;
    LUT4 i8154_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19702), 
         .D(n2838), .Z(n2854)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8154_3_lut_4_lut.init = 16'hf780;
    LUT4 i8019_3_lut (.A(n4342), .B(n18600), .C(led_0_6), .Z(n4358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i8019_3_lut.init = 16'hcaca;
    PFUMX mux_1568_i1 (.BLUT(n2848), .ALUT(n2854), .C0(n19299), .Z(n2857));
    LUT4 i8208_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19603), 
         .D(n2415), .Z(n2431)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8208_3_lut_4_lut.init = 16'hf780;
    LUT4 i4994_2_lut (.A(phase_increment_1__63__N_17[15]), .B(led_0_6), 
         .Z(n3674)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4994_2_lut.init = 16'heeee;
    L6MUX21 i8683 (.D0(n19736), .D1(n19733), .SD(n19822), .Z(n19737));
    LUT4 i4927_2_lut_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[44]), 
         .Z(n2326)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i4927_2_lut_2_lut.init = 16'h4444;
    LUT4 n3716_bdd_3_lut_8641 (.A(n3716), .B(rx_byte[2]), .C(rx_byte[3]), 
         .Z(n19685)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n3716_bdd_3_lut_8641.init = 16'hacac;
    LUT4 i4934_2_lut_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[41]), 
         .Z(n2467)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i4934_2_lut_2_lut.init = 16'h4444;
    LUT4 mux_644_i1_3_lut (.A(phase_increment_1__63__N_19[59]), .B(phase_increment_1__63__N_20[59]), 
         .C(rx_byte[0]), .Z(n1616)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_644_i1_3_lut.init = 16'hcaca;
    PFUMX i8681 (.BLUT(n19735), .ALUT(n19734), .C0(led_0_6), .Z(n19736));
    LUT4 i4903_4_lut_4_lut (.A(rx_byte[3]), .B(rx_byte[0]), .C(phase_increment_1__63__N_18[56]), 
         .D(phase_increment_1__63__N_16[56]), .Z(n1767)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(265[5] 289[6])
    defparam i4903_4_lut_4_lut.init = 16'hf7d5;
    LUT4 n3716_bdd_3_lut (.A(phase_increment_1__63__N_19[14]), .B(phase_increment_1__63__N_20[14]), 
         .C(rx_byte[0]), .Z(n19686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3716_bdd_3_lut.init = 16'hcaca;
    PFUMX mux_1984_i1 (.BLUT(n3407), .ALUT(n3392), .C0(rx_byte[2]), .Z(n3415));
    PFUMX i8431 (.BLUT(n19411), .ALUT(n19410), .C0(rx_byte[2]), .Z(n19412));
    LUT4 i4962_2_lut_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[29]), 
         .Z(n3031)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i4962_2_lut_2_lut.init = 16'h4444;
    LUT4 i4990_2_lut_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[17]), 
         .Z(n3595)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i4990_2_lut_2_lut.init = 16'h4444;
    LUT4 i8131_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19765), 
         .D(n3073), .Z(n3089)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8131_3_lut_4_lut.init = 16'hf780;
    LUT4 i5003_2_lut_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[12]), 
         .Z(n3830)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i5003_2_lut_2_lut.init = 16'h4444;
    LUT4 i8178_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19681), 
         .D(n2650), .Z(n2666)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8178_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1764_i1_3_lut (.A(phase_increment_1__63__N_19[27]), .B(phase_increment_1__63__N_20[27]), 
         .C(rx_byte[0]), .Z(n3120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1764_i1_3_lut.init = 16'hcaca;
    LUT4 i8226_3_lut_4_lut (.A(n26_adj_5299), .B(n19825), .C(n19552), 
         .D(n2227), .Z(n2243)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i8226_3_lut_4_lut.init = 16'hf780;
    PFUMX i8496 (.BLUT(n19479), .ALUT(n19478), .C0(rx_byte[2]), .Z(n19480));
    LUT4 i5000_2_lut_2_lut (.A(rx_byte[0]), .B(phase_increment_1__63__N_21[13]), 
         .Z(n3783)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i5000_2_lut_2_lut.init = 16'h4444;
    LUT4 mux_2649_i1_4_lut_4_lut (.A(rx_byte[0]), .B(rx_byte[2]), .C(led_0_6), 
         .D(phase_increment_1__63__N_21[2]), .Z(n4308)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam mux_2649_i1_4_lut_4_lut.init = 16'hd1c0;
    PFUMX mux_2511_i1 (.BLUT(n4107), .ALUT(n4117), .C0(led_0_6), .Z(n4123));
    LUT4 i1_2_lut_3_lut_3_lut (.A(rx_byte[0]), .B(rx_byte[3]), .C(led_0_6), 
         .Z(n18704)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam i1_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 i4886_4_lut (.A(phase_increment_1__63__N_16[57]), .B(rx_byte[3]), 
         .C(phase_increment_1__63__N_18[57]), .D(rx_byte[0]), .Z(n1720)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam i4886_4_lut.init = 16'hc088;
    LUT4 pwm_out_I_0_1_lut (.A(pwm_out_c), .Z(pwm_out_p_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(257[24:32])
    defparam pwm_out_I_0_1_lut.init = 16'h5555;
    PFUMX i8678 (.BLUT(n19732), .ALUT(n19731), .C0(rx_byte[2]), .Z(n19733));
    LUT4 mux_714_i1_3_lut (.A(phase_increment_1__63__N_19[57]), .B(phase_increment_1__63__N_20[57]), 
         .C(rx_byte[0]), .Z(n1710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_714_i1_3_lut.init = 16'hcaca;
    PFUMX mux_2196_i1 (.BLUT(n3684), .ALUT(n3694), .C0(led_0_6), .Z(n3700));
    MUX21 i8400 (.D0(n1820), .D1(n1817), .SD(n19822), .Z(n1823));
    MUX21 i8413 (.D0(n3888), .D1(n3885), .SD(n19822), .Z(n3891));
    PFUMX mux_1813_i1 (.BLUT(n3177), .ALUT(n3183), .C0(n19296), .Z(n3186));
    PFUMX mux_1778_i1 (.BLUT(n3130), .ALUT(n3136), .C0(n19294), .Z(n3139));
    MUX21 i8414 (.D0(n3841), .D1(n3838), .SD(n19822), .Z(n3844));
    MUX21 i8415 (.D0(n3418), .D1(n3415), .SD(n19822), .Z(n3421));
    PFUMX mux_2054_i1 (.BLUT(n3501), .ALUT(n3486), .C0(rx_byte[2]), .Z(n3509));
    LUT4 i1_3_lut_adj_241 (.A(rx_byte[3]), .B(phase_increment_1__63__N_18[1]), 
         .C(rx_byte[0]), .Z(n18600)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_241.init = 16'h8080;
    MUX21 i8416 (.D0(n3371), .D1(n3368), .SD(n19822), .Z(n3374));
    LUT4 mux_1834_i1_3_lut (.A(phase_increment_1__63__N_19[25]), .B(phase_increment_1__63__N_20[25]), 
         .C(rx_byte[0]), .Z(n3214)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1834_i1_3_lut.init = 16'hcaca;
    MUX21 i8401 (.D0(n3512), .D1(n3509), .SD(n19822), .Z(n3515));
    MUX21 i8417 (.D0(n1444), .D1(n1441), .SD(n19822), .Z(n1447));
    MUX21 i8418 (.D0(n1491), .D1(n1488), .SD(n19822), .Z(n1494));
    VLO i1 (.Z(GND_net));
    PFUMX mux_2266_i1 (.BLUT(n3778), .ALUT(n3788), .C0(led_0_6), .Z(n3794));
    MUX21 i8419 (.D0(n1538), .D1(n1535), .SD(n19822), .Z(n1541));
    PFUMX i8669 (.BLUT(n19722), .ALUT(n19721), .C0(rx_byte[2]), .Z(n19723));
    MUX21 i8420 (.D0(n1726), .D1(n1723), .SD(n19822), .Z(n1729));
    MUX21 i8421 (.D0(n3042), .D1(n3039), .SD(n19822), .Z(n3045));
    MUX21 i8402 (.D0(n4076), .D1(n4073), .SD(n19822), .Z(n4079));
    MUX21 i8403 (.D0(n1961), .D1(n1958), .SD(n19822), .Z(n1964));
    PFUMX i8666 (.BLUT(n19719), .ALUT(n19718), .C0(rx_byte[2]), .Z(n19720));
    MUX21 i8404 (.D0(n2102), .D1(n2099), .SD(n19822), .Z(n2105));
    PFUMX i8490 (.BLUT(n19473), .ALUT(n19472), .C0(rx_byte[2]), .Z(n19474));
    MUX21 i8405 (.D0(n2055), .D1(n2052), .SD(n19822), .Z(n2058));
    MUX21 i8406 (.D0(n4123), .D1(n4120), .SD(n19822), .Z(n4126));
    PFUMX mux_2124_i1 (.BLUT(n3595), .ALUT(n3580), .C0(rx_byte[2]), .Z(n3603));
    MUX21 i8399 (.D0(n1773), .D1(n1770), .SD(n19822), .Z(n1776));
    MUX21 i8407 (.D0(n2337), .D1(n2334), .SD(n19822), .Z(n2340));
    MUX21 i8408 (.D0(n3606), .D1(n3603), .SD(n19822), .Z(n3609));
    MUX21 i8409 (.D0(n2478), .D1(n2475), .SD(n19822), .Z(n2481));
    MUX21 i8410 (.D0(n2525), .D1(n2522), .SD(n19822), .Z(n2528));
    MUX21 i8411 (.D0(n3700), .D1(n3697), .SD(n19822), .Z(n3703));
    PFUMX mux_2373_i1 (.BLUT(n3929), .ALUT(n3935), .C0(n19295), .Z(n3938));
    PFUMX mux_2336_i1 (.BLUT(n3872), .ALUT(n3882), .C0(led_0_6), .Z(n3888));
    PFUMX mux_1848_i1 (.BLUT(n3224), .ALUT(n3230), .C0(n19295), .Z(n3233));
    PFUMX mux_2301_i1 (.BLUT(n3825), .ALUT(n3835), .C0(led_0_6), .Z(n3841));
    PFUMX i8663 (.BLUT(n19716), .ALUT(n19715), .C0(rx_byte[2]), .Z(n19717));
    PFUMX i8655 (.BLUT(n19701), .ALUT(n19700), .C0(rx_byte[2]), .Z(n19702));
    PFUMX mux_2194_i1 (.BLUT(n3689), .ALUT(n3674), .C0(rx_byte[2]), .Z(n3697));
    PFUMX i8767 (.BLUT(n19862), .ALUT(n19863), .C0(led_0_6), .Z(n26_adj_5299));
    LUT4 i5023_4_lut_4_lut (.A(rx_byte[3]), .B(rx_byte[0]), .C(phase_increment_1__63__N_18[6]), 
         .D(phase_increment_1__63__N_16[6]), .Z(n4117)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(265[5] 289[6])
    defparam i5023_4_lut_4_lut.init = 16'hf7d5;
    L6MUX21 i8644 (.D0(n19687), .D1(n19684), .SD(n19822), .Z(n19688));
    PFUMX i8642 (.BLUT(n19686), .ALUT(n19685), .C0(led_0_6), .Z(n19687));
    LUT4 mux_2674_i1_3_lut (.A(phase_increment_1__63__N_19[1]), .B(phase_increment_1__63__N_20[1]), 
         .C(rx_byte[0]), .Z(n4342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_2674_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3807_add_4_59 (.A0(\phase_increment[0] [57]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [58]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17659), .COUT(n17660), .S0(phase_increment_1__63__N_18[57]), 
          .S1(phase_increment_1__63__N_18[58]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_57 (.A0(\phase_increment[0] [55]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [56]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17658), .COUT(n17659), .S0(phase_increment_1__63__N_18[55]), 
          .S1(phase_increment_1__63__N_18[56]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_55 (.A0(\phase_increment[0] [53]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [54]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17657), .COUT(n17658), .S0(phase_increment_1__63__N_18[53]), 
          .S1(phase_increment_1__63__N_18[54]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_53 (.A0(\phase_increment[0] [51]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [52]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17656), .COUT(n17657), .S0(phase_increment_1__63__N_18[51]), 
          .S1(phase_increment_1__63__N_18[52]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_51 (.A0(\phase_increment[0] [49]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [50]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17655), .COUT(n17656), .S0(phase_increment_1__63__N_18[49]), 
          .S1(phase_increment_1__63__N_18[50]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_49 (.A0(\phase_increment[0] [47]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [48]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17654), .COUT(n17655), .S0(phase_increment_1__63__N_18[47]), 
          .S1(phase_increment_1__63__N_18[48]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_47 (.A0(\phase_increment[0] [45]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [46]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17653), .COUT(n17654), .S0(phase_increment_1__63__N_18[45]), 
          .S1(phase_increment_1__63__N_18[46]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_47.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_47.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_45 (.A0(\phase_increment[0] [43]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [44]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17652), .COUT(n17653), .S0(phase_increment_1__63__N_18[43]), 
          .S1(phase_increment_1__63__N_18[44]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_45.INIT1 = 16'haaa0;
    defparam _add_1_3807_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_43 (.A0(\phase_increment[0] [41]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [42]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17651), .COUT(n17652), .S0(phase_increment_1__63__N_18[41]), 
          .S1(phase_increment_1__63__N_18[42]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_43.INIT1 = 16'haaa0;
    defparam _add_1_3807_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_41 (.A0(\phase_increment[0] [39]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [40]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17650), .COUT(n17651), .S0(phase_increment_1__63__N_18[39]), 
          .S1(phase_increment_1__63__N_18[40]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_41.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_41.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_39 (.A0(\phase_increment[0] [37]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [38]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17649), .COUT(n17650), .S0(phase_increment_1__63__N_18[37]), 
          .S1(phase_increment_1__63__N_18[38]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_39.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_39.INJECT1_1 = "NO";
    PFUMX i8639 (.BLUT(n19683), .ALUT(n19682), .C0(rx_byte[2]), .Z(n19684));
    LUT4 i4890_4_lut_4_lut (.A(rx_byte[3]), .B(rx_byte[0]), .C(phase_increment_1__63__N_18[55]), 
         .D(phase_increment_1__63__N_16[55]), .Z(n1814)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(265[5] 289[6])
    defparam i4890_4_lut_4_lut.init = 16'hf7d5;
    PFUMX mux_2688_i1 (.BLUT(n4358), .ALUT(n4355), .C0(n19822), .Z(n4361));
    PFUMX mux_2653_i1 (.BLUT(n4311), .ALUT(n4308), .C0(n19822), .Z(n4314));
    PFUMX mux_1704_i1 (.BLUT(n3031), .ALUT(n3016), .C0(rx_byte[2]), .Z(n3039));
    PFUMX i8763 (.BLUT(n19856), .ALUT(n19857), .C0(rx_byte[4]), .Z(n45));
    CCU2C _add_1_3633_add_4_29 (.A0(comb7[62]), .B0(cout_adj_6543), .C0(n105_adj_5901), 
          .D0(n11_adj_5393), .A1(comb7[63]), .B1(cout_adj_6543), .C1(n102_adj_5900), 
          .D1(n10_adj_5392), .CIN(n17317), .COUT(n17318), .S0(comb8_71__N_2137[62]), 
          .S1(comb8_71__N_2137[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_29.INJECT1_1 = "NO";
    PFUMX i8636 (.BLUT(n19680), .ALUT(n19679), .C0(rx_byte[2]), .Z(n19681));
    CCU2C square_sum_add_4_16 (.A0(q_squared[14]), .B0(i_squared[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(q_squared[15]), .B1(i_squared[15]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17492), .COUT(n17493), .S0(n84), .S1(n81));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_16.INIT0 = 16'h666a;
    defparam square_sum_add_4_16.INIT1 = 16'h666a;
    defparam square_sum_add_4_16.INJECT1_0 = "NO";
    defparam square_sum_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_37 (.A0(\phase_increment[0] [35]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [36]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17648), .COUT(n17649), .S0(phase_increment_1__63__N_18[35]), 
          .S1(phase_increment_1__63__N_18[36]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_3807_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_35 (.A0(\phase_increment[0] [33]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [34]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17647), .COUT(n17648), .S0(phase_increment_1__63__N_18[33]), 
          .S1(phase_increment_1__63__N_18[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_35.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_35.INIT1 = 16'haaa0;
    defparam _add_1_3807_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3615_add_4_12 (.A0(amdemod_out_d_11__N_2399[7]), .B0(square_sum[25]), 
          .C0(n30_adj_6282), .D0(n13890), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2399[8]), .D1(VCC_net), .CIN(n17425), 
          .COUT(n17426), .S0(n51_adj_6464), .S1(n48_adj_6463));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3615_add_4_12.INIT0 = 16'h596a;
    defparam _add_1_3615_add_4_12.INIT1 = 16'he1e1;
    defparam _add_1_3615_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3615_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_33 (.A0(\phase_increment[0] [31]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [32]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17646), .COUT(n17647), .S0(phase_increment_1__63__N_18[31]), 
          .S1(phase_increment_1__63__N_18[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_33.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_33.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_31 (.A0(\phase_increment[0] [29]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [30]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17645), .COUT(n17646), .S0(phase_increment_1__63__N_18[29]), 
          .S1(phase_increment_1__63__N_18[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_31.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_31.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_29 (.A0(\phase_increment[0] [27]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [28]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17644), .COUT(n17645), .S0(phase_increment_1__63__N_18[27]), 
          .S1(phase_increment_1__63__N_18[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_29.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_29.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_8 (.A0(integrator5_adj_6562[41]), .B0(integrator4_adj_6561[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[42]), .B1(integrator4_adj_6561[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17405), .COUT(n17406), .S0(n168_adj_6504), 
          .S1(n165_adj_6503));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_27 (.A0(\phase_increment[0] [25]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [26]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17643), .COUT(n17644), .S0(phase_increment_1__63__N_18[25]), 
          .S1(phase_increment_1__63__N_18[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_27.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_27.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_14 (.A0(q_squared[12]), .B0(i_squared[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(q_squared[13]), .B1(i_squared[13]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17491), .COUT(n17492), .S0(n90), .S1(n87));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_14.INIT0 = 16'h666a;
    defparam square_sum_add_4_14.INIT1 = 16'h666a;
    defparam square_sum_add_4_14.INJECT1_0 = "NO";
    defparam square_sum_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_7 (.A0(comb7[40]), .B0(cout_adj_6543), .C0(n171_adj_5923), 
          .D0(n33_adj_5415), .A1(comb7[41]), .B1(cout_adj_6543), .C1(n168_adj_5922), 
          .D1(n32_adj_5414), .CIN(n17306), .COUT(n17307), .S0(comb8_71__N_2137[40]), 
          .S1(comb8_71__N_2137[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_7.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_12 (.A0(q_squared[10]), .B0(i_squared[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(q_squared[11]), .B1(i_squared[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17490), .COUT(n17491), .S0(n96_adj_5610), 
          .S1(n93_adj_5611));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_12.INIT0 = 16'h666a;
    defparam square_sum_add_4_12.INIT1 = 16'h666a;
    defparam square_sum_add_4_12.INJECT1_0 = "NO";
    defparam square_sum_add_4_12.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_10 (.A0(q_squared[8]), .B0(i_squared[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(q_squared[9]), .B1(i_squared[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17489), .COUT(n17490), .S0(n102_adj_5608), 
          .S1(n99_adj_5609));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_10.INIT0 = 16'h666a;
    defparam square_sum_add_4_10.INIT1 = 16'h666a;
    defparam square_sum_add_4_10.INJECT1_0 = "NO";
    defparam square_sum_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_31 (.A0(comb8[64]), .B0(cout_adj_6544), .C0(n99_adj_5862), 
          .D0(n9_adj_5427), .A1(comb8[65]), .B1(cout_adj_6544), .C1(n96_adj_5861), 
          .D1(n8_adj_5426), .CIN(n17296), .COUT(n17297), .S0(comb9_71__N_2209[64]), 
          .S1(comb9_71__N_2209[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_31.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_8 (.A0(q_squared[6]), .B0(i_squared[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(q_squared[7]), .B1(i_squared[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17488), .COUT(n17489), .S0(n108_adj_5606), 
          .S1(n105_adj_5607));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_8.INIT0 = 16'h666a;
    defparam square_sum_add_4_8.INIT1 = 16'h666a;
    defparam square_sum_add_4_8.INJECT1_0 = "NO";
    defparam square_sum_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_21 (.A0(comb8[54]), .B0(cout_adj_6544), .C0(n129_adj_5872), 
          .D0(n19_adj_5437), .A1(comb8[55]), .B1(cout_adj_6544), .C1(n126_adj_5871), 
          .D1(n18_adj_5436), .CIN(n17291), .COUT(n17292), .S0(comb9_71__N_2209[54]), 
          .S1(comb9_71__N_2209[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_21.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_6 (.A0(q_squared[4]), .B0(i_squared[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(q_squared[5]), .B1(i_squared[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17487), .COUT(n17488), .S0(n114_adj_5604), 
          .S1(n111_adj_5605));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_6.INIT0 = 16'h666a;
    defparam square_sum_add_4_6.INIT1 = 16'h666a;
    defparam square_sum_add_4_6.INJECT1_0 = "NO";
    defparam square_sum_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_13 (.A0(comb8[46]), .B0(cout_adj_6544), .C0(n153_adj_5880), 
          .D0(n27_adj_5445), .A1(comb8[47]), .B1(cout_adj_6544), .C1(n150_adj_5879), 
          .D1(n26_adj_5444), .CIN(n17287), .COUT(n17288), .S0(comb9_71__N_2209[46]), 
          .S1(comb9_71__N_2209[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_13.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_4 (.A0(q_squared[2]), .B0(i_squared[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(q_squared[3]), .B1(i_squared[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17486), .COUT(n17487), .S0(n120_adj_5602), 
          .S1(n117_adj_5603));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_4.INIT0 = 16'h666a;
    defparam square_sum_add_4_4.INIT1 = 16'h666a;
    defparam square_sum_add_4_4.INJECT1_0 = "NO";
    defparam square_sum_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_5 (.A0(comb8[38]), .B0(cout_adj_6544), .C0(n177_adj_5888), 
          .D0(n35_adj_5453), .A1(comb8[39]), .B1(cout_adj_6544), .C1(n174_adj_5887), 
          .D1(n34_adj_5452), .CIN(n17283), .COUT(n17284), .S0(comb9_71__N_2209[38]), 
          .S1(comb9_71__N_2209[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_5.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_2 (.A0(q_squared[0]), .B0(i_squared[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(q_squared[1]), .B1(i_squared[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17486), .S1(n123_adj_5601));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(97[22:43])
    defparam square_sum_add_4_2.INIT0 = 16'h0008;
    defparam square_sum_add_4_2.INIT1 = 16'h666a;
    defparam square_sum_add_4_2.INJECT1_0 = "NO";
    defparam square_sum_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3615_add_4_10 (.A0(n19815), .B0(amdemod_out_d_11__N_2399[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2399[6]), 
          .B1(amdemod_out_d_11__N_2370[11]), .C1(amdemod_out_d_11__N_2363), 
          .D1(amdemod_out_d_11__N_2369[11]), .CIN(n17424), .COUT(n17425), 
          .S0(n57_adj_6466), .S1(n54_adj_6465));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3615_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3615_add_4_10.INIT1 = 16'h656a;
    defparam _add_1_3615_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3615_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3600_add_4_13 (.A0(lo_sinewave[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17484), .S0(n28_adj_6350));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(51[25:37])
    defparam _add_1_3600_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_3600_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_3600_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3600_add_4_13.INJECT1_1 = "NO";
    PFUMX i8633 (.BLUT(n19677), .ALUT(n19676), .C0(rx_byte[2]), .Z(n19678));
    CCU2C _add_1_3807_add_4_25 (.A0(\phase_increment[0] [23]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [24]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17642), .COUT(n17643), .S0(phase_increment_1__63__N_18[23]), 
          .S1(phase_increment_1__63__N_18[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_25.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_25.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_23 (.A0(\phase_increment[0] [21]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [22]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17641), .COUT(n17642), .S0(phase_increment_1__63__N_18[21]), 
          .S1(phase_increment_1__63__N_18[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_23.INIT1 = 16'haaa0;
    defparam _add_1_3807_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_21 (.A0(\phase_increment[0] [19]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [20]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17640), .COUT(n17641), .S0(phase_increment_1__63__N_18[19]), 
          .S1(phase_increment_1__63__N_18[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_21.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_21.INJECT1_1 = "NO";
    PFUMX i8470 (.BLUT(n19448), .ALUT(n19447), .C0(rx_byte[2]), .Z(n19449));
    CCU2C _add_1_3807_add_4_19 (.A0(\phase_increment[0] [17]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [18]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17639), .COUT(n17640), .S0(phase_increment_1__63__N_18[17]), 
          .S1(phase_increment_1__63__N_18[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_19.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_3807_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3621_add_4_30 (.A0(comb_d9[27]), .B0(comb9[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[28]), .B1(comb9[28]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17398), .COUT(n17399));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_17 (.A0(\phase_increment[0] [15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [16]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17638), .COUT(n17639), .S0(phase_increment_1__63__N_18[15]), 
          .S1(phase_increment_1__63__N_18[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_3807_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_17.INJECT1_1 = "NO";
    FD1P3AX cic_gain__i1 (.D(cic_gain_7__N_544[0]), .SP(rx_data_valid), 
            .CK(clk_80mhz), .Q(cic_gain[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(260[8] 290[4])
    defparam cic_gain__i1.GSR = "ENABLED";
    CCU2C _add_1_3600_add_4_11 (.A0(lo_sinewave[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_sinewave[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17483), .COUT(n17484), .S0(n34_adj_6352), 
          .S1(n31_adj_6351));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(51[25:37])
    defparam _add_1_3600_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_3600_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_3600_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3600_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_15 (.A0(\phase_increment[0] [13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17637), .COUT(n17638), .S0(phase_increment_1__63__N_18[13]), 
          .S1(phase_increment_1__63__N_18[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3807_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_13 (.A0(\phase_increment[0] [11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17636), .COUT(n17637), .S0(phase_increment_1__63__N_18[11]), 
          .S1(phase_increment_1__63__N_18[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_13.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3807_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_13.INJECT1_1 = "NO";
    GSR GSR_INST (.GSR(VCC_net));
    CCU2C _add_1_3807_add_4_11 (.A0(\phase_increment[0] [9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17635), .COUT(n17636), .S0(phase_increment_1__63__N_18[9]), 
          .S1(phase_increment_1__63__N_18[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3807_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3621_add_4_28 (.A0(comb_d9[25]), .B0(comb9[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[26]), .B1(comb9[26]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17397), .COUT(n17398));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_9 (.A0(\phase_increment[0] [7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17634), .COUT(n17635), .S0(phase_increment_1__63__N_18[7]), 
          .S1(phase_increment_1__63__N_18[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_9.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_6 (.A0(integrator5_adj_6562[39]), .B0(integrator4_adj_6561[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[40]), .B1(integrator4_adj_6561[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17404), .COUT(n17405), .S0(n174_adj_6506), 
          .S1(n171_adj_6505));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_7 (.A0(\phase_increment[0] [5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17633), .COUT(n17634), .S0(phase_increment_1__63__N_18[5]), 
          .S1(phase_increment_1__63__N_18[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_3807_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_5 (.A0(phase_increment_1__63__N_17[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17632), .COUT(n17633), .S0(phase_increment_1__63__N_18[3]), 
          .S1(phase_increment_1__63__N_18[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_5.INIT0 = 16'h555f;
    defparam _add_1_3807_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_3807_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3615_add_4_8 (.A0(n19813), .B0(amdemod_out_d_11__N_2399[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2399[4]), 
          .B1(amdemod_out_d_11__N_2380[14]), .C1(n19815), .D1(amdemod_out_d_11__N_2379[14]), 
          .CIN(n17423), .COUT(n17424), .S0(n63_adj_6468), .S1(n60_adj_6467));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3615_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3615_add_4_8.INIT1 = 16'h656a;
    defparam _add_1_3615_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3615_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3600_add_4_9 (.A0(lo_sinewave[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_sinewave[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17482), .COUT(n17483), .S0(n40_adj_6354), 
          .S1(n37_adj_6353));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(51[25:37])
    defparam _add_1_3600_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_3600_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_3600_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3600_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_3 (.A0(phase_increment_1__63__N_17[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_increment_1__63__N_17[2]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17631), .COUT(n17632), 
          .S0(phase_increment_1__63__N_18[1]), .S1(phase_increment_1__63__N_18[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_3807_add_4_3.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_4 (.A0(integrator5_adj_6562[37]), .B0(integrator4_adj_6561[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[38]), .B1(integrator4_adj_6561[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17403), .COUT(n17404), .S0(n180_adj_6508), 
          .S1(n177_adj_6507));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3807_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_increment_1__63__N_21[0]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .COUT(n17631), .S1(phase_increment_1__63__N_18[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(284[40:78])
    defparam _add_1_3807_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3807_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3807_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3807_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_63 (.A0(\phase_increment[0] [62]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [63]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17629), .S0(phase_increment_1__63__N_20[62]), 
          .S1(phase_increment_1__63__N_20[63]));
    defparam _add_1_3813_add_4_63.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_63.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_63.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_63.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5_adj_6562[36]), .B1(integrator4_adj_6561[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n17403), .S1(n183_adj_6509));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3618_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_61 (.A0(\phase_increment[0] [60]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [61]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17628), .COUT(n17629), .S0(phase_increment_1__63__N_20[60]), 
          .S1(phase_increment_1__63__N_20[61]));
    defparam _add_1_3813_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_61.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_61.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_59 (.A0(\phase_increment[0] [58]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [59]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17627), .COUT(n17628), .S0(phase_increment_1__63__N_20[58]), 
          .S1(phase_increment_1__63__N_20[59]));
    defparam _add_1_3813_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_3621_add_4_38 (.A0(comb_d9[35]), .B0(comb9[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17402), .S1(cout_adj_6511));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3621_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3600_add_4_7 (.A0(lo_sinewave[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_sinewave[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17481), .COUT(n17482), .S0(n46_adj_6356), 
          .S1(n43_adj_6355));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(51[25:37])
    defparam _add_1_3600_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_3600_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_3600_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3600_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3600_add_4_5 (.A0(lo_sinewave[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_sinewave[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17480), .COUT(n17481), .S0(n52_adj_6358), 
          .S1(n49_adj_6357));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(51[25:37])
    defparam _add_1_3600_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_3600_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_3600_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3600_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_19 (.A0(comb7[52]), .B0(cout_adj_6543), .C0(n135_adj_5911), 
          .D0(n21_adj_5403), .A1(comb7[53]), .B1(cout_adj_6543), .C1(n132_adj_5910), 
          .D1(n20_adj_5402), .CIN(n17312), .COUT(n17313), .S0(comb8_71__N_2137[52]), 
          .S1(comb8_71__N_2137[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3600_add_4_3 (.A0(lo_sinewave[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_sinewave[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17479), .COUT(n17480), .S0(n58_adj_6360), 
          .S1(n55_adj_6359));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(51[25:37])
    defparam _add_1_3600_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_3600_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_3600_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3600_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_21 (.A0(comb7[54]), .B0(cout_adj_6543), .C0(n129_adj_5909), 
          .D0(n19_adj_5401), .A1(comb7[55]), .B1(cout_adj_6543), .C1(n126_adj_5908), 
          .D1(n18_adj_5400), .CIN(n17313), .COUT(n17314), .S0(comb8_71__N_2137[54]), 
          .S1(comb8_71__N_2137[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3600_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_sinewave[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17479), .S1(n61_adj_6361));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(51[25:37])
    defparam _add_1_3600_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3600_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_3600_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3600_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_15 (.A0(comb7[48]), .B0(cout_adj_6543), .C0(n147_adj_5915), 
          .D0(n25_adj_5407), .A1(comb7[49]), .B1(cout_adj_6543), .C1(n144_adj_5914), 
          .D1(n24_adj_5406), .CIN(n17310), .COUT(n17311), .S0(comb8_71__N_2137[48]), 
          .S1(comb8_71__N_2137[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3603_add_4_13 (.A0(lo_cosinewave[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17478), .S0(n28_adj_6362));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(52[25:39])
    defparam _add_1_3603_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_3603_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_3603_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3603_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_17 (.A0(comb7[50]), .B0(cout_adj_6543), .C0(n141_adj_5913), 
          .D0(n23_adj_5405), .A1(comb7[51]), .B1(cout_adj_6543), .C1(n138_adj_5912), 
          .D1(n22_adj_5404), .CIN(n17311), .COUT(n17312), .S0(comb8_71__N_2137[50]), 
          .S1(comb8_71__N_2137[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_9 (.A0(comb7[42]), .B0(cout_adj_6543), .C0(n165_adj_5921), 
          .D0(n31_adj_5413), .A1(comb7[43]), .B1(cout_adj_6543), .C1(n162_adj_5920), 
          .D1(n30_adj_5412), .CIN(n17307), .COUT(n17308), .S0(comb8_71__N_2137[42]), 
          .S1(comb8_71__N_2137[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3603_add_4_11 (.A0(lo_cosinewave[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_cosinewave[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17477), .COUT(n17478), .S0(n34_adj_6364), 
          .S1(n31_adj_6363));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(52[25:39])
    defparam _add_1_3603_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_3603_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_3603_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3603_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_11 (.A0(comb7[44]), .B0(cout_adj_6543), .C0(n159_adj_5919), 
          .D0(n29_adj_5411), .A1(comb7[45]), .B1(cout_adj_6543), .C1(n156_adj_5918), 
          .D1(n28_adj_5410), .CIN(n17308), .COUT(n17309), .S0(comb8_71__N_2137[44]), 
          .S1(comb8_71__N_2137[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3603_add_4_9 (.A0(lo_cosinewave[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_cosinewave[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17476), .COUT(n17477), .S0(n40_adj_6366), 
          .S1(n37_adj_6365));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(52[25:39])
    defparam _add_1_3603_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_3603_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_3603_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3603_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3615_add_4_6 (.A0(n19811), .B0(amdemod_out_d_11__N_2399[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2399[2]), 
          .B1(amdemod_out_d_11__N_2390[14]), .C1(n19813), .D1(amdemod_out_d_11__N_2389[14]), 
          .CIN(n17422), .COUT(n17423), .S0(n69_adj_6470), .S1(n66_adj_6469));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3615_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3615_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_3615_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3615_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_28 (.A0(integrator4_adj_6561[61]), .B0(integrator3_adj_6560[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[62]), .B1(integrator3_adj_6560[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17441), .COUT(n17442), .S0(n108_adj_6434), 
          .S1(n105_adj_6433));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3603_add_4_7 (.A0(lo_cosinewave[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_cosinewave[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17475), .COUT(n17476), .S0(n46_adj_6368), 
          .S1(n43_adj_6367));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(52[25:39])
    defparam _add_1_3603_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_3603_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_3603_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3603_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_13 (.A0(comb7[46]), .B0(cout_adj_6543), .C0(n153_adj_5917), 
          .D0(n27_adj_5409), .A1(comb7[47]), .B1(cout_adj_6543), .C1(n150_adj_5916), 
          .D1(n26_adj_5408), .CIN(n17309), .COUT(n17310), .S0(comb8_71__N_2137[46]), 
          .S1(comb8_71__N_2137[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_13.INJECT1_1 = "NO";
    L6MUX21 i8625 (.D0(n19667), .D1(n19664), .SD(n19822), .Z(n19668));
    PFUMX i8623 (.BLUT(n19666), .ALUT(n19665), .C0(led_0_6), .Z(n19667));
    PFUMX i8620 (.BLUT(n19663), .ALUT(n19662), .C0(rx_byte[2]), .Z(n19664));
    CCU2C _add_1_3603_add_4_5 (.A0(lo_cosinewave[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_cosinewave[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17474), .COUT(n17475), .S0(n52_adj_6370), 
          .S1(n49_adj_6369));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(52[25:39])
    defparam _add_1_3603_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_3603_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_3603_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3603_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_6543), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17304));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3633_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3633_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3603_add_4_3 (.A0(lo_cosinewave[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_cosinewave[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17473), .COUT(n17474), .S0(n58_adj_6372), 
          .S1(n55_adj_6371));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(52[25:39])
    defparam _add_1_3603_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_3603_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_3603_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3603_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_5 (.A0(comb7[38]), .B0(cout_adj_6543), .C0(n177_adj_5925), 
          .D0(n35_adj_5417), .A1(comb7[39]), .B1(cout_adj_6543), .C1(n174_adj_5924), 
          .D1(n34_adj_5416), .CIN(n17305), .COUT(n17306), .S0(comb8_71__N_2137[38]), 
          .S1(comb8_71__N_2137[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3633_add_4_3 (.A0(comb7[36]), .B0(cout_adj_6543), .C0(n183_adj_5927), 
          .D0(n37_adj_5419), .A1(comb7[37]), .B1(cout_adj_6543), .C1(n180_adj_5926), 
          .D1(n36_adj_5418), .CIN(n17304), .COUT(n17305), .S0(comb8_71__N_2137[36]), 
          .S1(comb8_71__N_2137[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam _add_1_3633_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3633_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3633_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3633_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_33 (.A0(comb8[66]), .B0(cout_adj_6544), .C0(n93_adj_5860), 
          .D0(n7_adj_5425), .A1(comb8[67]), .B1(cout_adj_6544), .C1(n90_adj_5859), 
          .D1(n6_adj_5424), .CIN(n17297), .COUT(n17298), .S0(comb9_71__N_2209[66]), 
          .S1(comb9_71__N_2209[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3603_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_cosinewave[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17473), .S1(n61_adj_6373));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(52[25:39])
    defparam _add_1_3603_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3603_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_3603_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3603_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_35 (.A0(comb8[68]), .B0(cout_adj_6544), .C0(n87_adj_5858), 
          .D0(n5_adj_5423), .A1(comb8[69]), .B1(cout_adj_6544), .C1(n84_adj_5857), 
          .D1(n4_adj_5422), .CIN(n17298), .COUT(n17299), .S0(comb9_71__N_2209[68]), 
          .S1(comb9_71__N_2209[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3606_add_4_16 (.A0(amdemod_out_d_11__N_2400[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2400[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17471), .S1(n36_adj_6374));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3606_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_3606_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3606_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3606_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3615_add_4_4 (.A0(n19810), .B0(square_sum[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_out_d_11__N_2399[0]), .B1(amdemod_out_d_11__N_2400[14]), 
          .C1(n19811), .D1(amdemod_out_d_11__N_2399[14]), .CIN(n17421), 
          .COUT(n17422), .S0(n75_adj_6472), .S1(n72_adj_6471));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3615_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3615_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_3615_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3615_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_26 (.A0(integrator4_adj_6561[59]), .B0(integrator3_adj_6560[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[60]), .B1(integrator3_adj_6560[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17440), .COUT(n17441), .S0(n114_adj_6436), 
          .S1(n111_adj_6435));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3606_add_4_14 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2400[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2400[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17470), .COUT(n17471), 
          .S0(n45_adj_6376), .S1(n42_adj_6375));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3606_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3606_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_3606_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3606_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_37 (.A0(comb8[70]), .B0(cout_adj_6544), .C0(n81_adj_5856), 
          .D0(n3_adj_5421), .A1(comb8[71]), .B1(cout_adj_6544), .C1(n78_adj_5855), 
          .D1(n2_adj_5420), .CIN(n17299), .S0(comb9_71__N_2209[70]), .S1(comb9_71__N_2209[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_23 (.A0(comb8[56]), .B0(cout_adj_6544), .C0(n123_adj_5870), 
          .D0(n17_adj_5435), .A1(comb8[57]), .B1(cout_adj_6544), .C1(n120_adj_5869), 
          .D1(n16_adj_5434), .CIN(n17292), .COUT(n17293), .S0(comb9_71__N_2209[56]), 
          .S1(comb9_71__N_2209[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3606_add_4_12 (.A0(amdemod_out_d_11__N_2400[7]), .B0(square_sum[25]), 
          .C0(n30_adj_6282), .D0(n13890), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2400[8]), .D1(VCC_net), .CIN(n17469), 
          .COUT(n17470), .S0(n51_adj_6378), .S1(n48_adj_6377));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3606_add_4_12.INIT0 = 16'h596a;
    defparam _add_1_3606_add_4_12.INIT1 = 16'he1e1;
    defparam _add_1_3606_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3606_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_25 (.A0(comb8[58]), .B0(cout_adj_6544), .C0(n117_adj_5868), 
          .D0(n15_adj_5433), .A1(comb8[59]), .B1(cout_adj_6544), .C1(n114_adj_5867), 
          .D1(n14_adj_5432), .CIN(n17293), .COUT(n17294), .S0(comb9_71__N_2209[58]), 
          .S1(comb9_71__N_2209[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3606_add_4_10 (.A0(n19815), .B0(amdemod_out_d_11__N_2400[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2400[6]), 
          .B1(amdemod_out_d_11__N_2370[11]), .C1(amdemod_out_d_11__N_2363), 
          .D1(amdemod_out_d_11__N_2369[11]), .CIN(n17468), .COUT(n17469), 
          .S0(n57_adj_6380), .S1(n54_adj_6379));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3606_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3606_add_4_10.INIT1 = 16'h656a;
    defparam _add_1_3606_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3606_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_29 (.A0(comb8[62]), .B0(cout_adj_6544), .C0(n105_adj_5864), 
          .D0(n11_adj_5429), .A1(comb8[63]), .B1(cout_adj_6544), .C1(n102_adj_5863), 
          .D1(n10_adj_5428), .CIN(n17295), .COUT(n17296), .S0(comb9_71__N_2209[62]), 
          .S1(comb9_71__N_2209[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_27 (.A0(comb8[60]), .B0(cout_adj_6544), .C0(n111_adj_5866), 
          .D0(n13_adj_5431), .A1(comb8[61]), .B1(cout_adj_6544), .C1(n108_adj_5865), 
          .D1(n12_adj_5430), .CIN(n17294), .COUT(n17295), .S0(comb9_71__N_2209[60]), 
          .S1(comb9_71__N_2209[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_15 (.A0(comb8[48]), .B0(cout_adj_6544), .C0(n147_adj_5878), 
          .D0(n25_adj_5443), .A1(comb8[49]), .B1(cout_adj_6544), .C1(n144_adj_5877), 
          .D1(n24_adj_5442), .CIN(n17288), .COUT(n17289), .S0(comb9_71__N_2209[48]), 
          .S1(comb9_71__N_2209[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3606_add_4_8 (.A0(n19813), .B0(amdemod_out_d_11__N_2400[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2400[4]), 
          .B1(amdemod_out_d_11__N_2380[14]), .C1(n19815), .D1(amdemod_out_d_11__N_2379[14]), 
          .CIN(n17467), .COUT(n17468), .S0(n63_adj_6382), .S1(n60_adj_6381));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3606_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3606_add_4_8.INIT1 = 16'h656a;
    defparam _add_1_3606_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3606_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_17 (.A0(comb8[50]), .B0(cout_adj_6544), .C0(n141_adj_5876), 
          .D0(n23_adj_5441), .A1(comb8[51]), .B1(cout_adj_6544), .C1(n138_adj_5875), 
          .D1(n22_adj_5440), .CIN(n17289), .COUT(n17290), .S0(comb9_71__N_2209[50]), 
          .S1(comb9_71__N_2209[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3606_add_4_6 (.A0(n19811), .B0(amdemod_out_d_11__N_2400[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2400[2]), 
          .B1(amdemod_out_d_11__N_2390[14]), .C1(n19813), .D1(amdemod_out_d_11__N_2389[14]), 
          .CIN(n17466), .COUT(n17467), .S0(n69_adj_6384), .S1(n66_adj_6383));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3606_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3606_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_3606_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3606_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_19 (.A0(comb8[52]), .B0(cout_adj_6544), .C0(n135_adj_5874), 
          .D0(n21_adj_5439), .A1(comb8[53]), .B1(cout_adj_6544), .C1(n132_adj_5873), 
          .D1(n20_adj_5438), .CIN(n17290), .COUT(n17291), .S0(comb9_71__N_2209[52]), 
          .S1(comb9_71__N_2209[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_19.INJECT1_1 = "NO";
    L6MUX21 i8467 (.D0(n19445), .D1(n19442), .SD(n19822), .Z(n19446));
    CCU2C _add_1_3636_add_4_7 (.A0(comb8[40]), .B0(cout_adj_6544), .C0(n171_adj_5886), 
          .D0(n33_adj_5451), .A1(comb8[41]), .B1(cout_adj_6544), .C1(n168_adj_5885), 
          .D1(n32_adj_5450), .CIN(n17284), .COUT(n17285), .S0(comb9_71__N_2209[40]), 
          .S1(comb9_71__N_2209[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3606_add_4_4 (.A0(n19810), .B0(square_sum[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_out_d_11__N_2400[0]), .B1(amdemod_out_d_11__N_2400[14]), 
          .C1(n19811), .D1(amdemod_out_d_11__N_2399[14]), .CIN(n17465), 
          .COUT(n17466), .S0(n75_adj_6386), .S1(n72_adj_6385));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3606_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3606_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_3606_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3606_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_9 (.A0(comb8[42]), .B0(cout_adj_6544), .C0(n165_adj_5884), 
          .D0(n31_adj_5449), .A1(comb8[43]), .B1(cout_adj_6544), .C1(n162_adj_5883), 
          .D1(n30_adj_5448), .CIN(n17285), .COUT(n17286), .S0(comb9_71__N_2209[42]), 
          .S1(comb9_71__N_2209[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3606_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17465), .S1(n78_adj_6387));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3606_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3606_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3606_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3606_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_11 (.A0(comb8[44]), .B0(cout_adj_6544), .C0(n159_adj_5882), 
          .D0(n29_adj_5447), .A1(comb8[45]), .B1(cout_adj_6544), .C1(n156_adj_5881), 
          .D1(n28_adj_5446), .CIN(n17286), .COUT(n17287), .S0(comb9_71__N_2209[44]), 
          .S1(comb9_71__N_2209[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_38 (.A0(integrator3_adj_6560[71]), .B0(integrator2_adj_6559[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17464), .S0(n78_adj_6388));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3609_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_38.INJECT1_1 = "NO";
    AMDemodulator AMDemodulator_inst (.cic_sine_clk(cic_sine_clk), .led_0_2(led_0_2), 
            .led_0_1(led_0_1), .n51(n51), .n51_adj_229(n51_adj_6517), 
            .n19813(n19813), .\amdemod_out_d_11__N_2379[14] (amdemod_out_d_11__N_2379[14]), 
            .\amdemod_out_d_11__N_2380[14] (amdemod_out_d_11__N_2380[14]), 
            .n19815(n19815), .led_0_0(led_0_0), .\cic_sine_out[5] (cic_sine_out[5]), 
            .n19816(n19816), .\cic_sine_out[4] (cic_sine_out[4]), .\cic_sine_out[3] (cic_sine_out[3]), 
            .\cic_sine_out[2] (cic_sine_out[2]), .\cic_sine_out[1] (cic_sine_out[1]), 
            .\data_in_reg_11__N_2898[7] (data_in_reg_11__N_2898[7]), .n46(n46_adj_6080), 
            .n46_adj_230(n46_adj_6066), .n48(n48), .n48_adj_231(n48_adj_6516), 
            .n43(n43_adj_6079), .n43_adj_232(n43_adj_6065), .n45(n45_adj_5665), 
            .n45_adj_233(n45_adj_6515), .n40(n40_adj_6078), .n40_adj_234(n40_adj_6064), 
            .n42(n42), .n42_adj_235(n42_adj_6514), .cic_cosine_out({cic_cosine_out}), 
            .\data_in_reg_11__N_2898[6] (data_in_reg_11__N_2898[6]), .n76(n76_adj_6062), 
            .n76_adj_236(n76_adj_6048), .n19811(n19811), .\data_in_reg_11__N_2898[5] (data_in_reg_11__N_2898[5]), 
            .\data_in_reg_11__N_2898[4] (data_in_reg_11__N_2898[4]), .\data_in_reg_11__N_2898[3] (data_in_reg_11__N_2898[3]), 
            .\data_in_reg_11__N_2898[2] (data_in_reg_11__N_2898[2]), .\data_in_reg_11__N_2898[1] (data_in_reg_11__N_2898[1]), 
            .n78(n78_adj_6473), .n78_adj_237(n78_adj_6387), .n73(n73_adj_6061), 
            .n73_adj_238(n73), .n75(n75_adj_6472), .n75_adj_239(n75_adj_6386), 
            .\cic_sine_out[0] (cic_sine_out[0]), .n70(n70_adj_6060), .n70_adj_240(n70_adj_6047), 
            .n72(n72_adj_6471), .n72_adj_241(n72_adj_6385), .n67(n67_adj_6059), 
            .n67_adj_242(n67_adj_6046), .n69(n69_adj_6470), .n69_adj_243(n69_adj_6384), 
            .n64(n64_adj_6058), .n64_adj_244(n64_adj_6045), .n66(n66_adj_6469), 
            .n66_adj_245(n66_adj_6383), .\data_in_reg_11__N_2898[0] (data_in_reg_11__N_2898[0]), 
            .n61(n61_adj_6057), .n61_adj_246(n61_adj_6044), .n63(n63_adj_6468), 
            .n63_adj_247(n63_adj_6382), .led_0_4(led_0_4), .led_0_5(led_0_5), 
            .n58(n58_adj_6056), .n58_adj_248(n58_adj_6043), .n36(n36_adj_5841), 
            .n36_adj_249(n36_adj_5811), .amdemod_out_d_11__N_2363(amdemod_out_d_11__N_2363), 
            .n60(n60_adj_6467), .n60_adj_250(n60_adj_6381), .n34(n34_adj_6185), 
            .n34_adj_251(n34_adj_6171), .n55(n55_adj_6055), .n55_adj_252(n55_adj_6042), 
            .n57(n57_adj_6466), .n57_adj_253(n57_adj_6380), .n52(n52_adj_6054), 
            .n52_adj_254(n52_adj_6041), .n54(n54_adj_6465), .n54_adj_255(n54_adj_6379), 
            .n36_adj_256(n36_adj_5797), .n36_adj_257(n36_adj_5711), .n49(n49_adj_6053), 
            .n49_adj_258(n49_adj_6040), .n34_adj_259(n34_adj_6157), .n34_adj_260(n34_adj_6143), 
            .n51_adj_261(n51_adj_6464), .n51_adj_262(n51_adj_6378), .n46_adj_263(n46_adj_6052), 
            .n46_adj_264(n46_adj_6039), .n48_adj_265(n48_adj_6463), .n48_adj_266(n48_adj_6377), 
            .n43_adj_267(n43_adj_6051), .n43_adj_268(n43_adj_6038), .n45_adj_269(n45_adj_6462), 
            .n45_adj_270(n45_adj_6376), .n40_adj_271(n40_adj_6050), .n40_adj_272(n40_adj_6037), 
            .n42_adj_273(n42_adj_6461), .n42_adj_274(n42_adj_6375), .n76_adj_275(n76_adj_6198), 
            .n76_adj_276(n76_adj_6184), .n36_adj_277(n36_adj_5664), .n36_adj_278(n36_adj_6513), 
            .n78_adj_279(n78_adj_5854), .n78_adj_280(n78_adj_5824), .n34_adj_281(n34_adj_6077), 
            .n34_adj_282(n34_adj_6063), .n36_adj_283(n36_adj_6460), .n36_adj_284(n36_adj_6374), 
            .n34_adj_285(n34_adj_6049), .n34_adj_286(n34_adj_6036), .\square_sum[23] (square_sum[23]), 
            .\square_sum[22] (square_sum[22]), .n4(n4_adj_6510), .n34_adj_287(n34_adj_6542), 
            .n34_adj_288(n34_adj_6200), .n19809(n19809), .\amdemod_out_d_11__N_2369[11] (amdemod_out_d_11__N_2369[11]), 
            .\amdemod_out_d_11__N_2370[11] (amdemod_out_d_11__N_2370[11]), 
            .n36_adj_289(n36_adj_6130), .n36_adj_290(n36_adj_5310), .n13878(n13878), 
            .n42_adj_291(n42_adj_6286), .\square_sum[25] (square_sum[25]), 
            .amdemod_out_d_11__N_2516(amdemod_out_d_11__N_2516), .n64_adj_292(n64_adj_6194), 
            .n64_adj_293(n64_adj_6180), .n66_adj_294(n66_adj_5850), .n66_adj_295(n66_adj_5820), 
            .n67_adj_296(n67_adj_6195), .n67_adj_297(n67_adj_6181), .n69_adj_298(n69_adj_5851), 
            .n69_adj_299(n69_adj_5821), .n58_adj_300(n58_adj_6192), .n58_adj_301(n58_adj_6178), 
            .n60_adj_302(n60_adj_5848), .n60_adj_303(n60_adj_5818), .n61_adj_304(n61_adj_6193), 
            .n61_adj_305(n61_adj_6179), .amdemod_out_d_11__N_2594(amdemod_out_d_11__N_2594), 
            .n63_adj_306(n63_adj_5849), .n63_adj_307(n63_adj_5819), .n55_adj_308(n55_adj_6191), 
            .n55_adj_309(n55_adj_6177), .n57_adj_310(n57_adj_5847), .n57_adj_311(n57_adj_5817), 
            .n52_adj_312(n52_adj_6190), .n52_adj_313(n52_adj_6176), .n54_adj_314(n54_adj_5846), 
            .n54_adj_315(n54_adj_5816), .\amdemod_out[9] (amdemod_out[9]), 
            .\data_in_reg_11__N_2898[8] (data_in_reg_11__N_2898[8]), .n39(n39_adj_6285), 
            .\amdemod_out_d_11__N_2365[3] (amdemod_out_d_11__N_2365[3]), .n39_adj_316(n39), 
            .n49_adj_317(n49_adj_6189), .n49_adj_318(n49_adj_6175), .n51_adj_319(n51_adj_5845), 
            .n51_adj_320(n51_adj_5815), .n46_adj_321(n46_adj_6188), .n46_adj_322(n46_adj_6174), 
            .n48_adj_323(n48_adj_5844), .n48_adj_324(n48_adj_5814), .n19810(n19810), 
            .n19828(n19828), .n19827(n19827), .\amdemod_out_d_11__N_2365[14] (amdemod_out_d_11__N_2365[14]), 
            .n24(n24_adj_6237), .n13890(n13890), .n43_adj_325(n43_adj_6187), 
            .n43_adj_326(n43_adj_6173), .n45_adj_327(n45_adj_5843), .n45_adj_328(n45_adj_5813), 
            .n40_adj_329(n40_adj_6186), .n40_adj_330(n40_adj_6172), .n30(n30_adj_6282), 
            .n76_adj_331(n76_adj_6170), .n76_adj_332(n76_adj_6156), .n78_adj_333(n78_adj_5810), 
            .n78_adj_334(n78_adj_5724), .n42_adj_335(n42_adj_5842), .n42_adj_336(n42_adj_5812), 
            .\amdemod_out_d_11__N_2409[14] (amdemod_out_d_11__N_2409[14]), 
            .\amdemod_out_d_11__N_2410[14] (amdemod_out_d_11__N_2410[14]), 
            .n19808(n19808), .\amdemod_out_d_11__N_2365[1] (amdemod_out_d_11__N_2365[1]), 
            .n45_adj_337(n45_adj_6243), .n13876(n13876), .\amdemod_out_d_11__N_2365[6] (amdemod_out_d_11__N_2365[6]), 
            .n30_adj_338(n30_adj_6239), .\amdemod_out_d_11__N_2365[2] (amdemod_out_d_11__N_2365[2]), 
            .n42_adj_339(n42_adj_6242), .amdemod_out_d_11__N_2597(amdemod_out_d_11__N_2597), 
            .n73_adj_340(n73_adj_6197), .n73_adj_341(n73_adj_6183), .n75_adj_342(n75_adj_5853), 
            .n75_adj_343(n75_adj_5823), .n70_adj_344(n70_adj_6196), .n70_adj_345(n70_adj_6182), 
            .n73_adj_346(n73_adj_6169), .n73_adj_347(n73_adj_6155), .n75_adj_348(n75_adj_5809), 
            .n75_adj_349(n75_adj_5723), .n70_adj_350(n70_adj_6168), .n70_adj_351(n70_adj_6154), 
            .n72_adj_352(n72_adj_5808), .n72_adj_353(n72_adj_5722), .n72_adj_354(n72_adj_5852), 
            .n72_adj_355(n72_adj_5822), .n67_adj_356(n67_adj_6167), .n67_adj_357(n67_adj_6153), 
            .\amdemod_out_d_11__N_2358[5] (amdemod_out_d_11__N_2358[5]), .n33(n33_adj_6283), 
            .n69_adj_358(n69_adj_5807), .n69_adj_359(n69_adj_5721), .n64_adj_360(n64_adj_6166), 
            .n64_adj_361(n64_adj_6152), .\amdemod_out_d_11__N_2365[4] (amdemod_out_d_11__N_2365[4]), 
            .n36_adj_362(n36_adj_6241), .\amdemod_out_d_11__N_2365[5] (amdemod_out_d_11__N_2365[5]), 
            .n33_adj_363(n33_adj_6240), .n66_adj_364(n66_adj_5806), .n66_adj_365(n66_adj_5720), 
            .n36_adj_366(n36_adj_6284), .n61_adj_367(n61_adj_6165), .n61_adj_368(n61_adj_6151), 
            .n63_adj_369(n63_adj_5805), .n63_adj_370(n63_adj_5719), .n58_adj_371(n58_adj_6164), 
            .n58_adj_372(n58_adj_6150), .n60_adj_373(n60_adj_5804), .n60_adj_374(n60_adj_5718), 
            .n55_adj_375(n55_adj_6163), .n55_adj_376(n55_adj_6149), .n57_adj_377(n57_adj_5803), 
            .n57_adj_378(n57_adj_5717), .n52_adj_379(n52_adj_6162), .n52_adj_380(n52_adj_6148), 
            .n54_adj_381(n54_adj_5802), .n54_adj_382(n54_adj_5716), .n49_adj_383(n49_adj_6161), 
            .n49_adj_384(n49_adj_6147), .n51_adj_385(n51_adj_5801), .n51_adj_386(n51_adj_5715), 
            .\amdemod_out_d_11__N_2365[7] (amdemod_out_d_11__N_2365[7]), .n27(n27_adj_6238), 
            .amdemod_out_d_11__N_2564(amdemod_out_d_11__N_2564), .n46_adj_387(n46_adj_6160), 
            .n46_adj_388(n46_adj_6146), .n48_adj_389(n48_adj_5800), .n48_adj_390(n48_adj_5714), 
            .amdemod_out_d_11__N_2567(amdemod_out_d_11__N_2567), .n46_adj_391(n46_adj_6199), 
            .n48_adj_392(n48_adj_6244), .n13821(n13821), .n13815(n13815), 
            .n43_adj_393(n43_adj_6159), .n43_adj_394(n43_adj_6145), .amdemod_out_d_11__N_2570(amdemod_out_d_11__N_2570), 
            .\amdemod_out_d_11__N_2399[14] (amdemod_out_d_11__N_2399[14]), 
            .\amdemod_out_d_11__N_2400[14] (amdemod_out_d_11__N_2400[14]), 
            .amdemod_out_d_11__N_2573(amdemod_out_d_11__N_2573), .n45_adj_395(n45_adj_5799), 
            .n45_adj_396(n45_adj_5713), .n40_adj_397(n40_adj_6158), .n40_adj_398(n40_adj_6144), 
            .n42_adj_399(n42_adj_5798), .n42_adj_400(n42_adj_5712), .amdemod_out_d_11__N_2576(amdemod_out_d_11__N_2576), 
            .n76_adj_401(n76_adj_6090), .n76_adj_402(n76_adj_6076), .n19812(n19812), 
            .amdemod_out_d_11__N_2579(amdemod_out_d_11__N_2579), .n78_adj_403(n78_adj_5674), 
            .n78_adj_404(n78_adj_6526), .n73_adj_405(n73_adj_6089), .n73_adj_406(n73_adj_6075), 
            .\amdemod_out_d_11__N_2389[14] (amdemod_out_d_11__N_2389[14]), 
            .\amdemod_out_d_11__N_2390[14] (amdemod_out_d_11__N_2390[14]), 
            .n75_adj_407(n75_adj_5673), .n75_adj_408(n75_adj_6525), .n70_adj_409(n70_adj_6088), 
            .n70_adj_410(n70_adj_6074), .amdemod_out_d_11__N_2585(amdemod_out_d_11__N_2585), 
            .n72_adj_411(n72_adj_5672), .n72_adj_412(n72_adj_6524), .n67_adj_413(n67_adj_6087), 
            .n67_adj_414(n67_adj_6073), .amdemod_out_d_11__N_2582(amdemod_out_d_11__N_2582), 
            .n69_adj_415(n69_adj_5671), .n69_adj_416(n69_adj_6523), .n19824(n19824), 
            .n64_adj_417(n64_adj_6086), .n64_adj_418(n64_adj_6072), .n66_adj_419(n66_adj_5670), 
            .n66_adj_420(n66_adj_6522), .n61_adj_421(n61_adj_6085), .n61_adj_422(n61_adj_6071), 
            .n63_adj_423(n63_adj_5669), .n63_adj_424(n63_adj_6521), .n58_adj_425(n58_adj_6084), 
            .n58_adj_426(n58_adj_6070), .n60_adj_427(n60_adj_5668), .n60_adj_428(n60_adj_6520), 
            .n19814(n19814), .n55_adj_429(n55_adj_6083), .n55_adj_430(n55_adj_6069), 
            .n57_adj_431(n57_adj_5667), .n57_adj_432(n57_adj_6519), .amdemod_out_d_11__N_2591(amdemod_out_d_11__N_2591), 
            .n52_adj_433(n52_adj_6082), .n52_adj_434(n52_adj_6068), .amdemod_out_d_11__N_2588(amdemod_out_d_11__N_2588), 
            .n54_adj_435(n54_adj_5666), .n54_adj_436(n54_adj_6518), .n49_adj_437(n49_adj_6081), 
            .n49_adj_438(n49_adj_6067), .amdemod_out_d_11__N_2600(amdemod_out_d_11__N_2600), 
            .amdemod_out_d_11__N_2798(amdemod_out_d_11__N_2798), .amdemod_out_d_11__N_2801(amdemod_out_d_11__N_2801), 
            .amdemod_out_d_11__N_2804(amdemod_out_d_11__N_2804), .amdemod_out_d_11__N_2807(amdemod_out_d_11__N_2807), 
            .amdemod_out_d_11__N_2810(amdemod_out_d_11__N_2810), .amdemod_out_d_11__N_2813(amdemod_out_d_11__N_2813), 
            .amdemod_out_d_11__N_2816(amdemod_out_d_11__N_2816), .amdemod_out_d_11__N_2819(amdemod_out_d_11__N_2819), 
            .amdemod_out_d_11__N_2822(amdemod_out_d_11__N_2822), .amdemod_out_d_11__N_2825(amdemod_out_d_11__N_2825), 
            .amdemod_out_d_11__N_2828(amdemod_out_d_11__N_2828), .amdemod_out_d_11__N_2831(amdemod_out_d_11__N_2831), 
            .amdemod_out_d_11__N_2834(amdemod_out_d_11__N_2834), .amdemod_out_d_11__N_2720(amdemod_out_d_11__N_2720), 
            .amdemod_out_d_11__N_2723(amdemod_out_d_11__N_2723), .amdemod_out_d_11__N_2726(amdemod_out_d_11__N_2726), 
            .amdemod_out_d_11__N_2729(amdemod_out_d_11__N_2729), .amdemod_out_d_11__N_2732(amdemod_out_d_11__N_2732), 
            .amdemod_out_d_11__N_2735(amdemod_out_d_11__N_2735), .amdemod_out_d_11__N_2738(amdemod_out_d_11__N_2738), 
            .amdemod_out_d_11__N_2741(amdemod_out_d_11__N_2741), .amdemod_out_d_11__N_2744(amdemod_out_d_11__N_2744), 
            .amdemod_out_d_11__N_2747(amdemod_out_d_11__N_2747), .amdemod_out_d_11__N_2750(amdemod_out_d_11__N_2750), 
            .amdemod_out_d_11__N_2753(amdemod_out_d_11__N_2753), .amdemod_out_d_11__N_2756(amdemod_out_d_11__N_2756), 
            .led_0_3(led_0_3), .amdemod_out_d_11__N_2642(amdemod_out_d_11__N_2642), 
            .amdemod_out_d_11__N_2645(amdemod_out_d_11__N_2645), .amdemod_out_d_11__N_2648(amdemod_out_d_11__N_2648), 
            .amdemod_out_d_11__N_2501(amdemod_out_d_11__N_2501), .amdemod_out_d_11__N_2651(amdemod_out_d_11__N_2651), 
            .amdemod_out_d_11__N_2654(amdemod_out_d_11__N_2654), .amdemod_out_d_11__N_2657(amdemod_out_d_11__N_2657), 
            .amdemod_out_d_11__N_2507(amdemod_out_d_11__N_2507), .amdemod_out_d_11__N_2660(amdemod_out_d_11__N_2660), 
            .amdemod_out_d_11__N_2663(amdemod_out_d_11__N_2663), .amdemod_out_d_11__N_2666(amdemod_out_d_11__N_2666), 
            .amdemod_out_d_11__N_2669(amdemod_out_d_11__N_2669), .amdemod_out_d_11__N_2504(amdemod_out_d_11__N_2504), 
            .amdemod_out_d_11__N_2672(amdemod_out_d_11__N_2672), .amdemod_out_d_11__N_2675(amdemod_out_d_11__N_2675), 
            .amdemod_out_d_11__N_2678(amdemod_out_d_11__N_2678), .amdemod_out_d_11__N_2513(amdemod_out_d_11__N_2513), 
            .amdemod_out_d_11__N_2510(amdemod_out_d_11__N_2510), .VCC_net(VCC_net), 
            .GND_net(GND_net), .q_squared({q_squared}), .i_squared({i_squared})) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(219[6] 224[5])
    CCU2C _add_1_3609_add_4_36 (.A0(integrator3_adj_6560[69]), .B0(integrator2_adj_6559[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[70]), .B1(integrator2_adj_6559[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17463), .COUT(n17464), .S0(n84_adj_6390), 
          .S1(n81_adj_6389));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3615_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17421), .S1(n78_adj_6473));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3615_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3615_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3615_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3615_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_24 (.A0(integrator4_adj_6561[57]), .B0(integrator3_adj_6560[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[58]), .B1(integrator3_adj_6560[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17439), .COUT(n17440), .S0(n120_adj_6438), 
          .S1(n117_adj_6437));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_34 (.A0(integrator3_adj_6560[67]), .B0(integrator2_adj_6559[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[68]), .B1(integrator2_adj_6559[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17462), .COUT(n17463), .S0(n90_adj_6392), 
          .S1(n87_adj_6391));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_3 (.A0(comb8[36]), .B0(cout_adj_6544), .C0(n183_adj_5890), 
          .D0(n37_adj_5455), .A1(comb8[37]), .B1(cout_adj_6544), .C1(n180_adj_5889), 
          .D1(n36_adj_5454), .CIN(n17282), .COUT(n17283), .S0(comb9_71__N_2209[36]), 
          .S1(comb9_71__N_2209[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3636_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3636_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3636_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_6544), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17282));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam _add_1_3636_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3636_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3636_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3636_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_32 (.A0(integrator3_adj_6560[65]), .B0(integrator2_adj_6559[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[66]), .B1(integrator2_adj_6559[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17461), .COUT(n17462), .S0(n96_adj_6394), 
          .S1(n93_adj_6393));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_30 (.A0(integrator3_adj_6560[63]), .B0(integrator2_adj_6559[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[64]), .B1(integrator2_adj_6559[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17460), .COUT(n17461), .S0(n102_adj_6396), 
          .S1(n99_adj_6395));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_30.INJECT1_1 = "NO";
    PFUMX i8465 (.BLUT(n19444), .ALUT(n19443), .C0(led_0_6), .Z(n19445));
    CCU2C _add_1_3609_add_4_28 (.A0(integrator3_adj_6560[61]), .B0(integrator2_adj_6559[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[62]), .B1(integrator2_adj_6559[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17459), .COUT(n17460), .S0(n108_adj_6398), 
          .S1(n105_adj_6397));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_26 (.A0(integrator3_adj_6560[59]), .B0(integrator2_adj_6559[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[60]), .B1(integrator2_adj_6559[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17458), .COUT(n17459), .S0(n114_adj_6400), 
          .S1(n111_adj_6399));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_26.INJECT1_1 = "NO";
    LUT4 i4917_4_lut_4_lut (.A(rx_byte[3]), .B(rx_byte[0]), .C(phase_increment_1__63__N_18[49]), 
         .D(phase_increment_1__63__N_16[49]), .Z(n2096)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(265[5] 289[6])
    defparam i4917_4_lut_4_lut.init = 16'hf7d5;
    PFUMX mux_2509_i1 (.BLUT(n4112), .ALUT(n4097), .C0(rx_byte[2]), .Z(n4120));
    PFUMX i8608 (.BLUT(n19648), .ALUT(n19647), .C0(rx_byte[2]), .Z(n19649));
    PFUMX i8603 (.BLUT(n19641), .ALUT(n19640), .C0(rx_byte[2]), .Z(n19642));
    CCU2C _add_1_3813_add_4_57 (.A0(\phase_increment[0] [56]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [57]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17626), .COUT(n17627), .S0(phase_increment_1__63__N_20[56]), 
          .S1(phase_increment_1__63__N_20[57]));
    defparam _add_1_3813_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_22 (.A0(integrator4_adj_6561[55]), .B0(integrator3_adj_6560[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[56]), .B1(integrator3_adj_6560[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17438), .COUT(n17439), .S0(n126_adj_6440), 
          .S1(n123_adj_6439));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_24 (.A0(integrator3_adj_6560[57]), .B0(integrator2_adj_6559[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[58]), .B1(integrator2_adj_6559[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17457), .COUT(n17458), .S0(n120_adj_6402), 
          .S1(n117_adj_6401));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_20 (.A0(integrator4_adj_6561[53]), .B0(integrator3_adj_6560[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[54]), .B1(integrator3_adj_6560[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17437), .COUT(n17438), .S0(n132_adj_6442), 
          .S1(n129_adj_6441));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_22 (.A0(integrator3_adj_6560[55]), .B0(integrator2_adj_6559[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[56]), .B1(integrator2_adj_6559[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17456), .COUT(n17457), .S0(n126_adj_6404), 
          .S1(n123_adj_6403));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_22.INJECT1_1 = "NO";
    LUT4 mux_1667_i1_3_lut (.A(rx_byte[2]), .B(n2964), .C(rx_byte[3]), 
         .Z(n2989)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(274[5] 288[12])
    defparam mux_1667_i1_3_lut.init = 16'hcaca;
    CCU2C _add_1_3618_add_4_38 (.A0(integrator5_adj_6562[71]), .B0(integrator4_adj_6561[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17420), .S0(n78_adj_6474));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3618_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_18 (.A0(integrator4_adj_6561[51]), .B0(integrator3_adj_6560[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[52]), .B1(integrator3_adj_6560[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17436), .COUT(n17437), .S0(n138_adj_6444), 
          .S1(n135_adj_6443));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_20 (.A0(integrator3_adj_6560[53]), .B0(integrator2_adj_6559[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[54]), .B1(integrator2_adj_6559[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17455), .COUT(n17456), .S0(n132_adj_6406), 
          .S1(n129_adj_6405));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_37 (.A0(integrator_tmp[70]), .B0(cout_adj_5271), 
          .C0(n81_adj_5965), .D0(n3), .A1(integrator_tmp[71]), .B1(cout_adj_5271), 
          .C1(n78_adj_5964), .D1(n2), .CIN(n17383), .S0(comb6_71__N_1993[70]), 
          .S1(comb6_71__N_1993[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_55 (.A0(\phase_increment[0] [54]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [55]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17625), .COUT(n17626), .S0(phase_increment_1__63__N_20[54]), 
          .S1(phase_increment_1__63__N_20[55]));
    defparam _add_1_3813_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_3621_add_4_26 (.A0(comb_d9[23]), .B0(comb9[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[24]), .B1(comb9[24]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17396), .COUT(n17397));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3621_add_4_36 (.A0(comb_d9[33]), .B0(comb9[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[34]), .B1(comb9[34]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17401), .COUT(n17402));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_53 (.A0(\phase_increment[0] [52]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [53]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17624), .COUT(n17625), .S0(phase_increment_1__63__N_20[52]), 
          .S1(phase_increment_1__63__N_20[53]));
    defparam _add_1_3813_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_3624_add_4_35 (.A0(integrator_tmp[68]), .B0(cout_adj_5271), 
          .C0(n87_adj_5967), .D0(n5), .A1(integrator_tmp[69]), .B1(cout_adj_5271), 
          .C1(n84_adj_5966), .D1(n4), .CIN(n17382), .COUT(n17383), .S0(comb6_71__N_1993[68]), 
          .S1(comb6_71__N_1993[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam _add_1_3624_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3624_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3624_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3624_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_51 (.A0(\phase_increment[0] [50]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [51]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17623), .COUT(n17624), .S0(phase_increment_1__63__N_20[50]), 
          .S1(phase_increment_1__63__N_20[51]));
    defparam _add_1_3813_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_36 (.A0(integrator5_adj_6562[69]), .B0(integrator4_adj_6561[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[70]), .B1(integrator4_adj_6561[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17419), .COUT(n17420), .S0(n84_adj_6476), 
          .S1(n81_adj_6475));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_16 (.A0(integrator4_adj_6561[49]), .B0(integrator3_adj_6560[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[50]), .B1(integrator3_adj_6560[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17435), .COUT(n17436), .S0(n144_adj_6446), 
          .S1(n141_adj_6445));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_18 (.A0(integrator3_adj_6560[51]), .B0(integrator2_adj_6559[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[52]), .B1(integrator2_adj_6559[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17454), .COUT(n17455), .S0(n138_adj_6408), 
          .S1(n135_adj_6407));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_34 (.A0(integrator5_adj_6562[67]), .B0(integrator4_adj_6561[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[68]), .B1(integrator4_adj_6561[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17418), .COUT(n17419), .S0(n90_adj_6478), 
          .S1(n87_adj_6477));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_14 (.A0(integrator4_adj_6561[47]), .B0(integrator3_adj_6560[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[48]), .B1(integrator3_adj_6560[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17434), .COUT(n17435), .S0(n150_adj_6448), 
          .S1(n147_adj_6447));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_16 (.A0(integrator3_adj_6560[49]), .B0(integrator2_adj_6559[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[50]), .B1(integrator2_adj_6559[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17453), .COUT(n17454), .S0(n144_adj_6410), 
          .S1(n141_adj_6409));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3621_add_4_24 (.A0(comb_d9[21]), .B0(comb9[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[22]), .B1(comb9[22]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17395), .COUT(n17396));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3621_add_4_34 (.A0(comb_d9[31]), .B0(comb9[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[32]), .B1(comb9[32]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17400), .COUT(n17401));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_49 (.A0(\phase_increment[0] [48]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [49]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17622), .COUT(n17623), .S0(phase_increment_1__63__N_20[48]), 
          .S1(phase_increment_1__63__N_20[49]));
    defparam _add_1_3813_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_3621_add_4_32 (.A0(comb_d9[29]), .B0(comb9[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[30]), .B1(comb9[30]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17399), .COUT(n17400));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam _add_1_3621_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_3621_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_3621_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3621_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_32 (.A0(integrator5_adj_6562[65]), .B0(integrator4_adj_6561[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[66]), .B1(integrator4_adj_6561[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17417), .COUT(n17418), .S0(n96_adj_6480), 
          .S1(n93_adj_6479));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_47 (.A0(\phase_increment[0] [46]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [47]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17621), .COUT(n17622), .S0(phase_increment_1__63__N_20[46]), 
          .S1(phase_increment_1__63__N_20[47]));
    defparam _add_1_3813_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_3813_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_45 (.A0(\phase_increment[0] [44]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [45]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17620), .COUT(n17621), .S0(phase_increment_1__63__N_20[44]), 
          .S1(phase_increment_1__63__N_20[45]));
    defparam _add_1_3813_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_45.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_30 (.A0(integrator5_adj_6562[63]), .B0(integrator4_adj_6561[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[64]), .B1(integrator4_adj_6561[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17416), .COUT(n17417), .S0(n102_adj_6482), 
          .S1(n99_adj_6481));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_12 (.A0(integrator4_adj_6561[45]), .B0(integrator3_adj_6560[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[46]), .B1(integrator3_adj_6560[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17433), .COUT(n17434), .S0(n156_adj_6450), 
          .S1(n153_adj_6449));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_14 (.A0(integrator3_adj_6560[47]), .B0(integrator2_adj_6559[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[48]), .B1(integrator2_adj_6559[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17452), .COUT(n17453), .S0(n150_adj_6412), 
          .S1(n147_adj_6411));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_28 (.A0(integrator5_adj_6562[61]), .B0(integrator4_adj_6561[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[62]), .B1(integrator4_adj_6561[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17415), .COUT(n17416), .S0(n108_adj_6484), 
          .S1(n105_adj_6483));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_43 (.A0(\phase_increment[0] [42]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [43]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17619), .COUT(n17620), .S0(phase_increment_1__63__N_20[42]), 
          .S1(phase_increment_1__63__N_20[43]));
    defparam _add_1_3813_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_43.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_12 (.A0(integrator3_adj_6560[45]), .B0(integrator2_adj_6559[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[46]), .B1(integrator2_adj_6559[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17451), .COUT(n17452), .S0(n156_adj_6414), 
          .S1(n153_adj_6413));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_26 (.A0(integrator5_adj_6562[59]), .B0(integrator4_adj_6561[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[60]), .B1(integrator4_adj_6561[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17414), .COUT(n17415), .S0(n114_adj_6486), 
          .S1(n111_adj_6485));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_41 (.A0(\phase_increment[0] [40]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [41]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17618), .COUT(n17619), .S0(phase_increment_1__63__N_20[40]), 
          .S1(phase_increment_1__63__N_20[41]));
    defparam _add_1_3813_add_4_41.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_24 (.A0(integrator5_adj_6562[57]), .B0(integrator4_adj_6561[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[58]), .B1(integrator4_adj_6561[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17413), .COUT(n17414), .S0(n120_adj_6488), 
          .S1(n117_adj_6487));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_39 (.A0(\phase_increment[0] [38]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [39]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17617), .COUT(n17618), .S0(phase_increment_1__63__N_20[38]), 
          .S1(phase_increment_1__63__N_20[39]));
    defparam _add_1_3813_add_4_39.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_37 (.A0(\phase_increment[0] [36]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [37]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17616), .COUT(n17617), .S0(phase_increment_1__63__N_20[36]), 
          .S1(phase_increment_1__63__N_20[37]));
    defparam _add_1_3813_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_3813_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_22 (.A0(integrator5_adj_6562[55]), .B0(integrator4_adj_6561[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[56]), .B1(integrator4_adj_6561[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17412), .COUT(n17413), .S0(n126_adj_6490), 
          .S1(n123_adj_6489));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_10 (.A0(integrator3_adj_6560[43]), .B0(integrator2_adj_6559[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[44]), .B1(integrator2_adj_6559[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17450), .COUT(n17451), .S0(n162_adj_6416), 
          .S1(n159_adj_6415));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3618_add_4_20 (.A0(integrator5_adj_6562[53]), .B0(integrator4_adj_6561[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[54]), .B1(integrator4_adj_6561[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17411), .COUT(n17412), .S0(n132_adj_6492), 
          .S1(n129_adj_6491));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_8 (.A0(integrator3_adj_6560[41]), .B0(integrator2_adj_6559[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[42]), .B1(integrator2_adj_6559[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17449), .COUT(n17450), .S0(n168_adj_6418), 
          .S1(n165_adj_6417));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_8.INJECT1_1 = "NO";
    \CIC(REGISTER_WIDTH=72,DECIMATION_RATIO=4096)  cic_sine_inst (.comb_d7({comb_d7}), 
            .n14(n14_adj_5396), .comb_d6({comb_d6}), .n20(n20_adj_5366), 
            .integrator_d_tmp({integrator_d_tmp}), .clk_80mhz(clk_80mhz), 
            .integrator_tmp({integrator_tmp}), .\cic_gain[0] (cic_gain[0]), 
            .integrator2({integrator2}), .integrator2_71__N_1032({integrator2_71__N_1032}), 
            .\cic_gain[1] (cic_gain[1]), .integrator3({integrator3}), .integrator3_71__N_1104({integrator3_71__N_1104}), 
            .integrator4({integrator4}), .integrator4_71__N_1176({integrator4_71__N_1176}), 
            .integrator5({integrator5}), .integrator5_71__N_1248({integrator5_71__N_1248}), 
            .comb6({comb6}), .comb6_71__N_1993({comb6_71__N_1993}), .cic_sine_clk(cic_sine_clk), 
            .n27(n27_adj_5373), .comb7({comb7}), .comb7_71__N_2065({comb7_71__N_2065}), 
            .comb8({comb8}), .comb8_71__N_2137({comb8_71__N_2137}), .comb_d8({comb_d8}), 
            .comb9({comb9}), .comb9_71__N_2209({comb9_71__N_2209}), .comb_d9({comb_d9}), 
            .integrator1({integrator1}), .integrator1_71__N_960({integrator1_71__N_960}), 
            .count({count}), .n26(n26_adj_5372), .n35(n35_adj_5381), .n34(n34_adj_5380), 
            .n17(n17_adj_5399), .n16(n16_adj_5398), .n29(n29_adj_5375), 
            .n28(n28_adj_5374), .n37(n37_adj_5383), .n9(n9_adj_5391), 
            .\comb10[67] (comb10_adj_6571[67]), .\comb10[69] (comb10_adj_6571[69]), 
            .n8(n8_adj_5390), .n36(n36_adj_5382), .n23(n23_adj_5369), 
            .\comb10[68] (comb10_adj_6571[68]), .\comb10[70] (comb10_adj_6571[70]), 
            .n22(n22_adj_5368), .n31(n31_adj_5377), .n30(n30_adj_5376), 
            .n25(n25_adj_5371), .n24(n24_adj_5370), .n33(n33_adj_5379), 
            .n32(n32_adj_5378), .n21(n21_adj_5403), .n20_adj_115(n20_adj_5402), 
            .n19(n19_adj_5401), .n18(n18_adj_5400), .n25_adj_116(n25_adj_5407), 
            .n24_adj_117(n24_adj_5406), .n23_adj_118(n23_adj_5405), .n22_adj_119(n22_adj_5404), 
            .n3(n3_adj_5385), .n31_adj_120(n31_adj_5413), .n30_adj_121(n30_adj_5412), 
            .n29_adj_122(n29_adj_5411), .n28_adj_123(n28_adj_5410), .n27_adj_124(n27_adj_5409), 
            .n26_adj_125(n26_adj_5408), .n35_adj_126(n35_adj_5417), .n34_adj_127(n34_adj_5416), 
            .n2(n2_adj_5384), .n37_adj_128(n37_adj_5419), .n36_adj_129(n36_adj_5418), 
            .n5(n5_adj_5387), .n7(n7_adj_5425), .n4(n4_adj_5386), .n6(n6_adj_5424), 
            .n5_adj_130(n5_adj_5423), .n4_adj_131(n4_adj_5422), .n3_adj_132(n3_adj_5421), 
            .n2_adj_133(n2_adj_5420), .n17_adj_134(n17_adj_5435), .n16_adj_135(n16_adj_5434), 
            .n15(n15_adj_5433), .n14_adj_136(n14_adj_5432), .n11(n11_adj_5429), 
            .n10(n10_adj_5428), .n13(n13_adj_5431), .n12(n12_adj_5430), 
            .n25_adj_137(n25_adj_5443), .n24_adj_138(n24_adj_5442), .n62(n62), 
            .\comb10[60] (comb10_adj_6571[60]), .n23_adj_139(n23_adj_5441), 
            .n22_adj_140(n22_adj_5440), .n21_adj_141(n21_adj_5439), .n20_adj_142(n20_adj_5438), 
            .n33_adj_143(n33_adj_5451), .n32_adj_144(n32_adj_5450), .n31_adj_145(n31_adj_5449), 
            .n30_adj_146(n30_adj_5448), .n29_adj_147(n29_adj_5447), .n28_adj_148(n28_adj_5446), 
            .n37_adj_149(n37_adj_5455), .n36_adj_150(n36_adj_5454), .n3_adj_151(n3), 
            .n2_adj_152(n2), .n5_adj_153(n5), .n4_adj_154(n4), .n68(n68), 
            .\comb10[66] (comb10_adj_6571[66]), .n67_adj_228({n28, n31, 
            n34, n37_adj_5270, n40, n43, n46, n49, n52, n55, 
            n58, n61}), .n76(n76_adj_6527), .n78(n78_adj_5825), .cout(cout_adj_6511), 
            .n79(n79_adj_6528), .n81(n81_adj_5826), .n82(n82_adj_6529), 
            .n84(n84_adj_5827), .n85(n85_adj_6530), .n87(n87_adj_5828), 
            .n88(n88_adj_6531), .n90(n90_adj_5829), .n91(n91_adj_6532), 
            .n93(n93_adj_5830), .led_0_2(led_0_2), .n94(n94_adj_6533), 
            .n96(n96_adj_5831), .n97(n97_adj_6534), .n99(n99_adj_5832), 
            .n100(n100_adj_6535), .n102(n102_adj_5833), .n103(n103_adj_6536), 
            .n105(n105_adj_5834), .n67(n67), .\comb10[65] (comb10_adj_6571[65]), 
            .n106(n106_adj_6537), .n108(n108_adj_5835), .n109(n109_adj_6538), 
            .n111(n111_adj_5836), .n66(n66_adj_5290), .\comb10[64] (comb10_adj_6571[64]), 
            .n112(n112_adj_6539), .n114(n114_adj_5837), .n115(n115_adj_6540), 
            .n117(n117_adj_5838), .n118(n118_adj_6541), .n120(n120_adj_5839), 
            .n64(n64), .\comb10[62] (comb10_adj_6571[62]), .n19_adj_159(n19_adj_5437), 
            .n63(n63_adj_5289), .\comb10[61] (comb10_adj_6571[61]), .n65(n65), 
            .\comb10[63] (comb10_adj_6571[63]), .n7_adj_160(n7), .n6_adj_161(n6), 
            .n13_adj_162(n13), .n12_adj_163(n12), .n21_adj_164(n21), .n20_adj_165(n20), 
            .n15_adj_166(n15), .n14_adj_167(n14), .n23_adj_168(n23), .n22_adj_169(n22), 
            .n9_adj_170(n9), .n8_adj_171(n8), .n17_adj_172(n17), .n16_adj_173(n16), 
            .n25_adj_174(n25), .n24_adj_175(n24), .n11_adj_176(n11), .n10_adj_177(n10), 
            .n19_adj_178(n19), .n18_adj_179(n18), .n27_adj_180(n27), .n26_adj_181(n26), 
            .n33_adj_182(n33), .n32_adj_183(n32), .n35_adj_184(n35), .n34_adj_185(n34_adj_5272), 
            .n29_adj_186(n29), .n28_adj_187(n28_adj_5274), .n37_adj_188(n37), 
            .n36_adj_189(n36), .n3_adj_190(n3_adj_5304), .n2_adj_191(n2_adj_5354), 
            .n31_adj_192(n31_adj_5273), .n30_adj_193(n30), .n5_adj_194(n5_adj_5300), 
            .n4_adj_195(n4_adj_5301), .n11_adj_196(n11_adj_5357), .n10_adj_197(n10_adj_5356), 
            .n17_adj_198(n17_adj_5363), .n16_adj_199(n16_adj_5362), .n13_adj_200(n13_adj_5359), 
            .n12_adj_201(n12_adj_5358), .n7_adj_202(n7_adj_5294), .n6_adj_203(n6_adj_5298), 
            .n15_adj_204(n15_adj_5361), .n14_adj_205(n14_adj_5360), .n61_adj_206(n61_adj_5288), 
            .\comb10[59] (comb10_adj_6571[59]), .n19_adj_207(n19_adj_5365), 
            .n18_adj_208(n18_adj_5364), .n9_adj_209(n9_adj_5355), .n8_adj_210(n8_adj_5286), 
            .n21_adj_211(n21_adj_5367), .led_0_1(led_0_1), .led_0_0(led_0_0), 
            .\cic_sine_out[5] (cic_sine_out[5]), .n7_adj_212(n7_adj_5389), 
            .n6_adj_213(n6_adj_5388), .n13_adj_214(n13_adj_5395), .n12_adj_215(n12_adj_5394), 
            .n15_adj_216(n15_adj_5397), .\cic_sine_out[4] (cic_sine_out[4]), 
            .\cic_sine_out[3] (cic_sine_out[3]), .\cic_sine_out[2] (cic_sine_out[2]), 
            .\comb10[71] (comb10_adj_6571[71]), .\cic_cosine_out[11] (cic_cosine_out[11]), 
            .n70(n70), .\cic_cosine_out[9] (cic_cosine_out[9]), .\cic_cosine_out[8] (cic_cosine_out[8]), 
            .\cic_cosine_out[7] (cic_cosine_out[7]), .\cic_cosine_out[6] (cic_cosine_out[6]), 
            .\cic_cosine_out[5] (cic_cosine_out[5]), .\cic_cosine_out[4] (cic_cosine_out[4]), 
            .\cic_cosine_out[3] (cic_cosine_out[3]), .\cic_cosine_out[2] (cic_cosine_out[2]), 
            .led_0_5(led_0_5), .led_0_3(led_0_3), .n18_adj_217(n18_adj_5436), 
            .n11_adj_218(n11_adj_5393), .n10_adj_219(n10_adj_5392), .n33_adj_220(n33_adj_5415), 
            .n32_adj_221(n32_adj_5414), .n9_adj_222(n9_adj_5427), .n8_adj_223(n8_adj_5426), 
            .\cic_cosine_out[10] (cic_cosine_out[10]), .led_0_4(led_0_4), 
            .\cic_sine_out[1] (cic_sine_out[1]), .\cic_sine_out[0] (cic_sine_out[0]), 
            .n27_adj_224(n27_adj_5445), .n26_adj_225(n26_adj_5444), .n35_adj_226(n35_adj_5453), 
            .n34_adj_227(n34_adj_5452)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(190[7] 196[6])
    CCU2C _add_1_3618_add_4_18 (.A0(integrator5_adj_6562[51]), .B0(integrator4_adj_6561[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[52]), .B1(integrator4_adj_6561[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17410), .COUT(n17411), .S0(n138_adj_6494), 
          .S1(n135_adj_6493));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_10 (.A0(integrator4_adj_6561[43]), .B0(integrator3_adj_6560[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[44]), .B1(integrator3_adj_6560[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17432), .COUT(n17433), .S0(n162_adj_6452), 
          .S1(n159_adj_6451));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_6 (.A0(integrator3_adj_6560[39]), .B0(integrator2_adj_6559[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[40]), .B1(integrator2_adj_6559[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17448), .COUT(n17449), .S0(n174_adj_6420), 
          .S1(n171_adj_6419));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_6.INJECT1_1 = "NO";
    PFUMX mux_2474_i1 (.BLUT(n4065), .ALUT(n4050), .C0(rx_byte[2]), .Z(n4073));
    CCU2C _add_1_3618_add_4_16 (.A0(integrator5_adj_6562[49]), .B0(integrator4_adj_6561[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6562[50]), .B1(integrator4_adj_6561[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17409), .COUT(n17410), .S0(n144_adj_6496), 
          .S1(n141_adj_6495));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(77[20:45])
    defparam _add_1_3618_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_3618_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_3618_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3618_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_8 (.A0(integrator4_adj_6561[41]), .B0(integrator3_adj_6560[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[42]), .B1(integrator3_adj_6560[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17431), .COUT(n17432), .S0(n168_adj_6454), 
          .S1(n165_adj_6453));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_4 (.A0(integrator3_adj_6560[37]), .B0(integrator2_adj_6559[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6560[38]), .B1(integrator2_adj_6559[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17447), .COUT(n17448), .S0(n180_adj_6422), 
          .S1(n177_adj_6421));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3609_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_6 (.A0(integrator4_adj_6561[39]), .B0(integrator3_adj_6560[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[40]), .B1(integrator3_adj_6560[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17430), .COUT(n17431), .S0(n174_adj_6456), 
          .S1(n171_adj_6455));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3609_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator3_adj_6560[36]), .B1(integrator2_adj_6559[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n17447), .S1(n183_adj_6423));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(75[20:45])
    defparam _add_1_3609_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3609_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3609_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3609_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3813_add_4_35 (.A0(\phase_increment[0] [34]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\phase_increment[0] [35]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17615), .COUT(n17616), .S0(phase_increment_1__63__N_20[34]), 
          .S1(phase_increment_1__63__N_20[35]));
    defparam _add_1_3813_add_4_35.INIT0 = 16'h555f;
    defparam _add_1_3813_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_3813_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3813_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_4 (.A0(integrator4_adj_6561[37]), .B0(integrator3_adj_6560[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[38]), .B1(integrator3_adj_6560[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17429), .COUT(n17430), .S0(n180_adj_6458), 
          .S1(n177_adj_6457));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_38 (.A0(integrator4_adj_6561[71]), .B0(integrator3_adj_6560[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17446), .S0(n78_adj_6424));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3612_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator4_adj_6561[36]), .B1(integrator3_adj_6560[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n17429), .S1(n183_adj_6459));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3612_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_36 (.A0(integrator4_adj_6561[69]), .B0(integrator3_adj_6560[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[70]), .B1(integrator3_adj_6560[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17445), .COUT(n17446), .S0(n84_adj_6426), 
          .S1(n81_adj_6425));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3615_add_4_16 (.A0(amdemod_out_d_11__N_2399[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2399[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17427), .S1(n36_adj_6460));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3615_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_3615_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3615_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3615_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_34 (.A0(integrator4_adj_6561[67]), .B0(integrator3_adj_6560[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[68]), .B1(integrator3_adj_6560[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17444), .COUT(n17445), .S0(n90_adj_6428), 
          .S1(n87_adj_6427));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3615_add_4_14 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2399[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2399[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17426), .COUT(n17427), 
          .S0(n45_adj_6462), .S1(n42_adj_6461));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3615_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_3615_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_3615_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3615_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3612_add_4_32 (.A0(integrator4_adj_6561[65]), .B0(integrator3_adj_6560[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6561[66]), .B1(integrator3_adj_6560[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17443), .COUT(n17444), .S0(n96_adj_6430), 
          .S1(n93_adj_6429));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(76[20:45])
    defparam _add_1_3612_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3612_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3612_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3612_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_26 (.A0(integrator2[59]), .B0(integrator1[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[60]), .B1(integrator1[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17841), .COUT(n17842), .S0(n114_adj_5333), 
          .S1(n111_adj_5339));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_28 (.A0(integrator2[61]), .B0(integrator1[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[62]), .B1(integrator1[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17842), .COUT(n17843), .S0(n108_adj_5313), 
          .S1(n105_adj_5319));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_30 (.A0(integrator2[63]), .B0(integrator1[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[64]), .B1(integrator1[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17843), .COUT(n17844), .S0(n102_adj_5335), 
          .S1(n99_adj_5340));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_32 (.A0(integrator2[65]), .B0(integrator1[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[66]), .B1(integrator1[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17844), .COUT(n17845), .S0(n96_adj_5334), 
          .S1(n93_adj_5337));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_34 (.A0(integrator2[67]), .B0(integrator1[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[68]), .B1(integrator1[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17845), .COUT(n17846), .S0(n90_adj_5331), 
          .S1(n87_adj_5336));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_36 (.A0(integrator2[69]), .B0(integrator1[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[70]), .B1(integrator1[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17846), .COUT(n17847), .S0(n84_adj_5322), 
          .S1(n81_adj_5323));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_3525_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_3525_add_4_38 (.A0(integrator2[71]), .B0(integrator1[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17847), .S0(n78_adj_5330));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3525_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_3525_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_3525_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_3525_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[18]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17848), .S1(amdemod_out_d_11__N_2370[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3759_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3759_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3759_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_3 (.A0(square_sum[19]), .B0(square_sum[25]), 
          .C0(n30_adj_6282), .D0(n13890), .A1(amdemod_out_d_11__N_2363), 
          .B1(n48_adj_6288), .C1(square_sum[25]), .D1(n13815), .CIN(n17848), 
          .COUT(n17849), .S0(amdemod_out_d_11__N_2370[1]), .S1(amdemod_out_d_11__N_2370[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3759_add_4_3.INIT0 = 16'h596a;
    defparam _add_1_3759_add_4_3.INIT1 = 16'h9a95;
    defparam _add_1_3759_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_5 (.A0(square_sum[25]), .B0(n19824), .C0(n45_adj_6287), 
          .D0(n13876), .A1(square_sum[25]), .B1(amdemod_out_d_11__N_2516), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17849), .COUT(n17850), .S0(amdemod_out_d_11__N_2370[3]), 
          .S1(amdemod_out_d_11__N_2370[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3759_add_4_5.INIT0 = 16'h1b4e;
    defparam _add_1_3759_add_4_5.INIT1 = 16'h666a;
    defparam _add_1_3759_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_7 (.A0(amdemod_out_d_11__N_2513), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2510), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17850), .COUT(n17851), .S0(amdemod_out_d_11__N_2370[5]), 
          .S1(amdemod_out_d_11__N_2370[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3759_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_9 (.A0(amdemod_out_d_11__N_2507), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2504), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17851), .COUT(n17852), .S0(amdemod_out_d_11__N_2370[7]), 
          .S1(amdemod_out_d_11__N_2370[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3759_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_11 (.A0(amdemod_out_d_11__N_2501), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2363), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17852), .COUT(n17853), .S0(amdemod_out_d_11__N_2370[9]), 
          .S1(amdemod_out_d_11__N_2370[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3759_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_13 (.A0(amdemod_out_d_11__N_2363), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17853), .S0(amdemod_out_d_11__N_2370[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3759_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_3759_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3756_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17854), .S1(n76_adj_6170));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3756_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3756_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3756_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3756_add_4_3 (.A0(square_sum[13]), .B0(amdemod_out_d_11__N_2380[14]), 
          .C0(n19815), .D0(amdemod_out_d_11__N_2379[14]), .A1(n19814), 
          .B1(amdemod_out_d_11__N_2379[0]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17854), .COUT(n17855), .S0(n73_adj_6169), .S1(n70_adj_6168));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3756_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_3756_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3756_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3756_add_4_5 (.A0(n19815), .B0(amdemod_out_d_11__N_2379[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n19816), .B1(amdemod_out_d_11__N_2379[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17855), .COUT(n17856), .S0(n67_adj_6167), 
          .S1(n64_adj_6166));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3756_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3756_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_3756_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3756_add_4_7 (.A0(amdemod_out_d_11__N_2363), .B0(amdemod_out_d_11__N_2379[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2379[4]), .D1(VCC_net), .CIN(n17856), 
          .COUT(n17857), .S0(n61_adj_6165), .S1(n58_adj_6164));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3756_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_3756_add_4_7.INIT1 = 16'h1e1e;
    defparam _add_1_3756_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3756_add_4_9 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2379[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2379[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17857), .COUT(n17858), 
          .S0(n55_adj_6163), .S1(n52_adj_6162));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3756_add_4_9.INIT0 = 16'h666a;
    defparam _add_1_3756_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_3756_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3756_add_4_11 (.A0(amdemod_out_d_11__N_2379[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2379[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17858), .COUT(n17859), 
          .S0(n49_adj_6161), .S1(n46_adj_6160));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3756_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3756_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3756_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3756_add_4_13 (.A0(amdemod_out_d_11__N_2379[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2379[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17859), .COUT(n17860), 
          .S0(n43_adj_6159), .S1(n40_adj_6158));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3756_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3756_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3756_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3756_add_4_15 (.A0(amdemod_out_d_11__N_2379[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2379[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17860), .S1(n34_adj_6157));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3756_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3756_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3756_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5318), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17865));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3753_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_3753_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_3 (.A0(integrator1[36]), .B0(cout_adj_5318), 
          .C0(n183_adj_5324), .D0(integrator2[36]), .A1(integrator1[37]), 
          .B1(cout_adj_5318), .C1(n180_adj_5325), .D1(integrator2[37]), 
          .CIN(n17865), .COUT(n17866), .S0(integrator2_71__N_1032[36]), 
          .S1(integrator2_71__N_1032[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_5 (.A0(integrator1[38]), .B0(cout_adj_5318), 
          .C0(n177_adj_5351), .D0(integrator2[38]), .A1(integrator1[39]), 
          .B1(cout_adj_5318), .C1(n174_adj_5303), .D1(integrator2[39]), 
          .CIN(n17866), .COUT(n17867), .S0(integrator2_71__N_1032[38]), 
          .S1(integrator2_71__N_1032[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_7 (.A0(integrator1[40]), .B0(cout_adj_5318), 
          .C0(n171_adj_5306), .D0(integrator2[40]), .A1(integrator1[41]), 
          .B1(cout_adj_5318), .C1(n168_adj_5350), .D1(integrator2[41]), 
          .CIN(n17867), .COUT(n17868), .S0(integrator2_71__N_1032[40]), 
          .S1(integrator2_71__N_1032[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_9 (.A0(integrator1[42]), .B0(cout_adj_5318), 
          .C0(n165_adj_5347), .D0(integrator2[42]), .A1(integrator1[43]), 
          .B1(cout_adj_5318), .C1(n162_adj_5309), .D1(integrator2[43]), 
          .CIN(n17868), .COUT(n17869), .S0(integrator2_71__N_1032[42]), 
          .S1(integrator2_71__N_1032[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_11 (.A0(integrator1[44]), .B0(cout_adj_5318), 
          .C0(n159_adj_5307), .D0(integrator2[44]), .A1(integrator1[45]), 
          .B1(cout_adj_5318), .C1(n156_adj_5352), .D1(integrator2[45]), 
          .CIN(n17869), .COUT(n17870), .S0(integrator2_71__N_1032[44]), 
          .S1(integrator2_71__N_1032[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_13 (.A0(integrator1[46]), .B0(cout_adj_5318), 
          .C0(n153_adj_5349), .D0(integrator2[46]), .A1(integrator1[47]), 
          .B1(cout_adj_5318), .C1(n150_adj_5346), .D1(integrator2[47]), 
          .CIN(n17870), .COUT(n17871), .S0(integrator2_71__N_1032[46]), 
          .S1(integrator2_71__N_1032[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_15 (.A0(integrator1[48]), .B0(cout_adj_5318), 
          .C0(n147_adj_5344), .D0(integrator2[48]), .A1(integrator1[49]), 
          .B1(cout_adj_5318), .C1(n144_adj_5348), .D1(integrator2[49]), 
          .CIN(n17871), .COUT(n17872), .S0(integrator2_71__N_1032[48]), 
          .S1(integrator2_71__N_1032[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_17 (.A0(integrator1[50]), .B0(cout_adj_5318), 
          .C0(n141), .D0(integrator2[50]), .A1(integrator1[51]), .B1(cout_adj_5318), 
          .C1(n138_adj_5345), .D1(integrator2[51]), .CIN(n17872), .COUT(n17873), 
          .S0(integrator2_71__N_1032[50]), .S1(integrator2_71__N_1032[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_19 (.A0(integrator1[52]), .B0(cout_adj_5318), 
          .C0(n135_adj_5343), .D0(integrator2[52]), .A1(integrator1[53]), 
          .B1(cout_adj_5318), .C1(n132_adj_5311), .D1(integrator2[53]), 
          .CIN(n17873), .COUT(n17874), .S0(integrator2_71__N_1032[52]), 
          .S1(integrator2_71__N_1032[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_21 (.A0(integrator1[54]), .B0(cout_adj_5318), 
          .C0(n129_adj_5312), .D0(integrator2[54]), .A1(integrator1[55]), 
          .B1(cout_adj_5318), .C1(n126_adj_5338), .D1(integrator2[55]), 
          .CIN(n17874), .COUT(n17875), .S0(integrator2_71__N_1032[54]), 
          .S1(integrator2_71__N_1032[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_23 (.A0(integrator1[56]), .B0(cout_adj_5318), 
          .C0(n123_adj_5342), .D0(integrator2[56]), .A1(integrator1[57]), 
          .B1(cout_adj_5318), .C1(n120_adj_5315), .D1(integrator2[57]), 
          .CIN(n17875), .COUT(n17876), .S0(integrator2_71__N_1032[56]), 
          .S1(integrator2_71__N_1032[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_25 (.A0(integrator1[58]), .B0(cout_adj_5318), 
          .C0(n117_adj_5316), .D0(integrator2[58]), .A1(integrator1[59]), 
          .B1(cout_adj_5318), .C1(n114_adj_5333), .D1(integrator2[59]), 
          .CIN(n17876), .COUT(n17877), .S0(integrator2_71__N_1032[58]), 
          .S1(integrator2_71__N_1032[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_27 (.A0(integrator1[60]), .B0(cout_adj_5318), 
          .C0(n111_adj_5339), .D0(integrator2[60]), .A1(integrator1[61]), 
          .B1(cout_adj_5318), .C1(n108_adj_5313), .D1(integrator2[61]), 
          .CIN(n17877), .COUT(n17878), .S0(integrator2_71__N_1032[60]), 
          .S1(integrator2_71__N_1032[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_29 (.A0(integrator1[62]), .B0(cout_adj_5318), 
          .C0(n105_adj_5319), .D0(integrator2[62]), .A1(integrator1[63]), 
          .B1(cout_adj_5318), .C1(n102_adj_5335), .D1(integrator2[63]), 
          .CIN(n17878), .COUT(n17879), .S0(integrator2_71__N_1032[62]), 
          .S1(integrator2_71__N_1032[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_31 (.A0(integrator1[64]), .B0(cout_adj_5318), 
          .C0(n99_adj_5340), .D0(integrator2[64]), .A1(integrator1[65]), 
          .B1(cout_adj_5318), .C1(n96_adj_5334), .D1(integrator2[65]), 
          .CIN(n17879), .COUT(n17880), .S0(integrator2_71__N_1032[64]), 
          .S1(integrator2_71__N_1032[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_33 (.A0(integrator1[66]), .B0(cout_adj_5318), 
          .C0(n93_adj_5337), .D0(integrator2[66]), .A1(integrator1[67]), 
          .B1(cout_adj_5318), .C1(n90_adj_5331), .D1(integrator2[67]), 
          .CIN(n17880), .COUT(n17881), .S0(integrator2_71__N_1032[66]), 
          .S1(integrator2_71__N_1032[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_35 (.A0(integrator1[68]), .B0(cout_adj_5318), 
          .C0(n87_adj_5336), .D0(integrator2[68]), .A1(integrator1[69]), 
          .B1(cout_adj_5318), .C1(n84_adj_5322), .D1(integrator2[69]), 
          .CIN(n17881), .COUT(n17882), .S0(integrator2_71__N_1032[68]), 
          .S1(integrator2_71__N_1032[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_37 (.A0(integrator1[70]), .B0(cout_adj_5318), 
          .C0(n81_adj_5323), .D0(integrator2[70]), .A1(integrator1[71]), 
          .B1(cout_adj_5318), .C1(n78_adj_5330), .D1(integrator2[71]), 
          .CIN(n17882), .S0(integrator2_71__N_1032[70]), .S1(integrator2_71__N_1032[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(74[20:45])
    defparam _add_1_3753_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_3753_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_3753_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17884), .S1(n76_adj_6156));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3750_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3750_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3750_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_3 (.A0(square_sum[13]), .B0(amdemod_out_d_11__N_2380[14]), 
          .C0(n19815), .D0(amdemod_out_d_11__N_2379[14]), .A1(n19814), 
          .B1(amdemod_out_d_11__N_2380[0]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17884), .COUT(n17885), .S0(n73_adj_6155), .S1(n70_adj_6154));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3750_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_3750_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_3750_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_5 (.A0(n19815), .B0(amdemod_out_d_11__N_2380[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n19816), .B1(amdemod_out_d_11__N_2380[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17885), .COUT(n17886), .S0(n67_adj_6153), 
          .S1(n64_adj_6152));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3750_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_3750_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_3750_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_7 (.A0(amdemod_out_d_11__N_2363), .B0(amdemod_out_d_11__N_2380[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2380[4]), .D1(VCC_net), .CIN(n17886), 
          .COUT(n17887), .S0(n61_adj_6151), .S1(n58_adj_6150));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3750_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_3750_add_4_7.INIT1 = 16'h1e1e;
    defparam _add_1_3750_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_9 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2380[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2380[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17887), .COUT(n17888), 
          .S0(n55_adj_6149), .S1(n52_adj_6148));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3750_add_4_9.INIT0 = 16'h666a;
    defparam _add_1_3750_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_3750_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_11 (.A0(amdemod_out_d_11__N_2380[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2380[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17888), .COUT(n17889), 
          .S0(n49_adj_6147), .S1(n46_adj_6146));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3750_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3750_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3750_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_13 (.A0(amdemod_out_d_11__N_2380[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2380[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17889), .COUT(n17890), 
          .S0(n43_adj_6145), .S1(n40_adj_6144));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3750_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3750_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3750_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_15 (.A0(amdemod_out_d_11__N_2380[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2380[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17890), .S1(n34_adj_6143));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam _add_1_3750_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3750_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3750_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3558_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_adj_6572[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17894), .S1(n61_adj_6142));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3558_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3558_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3558_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3558_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3558_add_4_3 (.A0(count_adj_6572[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_6572[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17894), .COUT(n17895), .S0(n58_adj_6141), 
          .S1(n55_adj_6140));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3558_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_3558_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_3558_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3558_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3558_add_4_5 (.A0(count_adj_6572[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_6572[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17895), .COUT(n17896), .S0(n52_adj_6139), 
          .S1(n49_adj_6138));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3558_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_3558_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_3558_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3558_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3558_add_4_7 (.A0(count_adj_6572[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_6572[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17896), .COUT(n17897), .S0(n46_adj_6137), 
          .S1(n43_adj_6136));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3558_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_3558_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_3558_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3558_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3558_add_4_9 (.A0(count_adj_6572[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_6572[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17897), .COUT(n17898), .S0(n40_adj_6135), 
          .S1(n37_adj_6134));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3558_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_3558_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_3558_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3558_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3558_add_4_11 (.A0(count_adj_6572[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_6572[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17898), .COUT(n17899), .S0(n34_adj_6133), 
          .S1(n31_adj_6132));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3558_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3558_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3558_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3558_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3558_add_4_13 (.A0(count_adj_6572[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17899), .S0(n28_adj_6131));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(93[25:34])
    defparam _add_1_3558_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3558_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_3558_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3558_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3555_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17900));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3555_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_3555_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_3555_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_3555_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_3555_add_4_4 (.A0(n19808), .B0(square_sum[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_out_d_11__N_2409[0]), .B1(amdemod_out_d_11__N_2410[14]), 
          .C1(n19809), .D1(amdemod_out_d_11__N_2409[14]), .CIN(n17900), 
          .COUT(n17901));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3555_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_3555_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_3555_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_3555_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_3555_add_4_6 (.A0(n19809), .B0(amdemod_out_d_11__N_2409[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2409[2]), 
          .B1(amdemod_out_d_11__N_2400[14]), .C1(n19811), .D1(amdemod_out_d_11__N_2399[14]), 
          .CIN(n17901), .COUT(n17902));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3555_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_3555_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_3555_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_3555_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_3555_add_4_8 (.A0(n19811), .B0(amdemod_out_d_11__N_2409[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2409[4]), 
          .B1(amdemod_out_d_11__N_2390[14]), .C1(n19813), .D1(amdemod_out_d_11__N_2389[14]), 
          .CIN(n17902), .COUT(n17903));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3555_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_3555_add_4_8.INIT1 = 16'h656a;
    defparam _add_1_3555_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_3555_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_3555_add_4_10 (.A0(n19813), .B0(amdemod_out_d_11__N_2409[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2409[6]), 
          .B1(amdemod_out_d_11__N_2380[14]), .C1(n19815), .D1(amdemod_out_d_11__N_2379[14]), 
          .CIN(n17903), .COUT(n17904));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3555_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_3555_add_4_10.INIT1 = 16'h656a;
    defparam _add_1_3555_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_3555_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_3555_add_4_12 (.A0(n19815), .B0(amdemod_out_d_11__N_2409[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2409[8]), 
          .B1(amdemod_out_d_11__N_2370[11]), .C1(amdemod_out_d_11__N_2363), 
          .D1(amdemod_out_d_11__N_2369[11]), .CIN(n17904), .COUT(n17905));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3555_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_3555_add_4_12.INIT1 = 16'h656a;
    defparam _add_1_3555_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_3555_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_3555_add_4_14 (.A0(amdemod_out_d_11__N_2409[9]), .B0(square_sum[25]), 
          .C0(n30_adj_6282), .D0(n13890), .A1(square_sum[25]), .B1(n19824), 
          .C1(amdemod_out_d_11__N_2409[10]), .D1(VCC_net), .CIN(n17905), 
          .COUT(n17906));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3555_add_4_14.INIT0 = 16'h596a;
    defparam _add_1_3555_add_4_14.INIT1 = 16'he1e1;
    defparam _add_1_3555_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_3555_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_3555_add_4_16 (.A0(square_sum[25]), .B0(amdemod_out_d_11__N_2409[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_out_d_11__N_2409[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n17906), .S1(n36_adj_6130));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3555_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_3555_add_4_16.INIT1 = 16'h555f;
    defparam _add_1_3555_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_3555_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_3810_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[20]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17908), .S1(n48_adj_6288));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3810_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3810_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3810_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3810_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3810_add_4_3 (.A0(square_sum[25]), .B0(n19824), .C0(square_sum[21]), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(n19824), .C1(square_sum[22]), 
          .D1(VCC_net), .CIN(n17908), .COUT(n17909), .S0(n45_adj_6287), 
          .S1(n42_adj_6286));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3810_add_4_3.INIT0 = 16'h1e1e;
    defparam _add_1_3810_add_4_3.INIT1 = 16'h1e11;
    defparam _add_1_3810_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3810_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3810_add_4_5 (.A0(square_sum[25]), .B0(n4_adj_6510), .C0(amdemod_out_d_11__N_2358[5]), 
          .D0(VCC_net), .A1(square_sum[22]), .B1(n13821), .C1(square_sum[25]), 
          .D1(square_sum[23]), .CIN(n17909), .COUT(n17910), .S0(n39_adj_6285), 
          .S1(n36_adj_6284));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3810_add_4_5.INIT0 = 16'h9696;
    defparam _add_1_3810_add_4_5.INIT1 = 16'h135f;
    defparam _add_1_3810_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3810_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3810_add_4_7 (.A0(square_sum[25]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17910), .S0(n33_adj_6283), .S1(n30_adj_6282));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam _add_1_3810_add_4_7.INIT0 = 16'haaaf;
    defparam _add_1_3810_add_4_7.INIT1 = 16'haaaf;
    defparam _add_1_3810_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3810_add_4_7.INJECT1_1 = "NO";
    CCU2C add_5422_1 (.A0(square_sum[0]), .B0(GND_net), .C0(GND_net), 
          .D0(square_sum[0]), .A1(square_sum[1]), .B1(amdemod_out_d_11__N_2410[14]), 
          .C1(n19809), .D1(amdemod_out_d_11__N_2409[14]), .COUT(n17912));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5422_1.INIT0 = 16'h000A;
    defparam add_5422_1.INIT1 = 16'h656a;
    defparam add_5422_1.INJECT1_0 = "NO";
    defparam add_5422_1.INJECT1_1 = "NO";
    CCU2C add_5422_3 (.A0(n19808), .B0(amdemod_out_d_11__N_2410[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19809), .B1(amdemod_out_d_11__N_2410[1]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17912), .COUT(n17913));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5422_3.INIT0 = 16'h9995;
    defparam add_5422_3.INIT1 = 16'h9995;
    defparam add_5422_3.INJECT1_0 = "NO";
    defparam add_5422_3.INJECT1_1 = "NO";
    CCU2C add_5422_5 (.A0(n19810), .B0(amdemod_out_d_11__N_2410[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19811), .B1(amdemod_out_d_11__N_2410[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17913), .COUT(n17914));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5422_5.INIT0 = 16'h9995;
    defparam add_5422_5.INIT1 = 16'h9995;
    defparam add_5422_5.INJECT1_0 = "NO";
    defparam add_5422_5.INJECT1_1 = "NO";
    CCU2C add_5422_7 (.A0(n19812), .B0(amdemod_out_d_11__N_2410[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19813), .B1(amdemod_out_d_11__N_2410[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17914), .COUT(n17915));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5422_7.INIT0 = 16'h9995;
    defparam add_5422_7.INIT1 = 16'h9995;
    defparam add_5422_7.INJECT1_0 = "NO";
    defparam add_5422_7.INJECT1_1 = "NO";
    CCU2C add_5422_9 (.A0(n19814), .B0(amdemod_out_d_11__N_2410[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(n19815), .B1(amdemod_out_d_11__N_2410[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17915), .COUT(n17916));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5422_9.INIT0 = 16'h9995;
    defparam add_5422_9.INIT1 = 16'h9995;
    defparam add_5422_9.INJECT1_0 = "NO";
    defparam add_5422_9.INJECT1_1 = "NO";
    CCU2C add_5422_11 (.A0(n19816), .B0(amdemod_out_d_11__N_2410[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_out_d_11__N_2363), .B1(amdemod_out_d_11__N_2410[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17916), .COUT(n17917));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5422_11.INIT0 = 16'h9995;
    defparam add_5422_11.INIT1 = 16'h9995;
    defparam add_5422_11.INJECT1_0 = "NO";
    defparam add_5422_11.INJECT1_1 = "NO";
    CCU2C add_5422_13 (.A0(square_sum[25]), .B0(n19824), .C0(amdemod_out_d_11__N_2410[10]), 
          .D0(VCC_net), .A1(square_sum[25]), .B1(amdemod_out_d_11__N_2410[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17917), .COUT(n17918));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5422_13.INIT0 = 16'h1e1e;
    defparam add_5422_13.INIT1 = 16'h666a;
    defparam add_5422_13.INJECT1_0 = "NO";
    defparam add_5422_13.INJECT1_1 = "NO";
    CCU2C add_5422_15 (.A0(amdemod_out_d_11__N_2410[12]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17918), .S0(n34_adj_6200));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam add_5422_15.INIT0 = 16'haaa0;
    defparam add_5422_15.INIT1 = 16'h0000;
    defparam add_5422_15.INJECT1_0 = "NO";
    defparam add_5422_15.INJECT1_1 = "NO";
    L6MUX21 i8598 (.D0(n19629), .D1(n19626), .SD(n19822), .Z(n19630));
    PFUMX i8462 (.BLUT(n19441), .ALUT(n19440), .C0(rx_byte[2]), .Z(n19442));
    PFUMX i8596 (.BLUT(n19628), .ALUT(n19627), .C0(led_0_6), .Z(n19629));
    PFUMX i8593 (.BLUT(n19625), .ALUT(n19624), .C0(rx_byte[2]), .Z(n19626));
    PWM pwm_inst (.\data_in_reg[0] (data_in_reg[0]), .clk_80mhz(clk_80mhz), 
        .\data_in_reg_11__N_2898[0] (data_in_reg_11__N_2898[0]), .\data_in_reg[9] (data_in_reg[9]), 
        .\data_in_reg[8] (data_in_reg[8]), .\data_in_reg_11__N_2898[8] (data_in_reg_11__N_2898[8]), 
        .\data_in_reg[7] (data_in_reg[7]), .\data_in_reg_11__N_2898[7] (data_in_reg_11__N_2898[7]), 
        .\data_in_reg[6] (data_in_reg[6]), .\data_in_reg_11__N_2898[6] (data_in_reg_11__N_2898[6]), 
        .\data_in_reg[5] (data_in_reg[5]), .\data_in_reg_11__N_2898[5] (data_in_reg_11__N_2898[5]), 
        .\data_in_reg[4] (data_in_reg[4]), .\data_in_reg_11__N_2898[4] (data_in_reg_11__N_2898[4]), 
        .\data_in_reg[3] (data_in_reg[3]), .\data_in_reg_11__N_2898[3] (data_in_reg_11__N_2898[3]), 
        .\data_in_reg[2] (data_in_reg[2]), .\data_in_reg_11__N_2898[2] (data_in_reg_11__N_2898[2]), 
        .\data_in_reg[1] (data_in_reg[1]), .\data_in_reg_11__N_2898[1] (data_in_reg_11__N_2898[1]), 
        .count({count_adj_6635}), .\amdemod_out[9] (amdemod_out[9]), .GND_net(GND_net), 
        .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(233[5] 237[5])
    PFUMX mux_1918_i1 (.BLUT(n3318), .ALUT(n3324), .C0(n19300), .Z(n3327));
    L6MUX21 i8456 (.D0(n19435), .D1(n19431), .SD(n19822), .Z(n19436));
    PFUMX i8454 (.BLUT(n19434), .ALUT(n19433), .C0(led_0_6), .Z(n19435));
    LUT4 phase_increment_1__63__N_21_43__bdd_2_lut_8578 (.A(phase_increment_1__63__N_17[43]), 
         .B(led_0_6), .Z(n19604)) /* synthesis lut_function=(A+(B)) */ ;
    defparam phase_increment_1__63__N_21_43__bdd_2_lut_8578.init = 16'heeee;
    PFUMX mux_516_i1 (.BLUT(n1428), .ALUT(n1438), .C0(led_0_6), .Z(n1444));
    PFUMX i8451 (.BLUT(n19430), .ALUT(n19429), .C0(rx_byte[2]), .Z(n19431));
    PFUMX mux_551_i1 (.BLUT(n1475), .ALUT(n1485), .C0(led_0_6), .Z(n1491));
    PFUMX mux_586_i1 (.BLUT(n1522), .ALUT(n1532), .C0(led_0_6), .Z(n1538));
    PFUMX mux_658_i1 (.BLUT(n1626), .ALUT(n1632), .C0(n19297), .Z(n1635));
    PFUMX mux_514_i1 (.BLUT(n1433), .ALUT(n1416), .C0(rx_byte[2]), .Z(n1441));
    PFUMX i8579 (.BLUT(n19605), .ALUT(n19604), .C0(rx_byte[2]), .Z(n19606));
    PFUMX mux_549_i1 (.BLUT(n1480), .ALUT(n1465), .C0(rx_byte[2]), .Z(n1488));
    \CIC(REGISTER_WIDTH=72,DECIMATION_RATIO=4096)_U2  cic_cosine_inst (.n67_adj_114({n28_adj_6131, 
            n31_adj_6132, n34_adj_6133, n37_adj_6134, n40_adj_6135, 
            n43_adj_6136, n46_adj_6137, n49_adj_6138, n52_adj_6139, 
            n55_adj_6140, n58_adj_6141, n61_adj_6142}), .\cic_gain[1] (cic_gain[1]), 
            .\comb10[60] (comb10_adj_6571[60]), .n62(n62), .\comb10[59] (comb10_adj_6571[59]), 
            .integrator_tmp({integrator_tmp_adj_6556}), .clk_80mhz(clk_80mhz), 
            .integrator5({integrator5_adj_6562}), .integrator_d_tmp({integrator_d_tmp_adj_6557}), 
            .integrator2({integrator2_adj_6559}), .integrator2_71__N_1032({integrator2_71__N_1032_adj_6574}), 
            .integrator3({integrator3_adj_6560}), .integrator3_71__N_1104({integrator3_71__N_1104_adj_6575}), 
            .integrator4({integrator4_adj_6561}), .integrator4_71__N_1176({integrator4_71__N_1176_adj_6576}), 
            .integrator5_71__N_1248({integrator5_71__N_1248_adj_6577}), .comb6({comb6_adj_6563}), 
            .comb6_71__N_1993({comb6_71__N_1993_adj_6589}), .comb_d6({comb_d6_adj_6564}), 
            .comb7({comb7_adj_6565}), .comb7_71__N_2065({comb7_71__N_2065_adj_6590}), 
            .comb_d7({comb_d7_adj_6566}), .comb8({comb8_adj_6567}), .comb8_71__N_2137({comb8_71__N_2137_adj_6591}), 
            .comb_d8({comb_d8_adj_6568}), .comb9({comb9_adj_6569}), .comb9_71__N_2209({comb9_71__N_2209_adj_6592}), 
            .comb_d9({comb_d9_adj_6570}), .integrator1({integrator1_adj_6558}), 
            .integrator1_71__N_960({integrator1_71__N_960_adj_6573}), .n19(n19_adj_5473), 
            .n18(n18_adj_5472), .n21(n21_adj_5475), .n20(n20_adj_5474), 
            .n23(n23_adj_5477), .n22(n22_adj_5476), .n25(n25_adj_5479), 
            .n24(n24_adj_5478), .n27(n27_adj_5481), .n3(n3_adj_5565), 
            .n2(n2_adj_5564), .n26(n26_adj_5480), .n5(n5_adj_5567), .n29(n29_adj_5483), 
            .n28_adj_1(n28_adj_5482), .n31_adj_2(n31_adj_5485), .\comb10[71] (comb10_adj_6571[71]), 
            .\comb10[70] (comb10_adj_6571[70]), .\comb10[69] (comb10_adj_6571[69]), 
            .\comb10[68] (comb10_adj_6571[68]), .\comb10[67] (comb10_adj_6571[67]), 
            .\comb10[66] (comb10_adj_6571[66]), .\comb10[65] (comb10_adj_6571[65]), 
            .\comb10[64] (comb10_adj_6571[64]), .\comb10[63] (comb10_adj_6571[63]), 
            .\comb10[62] (comb10_adj_6571[62]), .\comb10[61] (comb10_adj_6571[61]), 
            .n30(n30_adj_5484), .n33(n33_adj_5487), .n32(n32_adj_5486), 
            .n35(n35_adj_5489), .n4(n4_adj_5566), .n34_adj_3(n34_adj_5488), 
            .n37_adj_4(n37_adj_5491), .n36(n36_adj_5490), .n7(n7_adj_5569), 
            .n3_adj_5(n3_adj_5493), .n6(n6_adj_5568), .n2_adj_6(n2_adj_5492), 
            .n5_adj_7(n5_adj_5495), .n4_adj_8(n4_adj_5494), .n7_adj_9(n7_adj_5497), 
            .n6_adj_10(n6_adj_5496), .n9(n9_adj_5499), .n8(n8_adj_5498), 
            .n5_adj_11(n5_adj_5459), .n11(n11_adj_5501), .\cic_gain[0] (cic_gain[0]), 
            .n4_adj_12(n4_adj_5458), .n10(n10_adj_5500), .n13(n13_adj_5503), 
            .n12(n12_adj_5502), .n15(n15_adj_5505), .n14(n14_adj_5504), 
            .n17(n17_adj_5507), .n16(n16_adj_5506), .n19_adj_13(n19_adj_5509), 
            .n18_adj_14(n18_adj_5508), .n21_adj_15(n21_adj_5511), .n20_adj_16(n20_adj_5510), 
            .n23_adj_17(n23_adj_5513), .n22_adj_18(n22_adj_5512), .n25_adj_19(n25_adj_5515), 
            .n24_adj_20(n24_adj_5514), .n27_adj_21(n27_adj_5517), .n26_adj_22(n26_adj_5516), 
            .n29_adj_23(n29_adj_5519), .n28_adj_24(n28_adj_5518), .n7_adj_25(n7_adj_5461), 
            .n31_adj_26(n31_adj_5521), .n6_adj_27(n6_adj_5460), .n30_adj_28(n30_adj_5520), 
            .n33_adj_29(n33_adj_5523), .n32_adj_30(n32_adj_5522), .n35_adj_31(n35_adj_5525), 
            .n9_adj_32(n9_adj_5571), .n8_adj_33(n8_adj_5570), .n34_adj_34(n34_adj_5524), 
            .n37_adj_35(n37_adj_5527), .n36_adj_36(n36_adj_5526), .n3_adj_37(n3_adj_5529), 
            .n2_adj_38(n2_adj_5528), .n11_adj_39(n11_adj_5573), .n5_adj_40(n5_adj_5531), 
            .n4_adj_41(n4_adj_5530), .n7_adj_42(n7_adj_5533), .n6_adj_43(n6_adj_5532), 
            .n10_adj_44(n10_adj_5572), .n9_adj_45(n9_adj_5535), .n8_adj_46(n8_adj_5534), 
            .n11_adj_47(n11_adj_5537), .n10_adj_48(n10_adj_5536), .n13_adj_49(n13_adj_5539), 
            .n12_adj_50(n12_adj_5538), .n15_adj_51(n15_adj_5541), .n13_adj_52(n13_adj_5575), 
            .n14_adj_53(n14_adj_5540), .n17_adj_54(n17_adj_5543), .n16_adj_55(n16_adj_5542), 
            .n19_adj_56(n19_adj_5545), .n12_adj_57(n12_adj_5574), .n18_adj_58(n18_adj_5544), 
            .n15_adj_59(n15_adj_5577), .n21_adj_60(n21_adj_5547), .count({count_adj_6572}), 
            .n20_adj_61(n20_adj_5546), .n23_adj_62(n23_adj_5549), .n22_adj_63(n22_adj_5548), 
            .n25_adj_64(n25_adj_5551), .n24_adj_65(n24_adj_5550), .n27_adj_66(n27_adj_5553), 
            .n26_adj_67(n26_adj_5552), .n29_adj_68(n29_adj_5555), .n28_adj_69(n28_adj_5554), 
            .n31_adj_70(n31_adj_5557), .n30_adj_71(n30_adj_5556), .n9_adj_72(n9_adj_5463), 
            .n8_adj_73(n8_adj_5462), .n33_adj_74(n33_adj_5559), .n11_adj_75(n11_adj_5465), 
            .n10_adj_76(n10_adj_5464), .n32_adj_77(n32_adj_5558), .n35_adj_78(n35_adj_5561), 
            .n70(n70), .n68(n68), .n67(n67), .n66(n66_adj_5290), .n65(n65), 
            .n64(n64), .n63(n63_adj_5289), .n34_adj_79(n34_adj_5560), 
            .n37_adj_80(n37_adj_5563), .n36_adj_81(n36_adj_5562), .n13_adj_82(n13_adj_5467), 
            .n12_adj_83(n12_adj_5466), .n14_adj_84(n14_adj_5576), .n15_adj_85(n15_adj_5469), 
            .n17_adj_86(n17_adj_5579), .n16_adj_87(n16_adj_5578), .n14_adj_88(n14_adj_5468), 
            .n19_adj_89(n19_adj_5581), .n18_adj_90(n18_adj_5580), .n21_adj_91(n21_adj_5583), 
            .n20_adj_92(n20_adj_5582), .n61_adj_93(n61_adj_5288), .n23_adj_94(n23_adj_5585), 
            .n22_adj_95(n22_adj_5584), .n25_adj_96(n25_adj_5587), .n17_adj_97(n17_adj_5471), 
            .n16_adj_98(n16_adj_5470), .n24_adj_99(n24_adj_5586), .n27_adj_100(n27_adj_5589), 
            .n26_adj_101(n26_adj_5588), .n76(n76), .n78(n78_adj_5612), 
            .cout(cout_adj_6281), .n79(n79), .n81(n81_adj_5613), .n82(n82), 
            .n84(n84_adj_5614), .n85(n85), .n87(n87_adj_5615), .n88(n88), 
            .n90(n90_adj_5616), .n91(n91), .n93(n93_adj_5617), .n94(n94), 
            .n96(n96_adj_5618), .n97(n97), .n99(n99_adj_5619), .n100(n100), 
            .n102(n102_adj_5620), .n103(n103), .n105(n105_adj_5621), .n106(n106), 
            .n108(n108_adj_5622), .n109(n109), .n111(n111_adj_5623), .n112(n112), 
            .n114(n114_adj_5624), .n115(n115), .n117(n117_adj_5625), .n118(n118), 
            .n120(n120_adj_5626), .n29_adj_102(n29_adj_5591), .n28_adj_103(n28_adj_5590), 
            .n2_adj_104(n2_adj_5456), .n3_adj_105(n3_adj_5457), .n31_adj_106(n31_adj_5593), 
            .n30_adj_107(n30_adj_5592), .n33_adj_108(n33_adj_5595), .n32_adj_109(n32_adj_5594), 
            .n35_adj_110(n35_adj_5597), .n34_adj_111(n34_adj_5596), .n37_adj_112(n37_adj_5599), 
            .n36_adj_113(n36_adj_5598), .\cic_cosine_out[1] (cic_cosine_out[1]), 
            .\cic_cosine_out[0] (cic_cosine_out[0])) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(206[7] 212[6])
    
endmodule
//
// Verilog Description of module quarterwave_generator
//

module quarterwave_generator (clk_80mhz, \phase_accumulator[63] , \lo_sinewave[0] , 
            \lo_cosinewave[0] , \lo_cosinewave[9] , \lo_cosinewave[10] , 
            \lo_sinewave[5] , \lo_cosinewave[6] , \lo_cosinewave[7] , 
            \lo_cosinewave[4] , \lo_cosinewave[5] , \lo_sinewave[6] , 
            \lo_sinewave[9] , \lo_sinewave[10] , \lo_sinewave[12] , \lo_sinewave[8] , 
            \lo_sinewave[7] , \lo_sinewave[2] , \lo_sinewave[3] , \lo_sinewave[4] , 
            \lo_sinewave[1] , sine_table_value, n67, \phase_accumulator[62] , 
            cosine_table_value, n67_adj_464, \phase_accumulator[56] , 
            \phase_accumulator[57] , \phase_accumulator[58] , \phase_accumulator[59] , 
            \phase_accumulator[60] , \phase_accumulator[61] , \lo_cosinewave[12] , 
            \lo_cosinewave[8] , \lo_cosinewave[3] , \lo_cosinewave[2] , 
            \lo_cosinewave[1] , GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input clk_80mhz;
    input \phase_accumulator[63] ;
    output \lo_sinewave[0] ;
    output \lo_cosinewave[0] ;
    output \lo_cosinewave[9] ;
    output \lo_cosinewave[10] ;
    output \lo_sinewave[5] ;
    output \lo_cosinewave[6] ;
    output \lo_cosinewave[7] ;
    output \lo_cosinewave[4] ;
    output \lo_cosinewave[5] ;
    output \lo_sinewave[6] ;
    output \lo_sinewave[9] ;
    output \lo_sinewave[10] ;
    output \lo_sinewave[12] ;
    output \lo_sinewave[8] ;
    output \lo_sinewave[7] ;
    output \lo_sinewave[2] ;
    output \lo_sinewave[3] ;
    output \lo_sinewave[4] ;
    output \lo_sinewave[1] ;
    output [11:0]sine_table_value;
    input [11:0]n67;
    input \phase_accumulator[62] ;
    output [11:0]cosine_table_value;
    input [11:0]n67_adj_464;
    input \phase_accumulator[56] ;
    input \phase_accumulator[57] ;
    input \phase_accumulator[58] ;
    input \phase_accumulator[59] ;
    input \phase_accumulator[60] ;
    input \phase_accumulator[61] ;
    output \lo_cosinewave[12] ;
    output \lo_cosinewave[8] ;
    output \lo_cosinewave[3] ;
    output \lo_cosinewave[2] ;
    output \lo_cosinewave[1] ;
    input GND_net;
    input VCC_net;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(61[34:43])
    wire [1:0]sine_negate;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(15[32:43])
    wire [11:0]sinewave_11__N_733;
    wire [1:0]cosine_negate;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(19[32:45])
    
    wire cosine_negate_1__N_720;
    wire [11:0]cosinewave_11__N_745;
    wire [5:0]sine_index_5__N_721;
    wire [5:0]cosine_index_5__N_727;
    
    FD1S3AX sine_negate_i0 (.D(\phase_accumulator[63] ), .CK(clk_80mhz), 
            .Q(sine_negate[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sine_negate_i0.GSR = "ENABLED";
    FD1S3AX sinewave_i1 (.D(sinewave_11__N_733[0]), .CK(clk_80mhz), .Q(\lo_sinewave[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sinewave_i1.GSR = "ENABLED";
    FD1S3AX cosine_negate_i0 (.D(cosine_negate_1__N_720), .CK(clk_80mhz), 
            .Q(cosine_negate[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosine_negate_i0.GSR = "ENABLED";
    FD1S3AX cosinewave_i1 (.D(cosinewave_11__N_745[0]), .CK(clk_80mhz), 
            .Q(\lo_cosinewave[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosinewave_i1.GSR = "ENABLED";
    FD1S3AX cosinewave_i10 (.D(cosinewave_11__N_745[9]), .CK(clk_80mhz), 
            .Q(\lo_cosinewave[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosinewave_i10.GSR = "ENABLED";
    FD1S3AX cosinewave_i11 (.D(cosinewave_11__N_745[10]), .CK(clk_80mhz), 
            .Q(\lo_cosinewave[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosinewave_i11.GSR = "ENABLED";
    FD1S3AX sinewave_i6 (.D(sinewave_11__N_733[5]), .CK(clk_80mhz), .Q(\lo_sinewave[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sinewave_i6.GSR = "ENABLED";
    FD1S3AX cosinewave_i7 (.D(cosinewave_11__N_745[6]), .CK(clk_80mhz), 
            .Q(\lo_cosinewave[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosinewave_i7.GSR = "ENABLED";
    FD1S3AX cosinewave_i8 (.D(cosinewave_11__N_745[7]), .CK(clk_80mhz), 
            .Q(\lo_cosinewave[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosinewave_i8.GSR = "ENABLED";
    FD1S3AX cosinewave_i5 (.D(cosinewave_11__N_745[4]), .CK(clk_80mhz), 
            .Q(\lo_cosinewave[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosinewave_i5.GSR = "ENABLED";
    FD1S3AX cosinewave_i6 (.D(cosinewave_11__N_745[5]), .CK(clk_80mhz), 
            .Q(\lo_cosinewave[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosinewave_i6.GSR = "ENABLED";
    FD1S3AX sinewave_i7 (.D(sinewave_11__N_733[6]), .CK(clk_80mhz), .Q(\lo_sinewave[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sinewave_i7.GSR = "ENABLED";
    FD1S3AX sinewave_i10 (.D(sinewave_11__N_733[9]), .CK(clk_80mhz), .Q(\lo_sinewave[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sinewave_i10.GSR = "ENABLED";
    FD1S3AX sinewave_i11 (.D(sinewave_11__N_733[10]), .CK(clk_80mhz), .Q(\lo_sinewave[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sinewave_i11.GSR = "ENABLED";
    FD1S3AX sinewave_i12 (.D(sinewave_11__N_733[11]), .CK(clk_80mhz), .Q(\lo_sinewave[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sinewave_i12.GSR = "ENABLED";
    FD1S3AX cosine_negate_i1 (.D(cosine_negate[0]), .CK(clk_80mhz), .Q(cosine_negate[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosine_negate_i1.GSR = "ENABLED";
    FD1S3AX sinewave_i9 (.D(sinewave_11__N_733[8]), .CK(clk_80mhz), .Q(\lo_sinewave[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sinewave_i9.GSR = "ENABLED";
    FD1S3AX sinewave_i8 (.D(sinewave_11__N_733[7]), .CK(clk_80mhz), .Q(\lo_sinewave[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sinewave_i8.GSR = "ENABLED";
    FD1S3AX sinewave_i3 (.D(sinewave_11__N_733[2]), .CK(clk_80mhz), .Q(\lo_sinewave[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sinewave_i3.GSR = "ENABLED";
    FD1S3AX sinewave_i4 (.D(sinewave_11__N_733[3]), .CK(clk_80mhz), .Q(\lo_sinewave[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sinewave_i4.GSR = "ENABLED";
    FD1S3AX sinewave_i5 (.D(sinewave_11__N_733[4]), .CK(clk_80mhz), .Q(\lo_sinewave[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sinewave_i5.GSR = "ENABLED";
    FD1S3AX sinewave_i2 (.D(sinewave_11__N_733[1]), .CK(clk_80mhz), .Q(\lo_sinewave[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sinewave_i2.GSR = "ENABLED";
    FD1S3AX sine_negate_i1 (.D(sine_negate[0]), .CK(clk_80mhz), .Q(sine_negate[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam sine_negate_i1.GSR = "ENABLED";
    LUT4 mux_16_i1_3_lut (.A(sine_table_value[0]), .B(n67[0]), .C(sine_negate[1]), 
         .Z(sinewave_11__N_733[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[29:86])
    defparam mux_16_i1_3_lut.init = 16'hcaca;
    LUT4 phase_accumulator_63__I_0_2_lut (.A(\phase_accumulator[63] ), .B(\phase_accumulator[62] ), 
         .Z(cosine_negate_1__N_720)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(53[29:96])
    defparam phase_accumulator_63__I_0_2_lut.init = 16'h6666;
    LUT4 mux_18_i1_3_lut (.A(cosine_table_value[0]), .B(n67_adj_464[0]), 
         .C(cosine_negate[1]), .Z(cosinewave_11__N_745[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[29:88])
    defparam mux_18_i1_3_lut.init = 16'hcaca;
    LUT4 i4012_2_lut (.A(\phase_accumulator[56] ), .B(\phase_accumulator[62] ), 
         .Z(sine_index_5__N_721[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(58[16] 61[10])
    defparam i4012_2_lut.init = 16'h6666;
    LUT4 i4014_2_lut (.A(\phase_accumulator[57] ), .B(\phase_accumulator[62] ), 
         .Z(sine_index_5__N_721[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(58[16] 61[10])
    defparam i4014_2_lut.init = 16'h6666;
    LUT4 i4021_2_lut (.A(\phase_accumulator[58] ), .B(\phase_accumulator[62] ), 
         .Z(sine_index_5__N_721[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(58[16] 61[10])
    defparam i4021_2_lut.init = 16'h6666;
    LUT4 i4020_2_lut (.A(\phase_accumulator[59] ), .B(\phase_accumulator[62] ), 
         .Z(sine_index_5__N_721[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(58[16] 61[10])
    defparam i4020_2_lut.init = 16'h6666;
    LUT4 i4017_2_lut (.A(\phase_accumulator[60] ), .B(\phase_accumulator[62] ), 
         .Z(sine_index_5__N_721[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(58[16] 61[10])
    defparam i4017_2_lut.init = 16'h6666;
    LUT4 i4018_2_lut (.A(\phase_accumulator[61] ), .B(\phase_accumulator[62] ), 
         .Z(sine_index_5__N_721[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(58[16] 61[10])
    defparam i4018_2_lut.init = 16'h6666;
    LUT4 i8326_2_lut (.A(\phase_accumulator[56] ), .B(\phase_accumulator[62] ), 
         .Z(cosine_index_5__N_727[0])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(58[16] 61[10])
    defparam i8326_2_lut.init = 16'h9999;
    LUT4 i8332_2_lut (.A(\phase_accumulator[57] ), .B(\phase_accumulator[62] ), 
         .Z(cosine_index_5__N_727[1])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(58[16] 61[10])
    defparam i8332_2_lut.init = 16'h9999;
    LUT4 i8336_2_lut (.A(\phase_accumulator[58] ), .B(\phase_accumulator[62] ), 
         .Z(cosine_index_5__N_727[2])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(58[16] 61[10])
    defparam i8336_2_lut.init = 16'h9999;
    LUT4 i8334_2_lut (.A(\phase_accumulator[59] ), .B(\phase_accumulator[62] ), 
         .Z(cosine_index_5__N_727[3])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(58[16] 61[10])
    defparam i8334_2_lut.init = 16'h9999;
    LUT4 i8330_2_lut (.A(\phase_accumulator[60] ), .B(\phase_accumulator[62] ), 
         .Z(cosine_index_5__N_727[4])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(58[16] 61[10])
    defparam i8330_2_lut.init = 16'h9999;
    LUT4 i8328_2_lut (.A(\phase_accumulator[61] ), .B(\phase_accumulator[62] ), 
         .Z(cosine_index_5__N_727[5])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(58[16] 61[10])
    defparam i8328_2_lut.init = 16'h9999;
    FD1S3AX cosinewave_i12 (.D(cosinewave_11__N_745[11]), .CK(clk_80mhz), 
            .Q(\lo_cosinewave[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosinewave_i12.GSR = "ENABLED";
    FD1S3AX cosinewave_i9 (.D(cosinewave_11__N_745[8]), .CK(clk_80mhz), 
            .Q(\lo_cosinewave[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosinewave_i9.GSR = "ENABLED";
    FD1S3AX cosinewave_i4 (.D(cosinewave_11__N_745[3]), .CK(clk_80mhz), 
            .Q(\lo_cosinewave[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosinewave_i4.GSR = "ENABLED";
    FD1S3AX cosinewave_i3 (.D(cosinewave_11__N_745[2]), .CK(clk_80mhz), 
            .Q(\lo_cosinewave[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosinewave_i3.GSR = "ENABLED";
    FD1S3AX cosinewave_i2 (.D(cosinewave_11__N_745[1]), .CK(clk_80mhz), 
            .Q(\lo_cosinewave[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=158, LSE_RLINE=165 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(50[14] 68[8])
    defparam cosinewave_i2.GSR = "ENABLED";
    LUT4 mux_18_i10_3_lut (.A(cosine_table_value[9]), .B(n67_adj_464[9]), 
         .C(cosine_negate[1]), .Z(cosinewave_11__N_745[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[29:88])
    defparam mux_18_i10_3_lut.init = 16'hcaca;
    LUT4 mux_18_i11_3_lut (.A(cosine_table_value[10]), .B(n67_adj_464[10]), 
         .C(cosine_negate[1]), .Z(cosinewave_11__N_745[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[29:88])
    defparam mux_18_i11_3_lut.init = 16'hcaca;
    LUT4 mux_16_i6_3_lut (.A(sine_table_value[5]), .B(n67[5]), .C(sine_negate[1]), 
         .Z(sinewave_11__N_733[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[29:86])
    defparam mux_16_i6_3_lut.init = 16'hcaca;
    LUT4 mux_18_i7_3_lut (.A(cosine_table_value[6]), .B(n67_adj_464[6]), 
         .C(cosine_negate[1]), .Z(cosinewave_11__N_745[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[29:88])
    defparam mux_18_i7_3_lut.init = 16'hcaca;
    LUT4 mux_18_i8_3_lut (.A(cosine_table_value[7]), .B(n67_adj_464[7]), 
         .C(cosine_negate[1]), .Z(cosinewave_11__N_745[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[29:88])
    defparam mux_18_i8_3_lut.init = 16'hcaca;
    LUT4 mux_18_i5_3_lut (.A(cosine_table_value[4]), .B(n67_adj_464[4]), 
         .C(cosine_negate[1]), .Z(cosinewave_11__N_745[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[29:88])
    defparam mux_18_i5_3_lut.init = 16'hcaca;
    LUT4 mux_18_i6_3_lut (.A(cosine_table_value[5]), .B(n67_adj_464[5]), 
         .C(cosine_negate[1]), .Z(cosinewave_11__N_745[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[29:88])
    defparam mux_18_i6_3_lut.init = 16'hcaca;
    LUT4 mux_16_i7_3_lut (.A(sine_table_value[6]), .B(n67[6]), .C(sine_negate[1]), 
         .Z(sinewave_11__N_733[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[29:86])
    defparam mux_16_i7_3_lut.init = 16'hcaca;
    LUT4 mux_16_i10_3_lut (.A(sine_table_value[9]), .B(n67[9]), .C(sine_negate[1]), 
         .Z(sinewave_11__N_733[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[29:86])
    defparam mux_16_i10_3_lut.init = 16'hcaca;
    LUT4 mux_16_i11_3_lut (.A(sine_table_value[10]), .B(n67[10]), .C(sine_negate[1]), 
         .Z(sinewave_11__N_733[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[29:86])
    defparam mux_16_i11_3_lut.init = 16'hcaca;
    LUT4 mux_16_i12_3_lut (.A(sine_table_value[11]), .B(n67[11]), .C(sine_negate[1]), 
         .Z(sinewave_11__N_733[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[29:86])
    defparam mux_16_i12_3_lut.init = 16'hcaca;
    LUT4 mux_16_i9_3_lut (.A(sine_table_value[8]), .B(n67[8]), .C(sine_negate[1]), 
         .Z(sinewave_11__N_733[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[29:86])
    defparam mux_16_i9_3_lut.init = 16'hcaca;
    LUT4 mux_16_i8_3_lut (.A(sine_table_value[7]), .B(n67[7]), .C(sine_negate[1]), 
         .Z(sinewave_11__N_733[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[29:86])
    defparam mux_16_i8_3_lut.init = 16'hcaca;
    LUT4 mux_16_i3_3_lut (.A(sine_table_value[2]), .B(n67[2]), .C(sine_negate[1]), 
         .Z(sinewave_11__N_733[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[29:86])
    defparam mux_16_i3_3_lut.init = 16'hcaca;
    LUT4 mux_16_i4_3_lut (.A(sine_table_value[3]), .B(n67[3]), .C(sine_negate[1]), 
         .Z(sinewave_11__N_733[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[29:86])
    defparam mux_16_i4_3_lut.init = 16'hcaca;
    LUT4 mux_16_i5_3_lut (.A(sine_table_value[4]), .B(n67[4]), .C(sine_negate[1]), 
         .Z(sinewave_11__N_733[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[29:86])
    defparam mux_16_i5_3_lut.init = 16'hcaca;
    LUT4 mux_16_i2_3_lut (.A(sine_table_value[1]), .B(n67[1]), .C(sine_negate[1]), 
         .Z(sinewave_11__N_733[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(66[29:86])
    defparam mux_16_i2_3_lut.init = 16'hcaca;
    LUT4 mux_18_i12_3_lut (.A(cosine_table_value[11]), .B(n67_adj_464[11]), 
         .C(cosine_negate[1]), .Z(cosinewave_11__N_745[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[29:88])
    defparam mux_18_i12_3_lut.init = 16'hcaca;
    LUT4 mux_18_i9_3_lut (.A(cosine_table_value[8]), .B(n67_adj_464[8]), 
         .C(cosine_negate[1]), .Z(cosinewave_11__N_745[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[29:88])
    defparam mux_18_i9_3_lut.init = 16'hcaca;
    LUT4 mux_18_i4_3_lut (.A(cosine_table_value[3]), .B(n67_adj_464[3]), 
         .C(cosine_negate[1]), .Z(cosinewave_11__N_745[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[29:88])
    defparam mux_18_i4_3_lut.init = 16'hcaca;
    LUT4 mux_18_i3_3_lut (.A(cosine_table_value[2]), .B(n67_adj_464[2]), 
         .C(cosine_negate[1]), .Z(cosinewave_11__N_745[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[29:88])
    defparam mux_18_i3_3_lut.init = 16'hcaca;
    LUT4 mux_18_i2_3_lut (.A(cosine_table_value[1]), .B(n67_adj_464[1]), 
         .C(cosine_negate[1]), .Z(cosinewave_11__N_745[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(67[29:88])
    defparam mux_18_i2_3_lut.init = 16'hcaca;
    quarterwave_table sinewave_inst (.sine_index_5__N_721({sine_index_5__N_721}), 
            .sine_table_value({sine_table_value}), .clk_80mhz(clk_80mhz), 
            .GND_net(GND_net), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(26[75] 29[4])
    quarterwave_table_U0 cosinewave_inst (.cosine_index_5__N_727({cosine_index_5__N_727}), 
            .cosine_table_value({cosine_table_value}), .clk_80mhz(clk_80mhz), 
            .GND_net(GND_net), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/quarterwave_generator.v(31[75] 34[4])
    
endmodule
//
// Verilog Description of module quarterwave_table
//

module quarterwave_table (sine_index_5__N_721, sine_table_value, clk_80mhz, 
            GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input [5:0]sine_index_5__N_721;
    output [11:0]sine_table_value;
    input clk_80mhz;
    input GND_net;
    input VCC_net;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(61[34:43])
    
    PDPW16KD address_5__I_0 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), 
            .DI3(GND_net), .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .DI18(GND_net), 
            .DI19(GND_net), .DI20(GND_net), .DI21(GND_net), .DI22(GND_net), 
            .DI23(GND_net), .DI24(GND_net), .DI25(GND_net), .DI26(GND_net), 
            .DI27(GND_net), .DI28(GND_net), .DI29(GND_net), .DI30(GND_net), 
            .DI31(GND_net), .DI32(GND_net), .DI33(GND_net), .DI34(GND_net), 
            .DI35(GND_net), .ADW0(GND_net), .ADW1(GND_net), .ADW2(GND_net), 
            .ADW3(GND_net), .ADW4(GND_net), .ADW5(GND_net), .ADW6(GND_net), 
            .ADW7(GND_net), .ADW8(GND_net), .BE0(GND_net), .BE1(GND_net), 
            .BE2(GND_net), .BE3(GND_net), .CEW(VCC_net), .CLKW(GND_net), 
            .CSW0(GND_net), .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), 
            .ADR1(GND_net), .ADR2(GND_net), .ADR3(GND_net), .ADR4(sine_index_5__N_721[0]), 
            .ADR5(sine_index_5__N_721[1]), .ADR6(sine_index_5__N_721[2]), 
            .ADR7(sine_index_5__N_721[3]), .ADR8(sine_index_5__N_721[4]), 
            .ADR9(sine_index_5__N_721[5]), .ADR10(GND_net), .ADR11(GND_net), 
            .ADR12(GND_net), .ADR13(GND_net), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(clk_80mhz), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(sine_table_value[0]), .DO1(sine_table_value[1]), 
            .DO2(sine_table_value[2]), .DO3(sine_table_value[3]), .DO4(sine_table_value[4]), 
            .DO5(sine_table_value[5]), .DO6(sine_table_value[6]), .DO7(sine_table_value[7]), 
            .DO8(sine_table_value[8]), .DO9(sine_table_value[9]), .DO10(sine_table_value[10]), 
            .DO11(sine_table_value[11]));
    defparam address_5__I_0.DATA_WIDTH_W = 36;
    defparam address_5__I_0.DATA_WIDTH_R = 18;
    defparam address_5__I_0.GSR = "DISABLED";
    defparam address_5__I_0.REGMODE = "NOREG";
    defparam address_5__I_0.RESETMODE = "ASYNC";
    defparam address_5__I_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam address_5__I_0.CSDECODE_W = "0b000";
    defparam address_5__I_0.CSDECODE_R = "0b000";
    defparam address_5__I_0.INITVAL_00 = "0x002F8002C9002990026A0023A00209001D8001A7001760014500113000E1000AF0007D0004B00019";
    defparam address_5__I_0.INITVAL_01 = "0x00595005710054B00525004FF004D7004AF004860045C0043100406003DB003AE003810035400326";
    defparam address_5__I_0.INITVAL_02 = "0x00759007450072F0071800701006E8006CE006B3006970067B0065D0063E0061E005FD005DB005B9";
    defparam address_5__I_0.INITVAL_03 = "0x007FE007FD007FB007F7007F2007EC007E5007DC007D2007C7007BB007AE0079F0078F0077E0076C";
    defparam address_5__I_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INIT_DATA = "STATIC";
    
endmodule
//
// Verilog Description of module quarterwave_table_U0
//

module quarterwave_table_U0 (cosine_index_5__N_727, cosine_table_value, 
            clk_80mhz, GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input [5:0]cosine_index_5__N_727;
    output [11:0]cosine_table_value;
    input clk_80mhz;
    input GND_net;
    input VCC_net;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(61[34:43])
    
    PDPW16KD address_5__I_0 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), 
            .DI3(GND_net), .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .DI18(GND_net), 
            .DI19(GND_net), .DI20(GND_net), .DI21(GND_net), .DI22(GND_net), 
            .DI23(GND_net), .DI24(GND_net), .DI25(GND_net), .DI26(GND_net), 
            .DI27(GND_net), .DI28(GND_net), .DI29(GND_net), .DI30(GND_net), 
            .DI31(GND_net), .DI32(GND_net), .DI33(GND_net), .DI34(GND_net), 
            .DI35(GND_net), .ADW0(GND_net), .ADW1(GND_net), .ADW2(GND_net), 
            .ADW3(GND_net), .ADW4(GND_net), .ADW5(GND_net), .ADW6(GND_net), 
            .ADW7(GND_net), .ADW8(GND_net), .BE0(GND_net), .BE1(GND_net), 
            .BE2(GND_net), .BE3(GND_net), .CEW(VCC_net), .CLKW(GND_net), 
            .CSW0(GND_net), .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), 
            .ADR1(GND_net), .ADR2(GND_net), .ADR3(GND_net), .ADR4(cosine_index_5__N_727[0]), 
            .ADR5(cosine_index_5__N_727[1]), .ADR6(cosine_index_5__N_727[2]), 
            .ADR7(cosine_index_5__N_727[3]), .ADR8(cosine_index_5__N_727[4]), 
            .ADR9(cosine_index_5__N_727[5]), .ADR10(GND_net), .ADR11(GND_net), 
            .ADR12(GND_net), .ADR13(GND_net), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(clk_80mhz), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(cosine_table_value[0]), .DO1(cosine_table_value[1]), 
            .DO2(cosine_table_value[2]), .DO3(cosine_table_value[3]), .DO4(cosine_table_value[4]), 
            .DO5(cosine_table_value[5]), .DO6(cosine_table_value[6]), .DO7(cosine_table_value[7]), 
            .DO8(cosine_table_value[8]), .DO9(cosine_table_value[9]), .DO10(cosine_table_value[10]), 
            .DO11(cosine_table_value[11]));
    defparam address_5__I_0.DATA_WIDTH_W = 36;
    defparam address_5__I_0.DATA_WIDTH_R = 18;
    defparam address_5__I_0.GSR = "DISABLED";
    defparam address_5__I_0.REGMODE = "NOREG";
    defparam address_5__I_0.RESETMODE = "ASYNC";
    defparam address_5__I_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam address_5__I_0.CSDECODE_W = "0b000";
    defparam address_5__I_0.CSDECODE_R = "0b000";
    defparam address_5__I_0.INITVAL_00 = "0x002F8002C9002990026A0023A00209001D8001A7001760014500113000E1000AF0007D0004B00019";
    defparam address_5__I_0.INITVAL_01 = "0x00595005710054B00525004FF004D7004AF004860045C0043100406003DB003AE003810035400326";
    defparam address_5__I_0.INITVAL_02 = "0x00759007450072F0071800701006E8006CE006B3006970067B0065D0063E0061E005FD005DB005B9";
    defparam address_5__I_0.INITVAL_03 = "0x007FE007FD007FB007F7007F2007EC007E5007DC007D2007C7007BB007AE0079F0078F0077E0076C";
    defparam address_5__I_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam address_5__I_0.INIT_DATA = "STATIC";
    
endmodule
//
// Verilog Description of module Mixer
//

module Mixer (mix_sinewave, clk_80mhz, mix_cosinewave, diff_out_c, rf_in_c, 
            \lo_sinewave[0] , n67, \lo_sinewave[8] , \lo_cosinewave[0] , 
            n67_adj_451, \lo_sinewave[9] , \lo_sinewave[12] , \lo_sinewave[10] , 
            \lo_sinewave[6] , \lo_sinewave[3] , \lo_cosinewave[12] , \lo_cosinewave[10] , 
            \lo_cosinewave[9] , \lo_cosinewave[8] , \lo_cosinewave[7] , 
            \lo_cosinewave[6] , \lo_cosinewave[5] , \lo_cosinewave[4] , 
            \lo_cosinewave[3] , \lo_cosinewave[2] , \lo_cosinewave[1] , 
            \lo_sinewave[1] , \lo_sinewave[2] , \lo_sinewave[4] , \lo_sinewave[5] , 
            \lo_sinewave[7] ) /* synthesis syn_module_defined=1 */ ;
    output [11:0]mix_sinewave;
    input clk_80mhz;
    output [11:0]mix_cosinewave;
    output diff_out_c;
    input rf_in_c;
    input \lo_sinewave[0] ;
    input [11:0]n67;
    input \lo_sinewave[8] ;
    input \lo_cosinewave[0] ;
    input [11:0]n67_adj_451;
    input \lo_sinewave[9] ;
    input \lo_sinewave[12] ;
    input \lo_sinewave[10] ;
    input \lo_sinewave[6] ;
    input \lo_sinewave[3] ;
    input \lo_cosinewave[12] ;
    input \lo_cosinewave[10] ;
    input \lo_cosinewave[9] ;
    input \lo_cosinewave[8] ;
    input \lo_cosinewave[7] ;
    input \lo_cosinewave[6] ;
    input \lo_cosinewave[5] ;
    input \lo_cosinewave[4] ;
    input \lo_cosinewave[3] ;
    input \lo_cosinewave[2] ;
    input \lo_cosinewave[1] ;
    input \lo_sinewave[1] ;
    input \lo_sinewave[2] ;
    input \lo_sinewave[4] ;
    input \lo_sinewave[5] ;
    input \lo_sinewave[7] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(61[34:43])
    wire [11:0]sinewave_out_11__N_757;
    wire [11:0]cosinewave_out_11__N_769;
    wire [1:0]rf_in_d;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(32[13:20])
    
    FD1S3AX sinewave_out_i7 (.D(sinewave_out_11__N_757[7]), .CK(clk_80mhz), 
            .Q(mix_sinewave[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam sinewave_out_i7.GSR = "ENABLED";
    FD1S3AX sinewave_out_i0 (.D(sinewave_out_11__N_757[0]), .CK(clk_80mhz), 
            .Q(mix_sinewave[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam sinewave_out_i0.GSR = "ENABLED";
    FD1S3AX sinewave_out_i8 (.D(sinewave_out_11__N_757[8]), .CK(clk_80mhz), 
            .Q(mix_sinewave[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam sinewave_out_i8.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i0 (.D(cosinewave_out_11__N_769[0]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam cosinewave_out_i0.GSR = "ENABLED";
    FD1S3AY rf_in_d_i1 (.D(rf_in_c), .CK(clk_80mhz), .Q(diff_out_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(35[10] 38[6])
    defparam rf_in_d_i1.GSR = "ENABLED";
    FD1S3AX sinewave_out_i9 (.D(sinewave_out_11__N_757[9]), .CK(clk_80mhz), 
            .Q(mix_sinewave[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam sinewave_out_i9.GSR = "ENABLED";
    FD1S3AX sinewave_out_i11 (.D(sinewave_out_11__N_757[11]), .CK(clk_80mhz), 
            .Q(mix_sinewave[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam sinewave_out_i11.GSR = "ENABLED";
    FD1S3AX sinewave_out_i10 (.D(sinewave_out_11__N_757[10]), .CK(clk_80mhz), 
            .Q(mix_sinewave[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam sinewave_out_i10.GSR = "ENABLED";
    FD1S3AX sinewave_out_i6 (.D(sinewave_out_11__N_757[6]), .CK(clk_80mhz), 
            .Q(mix_sinewave[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam sinewave_out_i6.GSR = "ENABLED";
    FD1S3AX sinewave_out_i3 (.D(sinewave_out_11__N_757[3]), .CK(clk_80mhz), 
            .Q(mix_sinewave[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam sinewave_out_i3.GSR = "ENABLED";
    LUT4 mux_8_i1_3_lut (.A(\lo_sinewave[0] ), .B(n67[0]), .C(rf_in_d[1]), 
         .Z(sinewave_out_11__N_757[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_8_i1_3_lut.init = 16'hcaca;
    LUT4 mux_8_i9_3_lut (.A(\lo_sinewave[8] ), .B(n67[8]), .C(rf_in_d[1]), 
         .Z(sinewave_out_11__N_757[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_8_i9_3_lut.init = 16'hcaca;
    LUT4 mux_9_i1_3_lut (.A(\lo_cosinewave[0] ), .B(n67_adj_451[0]), .C(rf_in_d[1]), 
         .Z(cosinewave_out_11__N_769[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_9_i1_3_lut.init = 16'hcaca;
    LUT4 mux_8_i10_3_lut (.A(\lo_sinewave[9] ), .B(n67[9]), .C(rf_in_d[1]), 
         .Z(sinewave_out_11__N_757[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_8_i10_3_lut.init = 16'hcaca;
    FD1S3AY rf_in_d_i2 (.D(diff_out_c), .CK(clk_80mhz), .Q(rf_in_d[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(35[10] 38[6])
    defparam rf_in_d_i2.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i11 (.D(cosinewave_out_11__N_769[11]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam cosinewave_out_i11.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i10 (.D(cosinewave_out_11__N_769[10]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam cosinewave_out_i10.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i9 (.D(cosinewave_out_11__N_769[9]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam cosinewave_out_i9.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i8 (.D(cosinewave_out_11__N_769[8]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam cosinewave_out_i8.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i7 (.D(cosinewave_out_11__N_769[7]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam cosinewave_out_i7.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i6 (.D(cosinewave_out_11__N_769[6]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam cosinewave_out_i6.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i5 (.D(cosinewave_out_11__N_769[5]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam cosinewave_out_i5.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i4 (.D(cosinewave_out_11__N_769[4]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam cosinewave_out_i4.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i3 (.D(cosinewave_out_11__N_769[3]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam cosinewave_out_i3.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i2 (.D(cosinewave_out_11__N_769[2]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam cosinewave_out_i2.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i1 (.D(cosinewave_out_11__N_769[1]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam cosinewave_out_i1.GSR = "ENABLED";
    FD1S3AX sinewave_out_i1 (.D(sinewave_out_11__N_757[1]), .CK(clk_80mhz), 
            .Q(mix_sinewave[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam sinewave_out_i1.GSR = "ENABLED";
    FD1S3AX sinewave_out_i2 (.D(sinewave_out_11__N_757[2]), .CK(clk_80mhz), 
            .Q(mix_sinewave[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam sinewave_out_i2.GSR = "ENABLED";
    FD1S3AX sinewave_out_i4 (.D(sinewave_out_11__N_757[4]), .CK(clk_80mhz), 
            .Q(mix_sinewave[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam sinewave_out_i4.GSR = "ENABLED";
    FD1S3AX sinewave_out_i5 (.D(sinewave_out_11__N_757[5]), .CK(clk_80mhz), 
            .Q(mix_sinewave[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=172, LSE_RLINE=180 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(46[10] 54[6])
    defparam sinewave_out_i5.GSR = "ENABLED";
    LUT4 mux_8_i12_3_lut (.A(\lo_sinewave[12] ), .B(n67[11]), .C(rf_in_d[1]), 
         .Z(sinewave_out_11__N_757[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_8_i12_3_lut.init = 16'hcaca;
    LUT4 mux_8_i11_3_lut (.A(\lo_sinewave[10] ), .B(n67[10]), .C(rf_in_d[1]), 
         .Z(sinewave_out_11__N_757[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_8_i11_3_lut.init = 16'hcaca;
    LUT4 mux_8_i7_3_lut (.A(\lo_sinewave[6] ), .B(n67[6]), .C(rf_in_d[1]), 
         .Z(sinewave_out_11__N_757[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_8_i7_3_lut.init = 16'hcaca;
    LUT4 mux_8_i4_3_lut (.A(\lo_sinewave[3] ), .B(n67[3]), .C(rf_in_d[1]), 
         .Z(sinewave_out_11__N_757[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_8_i4_3_lut.init = 16'hcaca;
    LUT4 mux_9_i12_3_lut (.A(\lo_cosinewave[12] ), .B(n67_adj_451[11]), 
         .C(rf_in_d[1]), .Z(cosinewave_out_11__N_769[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_9_i12_3_lut.init = 16'hcaca;
    LUT4 mux_9_i11_3_lut (.A(\lo_cosinewave[10] ), .B(n67_adj_451[10]), 
         .C(rf_in_d[1]), .Z(cosinewave_out_11__N_769[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_9_i11_3_lut.init = 16'hcaca;
    LUT4 mux_9_i10_3_lut (.A(\lo_cosinewave[9] ), .B(n67_adj_451[9]), .C(rf_in_d[1]), 
         .Z(cosinewave_out_11__N_769[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_9_i10_3_lut.init = 16'hcaca;
    LUT4 mux_9_i9_3_lut (.A(\lo_cosinewave[8] ), .B(n67_adj_451[8]), .C(rf_in_d[1]), 
         .Z(cosinewave_out_11__N_769[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_9_i9_3_lut.init = 16'hcaca;
    LUT4 mux_9_i8_3_lut (.A(\lo_cosinewave[7] ), .B(n67_adj_451[7]), .C(rf_in_d[1]), 
         .Z(cosinewave_out_11__N_769[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_9_i8_3_lut.init = 16'hcaca;
    LUT4 mux_9_i7_3_lut (.A(\lo_cosinewave[6] ), .B(n67_adj_451[6]), .C(rf_in_d[1]), 
         .Z(cosinewave_out_11__N_769[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_9_i7_3_lut.init = 16'hcaca;
    LUT4 mux_9_i6_3_lut (.A(\lo_cosinewave[5] ), .B(n67_adj_451[5]), .C(rf_in_d[1]), 
         .Z(cosinewave_out_11__N_769[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_9_i6_3_lut.init = 16'hcaca;
    LUT4 mux_9_i5_3_lut (.A(\lo_cosinewave[4] ), .B(n67_adj_451[4]), .C(rf_in_d[1]), 
         .Z(cosinewave_out_11__N_769[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_9_i5_3_lut.init = 16'hcaca;
    LUT4 mux_9_i4_3_lut (.A(\lo_cosinewave[3] ), .B(n67_adj_451[3]), .C(rf_in_d[1]), 
         .Z(cosinewave_out_11__N_769[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_9_i4_3_lut.init = 16'hcaca;
    LUT4 mux_9_i3_3_lut (.A(\lo_cosinewave[2] ), .B(n67_adj_451[2]), .C(rf_in_d[1]), 
         .Z(cosinewave_out_11__N_769[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_9_i3_3_lut.init = 16'hcaca;
    LUT4 mux_9_i2_3_lut (.A(\lo_cosinewave[1] ), .B(n67_adj_451[1]), .C(rf_in_d[1]), 
         .Z(cosinewave_out_11__N_769[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_9_i2_3_lut.init = 16'hcaca;
    LUT4 mux_8_i2_3_lut (.A(\lo_sinewave[1] ), .B(n67[1]), .C(rf_in_d[1]), 
         .Z(sinewave_out_11__N_757[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_8_i2_3_lut.init = 16'hcaca;
    LUT4 mux_8_i3_3_lut (.A(\lo_sinewave[2] ), .B(n67[2]), .C(rf_in_d[1]), 
         .Z(sinewave_out_11__N_757[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_8_i3_3_lut.init = 16'hcaca;
    LUT4 mux_8_i5_3_lut (.A(\lo_sinewave[4] ), .B(n67[4]), .C(rf_in_d[1]), 
         .Z(sinewave_out_11__N_757[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_8_i5_3_lut.init = 16'hcaca;
    LUT4 mux_8_i6_3_lut (.A(\lo_sinewave[5] ), .B(n67[5]), .C(rf_in_d[1]), 
         .Z(sinewave_out_11__N_757[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_8_i6_3_lut.init = 16'hcaca;
    LUT4 mux_8_i8_3_lut (.A(\lo_sinewave[7] ), .B(n67[7]), .C(rf_in_d[1]), 
         .Z(sinewave_out_11__N_757[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Mixer.v(50[14] 53[8])
    defparam mux_8_i8_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=87) 
//

module \uart_rx(CLKS_PER_BIT=87)  (rx_byte1, clk_80mhz, rx_serial_c, GND_net, 
            VCC_net, rx_data_valid1) /* synthesis syn_module_defined=1 */ ;
    output [7:0]rx_byte1;
    input clk_80mhz;
    input rx_serial_c;
    input GND_net;
    input VCC_net;
    output rx_data_valid1;
    
    wire [7:0]UartClk /* synthesis SET_AS_NETWORK=\uart_rx_inst/UartClk[2], is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(37[14:21])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(61[34:43])
    wire [15:0]r_Clock_Count;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(39[18:31])
    
    wire UartClk_2_enable_34, n14275;
    wire [15:0]n69;
    wire [7:0]r_Rx_Byte;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(41[17:26])
    
    wire UartClk_2_enable_2, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(40[17:28])
    
    wire UartClk_2_enable_36, n18685, UartClk_2_enable_4, UartClk_2_enable_17, 
        UartClk_2_enable_13, n19817, UartClk_2_enable_14, UartClk_2_enable_15;
    wire [2:0]r_SM_Main;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(43[17:26])
    
    wire n19415, r_Rx_DV_last, r_Rx_DV, r_Rx_Data_R, UartClk_2_enable_16, 
        UartClk_2_enable_19, n18523, n19820, n18566, n18579;
    wire [2:0]r_SM_Main_2__N_2965;
    
    wire n18732, n24, n19821, n17972, n18744, n18528, n18736, 
        n26, n18623, n18714, n18716, n18708, n18712, n14677, n14691, 
        n19414, n19849, n14667, n18750, n18560;
    wire [2:0]n30;
    wire [2:0]n17;
    
    wire n19413, n19848, n18550, n19847, n17064, n17063, n17062, 
        n17061, n17060, n17059, n17058, n17057, n19829, UartClk_2_enable_35, 
        UartClk_2_enable_29, UartClk_2_enable_28, n14269, r_Rx_DV_last_N_3024, 
        r_Rx_DV_N_3025, n17892;
    
    FD1P3IX r_Clock_Count_3041__i9 (.D(n69[9]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i9.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i2 (.D(r_Rx_Data), .SP(UartClk_2_enable_2), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i2 (.D(n18685), .SP(UartClk_2_enable_36), .CK(UartClk[2]), 
            .Q(r_Bit_Index[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i2.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i3 (.D(r_Rx_Data), .SP(UartClk_2_enable_4), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i3.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i7 (.D(r_Rx_Byte[7]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(rx_byte1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i6 (.D(r_Rx_Byte[6]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(rx_byte1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i5 (.D(r_Rx_Byte[5]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(rx_byte1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i4 (.D(r_Rx_Byte[4]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(rx_byte1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i3 (.D(r_Rx_Byte[3]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(rx_byte1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i2 (.D(r_Rx_Byte[2]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(rx_byte1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i1 (.D(r_Rx_Byte[1]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(rx_byte1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_3041__i8 (.D(n69[8]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i8.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i4 (.D(r_Rx_Data), .SP(UartClk_2_enable_13), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i4.GSR = "ENABLED";
    LUT4 i8355_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n19817), .C(r_Bit_Index[1]), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_2)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(114[17:39])
    defparam i8355_2_lut_3_lut_4_lut.init = 16'h0010;
    FD1P3AX r_Rx_Byte_i5 (.D(r_Rx_Data), .SP(UartClk_2_enable_14), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i6 (.D(r_Rx_Data), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i6.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i0 (.D(n19415), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i0.GSR = "ENABLED";
    FD1S3AX r_Rx_DV_last_60 (.D(r_Rx_DV), .CK(clk_80mhz), .Q(r_Rx_DV_last)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(47[11] 52[8])
    defparam r_Rx_DV_last_60.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_R_61 (.D(rx_serial_c), .CK(UartClk[2]), .Q(r_Rx_Data_R)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(57[11] 62[8])
    defparam r_Rx_Data_R_61.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_62 (.D(r_Rx_Data_R), .CK(UartClk[2]), .Q(r_Rx_Data)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(57[11] 62[8])
    defparam r_Rx_Data_62.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i7 (.D(r_Rx_Data), .SP(UartClk_2_enable_16), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i7.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i0 (.D(r_Rx_Byte[0]), .SP(UartClk_2_enable_17), .CK(UartClk[2]), 
            .Q(rx_byte1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i0.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_3041__i7 (.D(n69[7]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i7.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i0 (.D(n18523), .SP(UartClk_2_enable_19), .CK(UartClk[2]), 
            .Q(r_Bit_Index[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i0.GSR = "ENABLED";
    LUT4 i8351_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n19820), .C(n18566), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_13)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(69[7] 161[14])
    defparam i8351_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i8346_3_lut_4_lut (.A(r_SM_Main[0]), .B(n19820), .C(r_Bit_Index[1]), 
         .D(n18566), .Z(UartClk_2_enable_15)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(69[7] 161[14])
    defparam i8346_3_lut_4_lut.init = 16'h0010;
    FD1P3IX r_Clock_Count_3041__i6 (.D(n69[6]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i6.GSR = "ENABLED";
    LUT4 i8343_3_lut_4_lut (.A(r_SM_Main[0]), .B(n19820), .C(r_Bit_Index[2]), 
         .D(n18579), .Z(UartClk_2_enable_16)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(69[7] 161[14])
    defparam i8343_3_lut_4_lut.init = 16'h1000;
    LUT4 i8376_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(r_SM_Main_2__N_2965[0]), 
         .D(n18732), .Z(UartClk_2_enable_34)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(69[7] 161[14])
    defparam i8376_4_lut.init = 16'h5455;
    LUT4 i1_2_lut (.A(r_Rx_Data), .B(r_SM_Main[0]), .Z(n18732)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(r_SM_Main[2]), .B(n24), .C(n19821), .D(r_SM_Main[1]), 
         .Z(n14275)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i1_4_lut.init = 16'h5044;
    LUT4 i1_4_lut_adj_225 (.A(r_Rx_Data), .B(r_SM_Main[0]), .C(n17972), 
         .D(n18744), .Z(n24)) /* synthesis lut_function=(!(A (B)+!A (B (C+!(D))))) */ ;
    defparam i1_4_lut_adj_225.init = 16'h3733;
    FD1P3IX r_Clock_Count_3041__i5 (.D(n69[5]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i5.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_3041__i4 (.D(n69[4]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i4.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(r_Clock_Count[5]), .B(r_Clock_Count[3]), .C(r_Clock_Count[0]), 
         .Z(n18744)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_226 (.A(r_Clock_Count[1]), .B(n18528), .C(n18736), 
         .D(r_Clock_Count[6]), .Z(n17972)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(85[17:52])
    defparam i1_4_lut_adj_226.init = 16'hfffd;
    LUT4 i1_2_lut_adj_227 (.A(r_Clock_Count[2]), .B(r_Clock_Count[4]), .Z(n18736)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_227.init = 16'heeee;
    LUT4 i1_4_lut_adj_228 (.A(n26), .B(n19821), .C(r_SM_Main[0]), .D(r_SM_Main[1]), 
         .Z(n18623)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_228.init = 16'h0800;
    LUT4 i39_2_lut (.A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .Z(n26)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i39_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_229 (.A(n18714), .B(n18716), .C(n18708), .D(n18712), 
         .Z(n18528)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(85[17:52])
    defparam i1_4_lut_adj_229.init = 16'hfffe;
    LUT4 i1_2_lut_adj_230 (.A(r_Clock_Count[11]), .B(r_Clock_Count[15]), 
         .Z(n18714)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_230.init = 16'heeee;
    LUT4 i1_3_lut_adj_231 (.A(r_Clock_Count[13]), .B(r_Clock_Count[8]), 
         .C(r_Clock_Count[7]), .Z(n18716)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(85[17:52])
    defparam i1_3_lut_adj_231.init = 16'hfefe;
    LUT4 i1_2_lut_adj_232 (.A(r_Clock_Count[14]), .B(r_Clock_Count[10]), 
         .Z(n18708)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_232.init = 16'heeee;
    LUT4 i1_2_lut_adj_233 (.A(r_Clock_Count[9]), .B(r_Clock_Count[12]), 
         .Z(n18712)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_233.init = 16'heeee;
    LUT4 i5127_4_lut (.A(n14677), .B(r_Clock_Count[6]), .C(r_Clock_Count[5]), 
         .D(r_Clock_Count[4]), .Z(n14691)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i5127_4_lut.init = 16'hc8c0;
    LUT4 i5113_3_lut (.A(r_Clock_Count[1]), .B(r_Clock_Count[3]), .C(r_Clock_Count[2]), 
         .Z(n14677)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i5113_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_234 (.A(r_Clock_Count[3]), .B(n17972), .C(r_Clock_Count[5]), 
         .D(r_Clock_Count[0]), .Z(r_SM_Main_2__N_2965[0])) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;
    defparam i1_4_lut_adj_234.init = 16'hdfff;
    LUT4 i8353_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n19820), .C(n18579), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_4)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(69[7] 161[14])
    defparam i8353_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 r_SM_Main_2__N_2959_2__bdd_3_lut (.A(r_SM_Main_2__N_2965[0]), .B(r_Rx_Data), 
         .C(r_SM_Main[0]), .Z(n19414)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+(C))) */ ;
    defparam r_SM_Main_2__N_2959_2__bdd_3_lut.init = 16'ha3a3;
    FD1P3IX r_Clock_Count_3041__i3 (.D(n69[3]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i3.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i1 (.D(n19849), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i1.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut (.A(n14691), .B(n18528), .C(n14667), .D(n18750), 
         .Z(n18685)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0e00;
    LUT4 i8373_4_lut (.A(n18528), .B(n18560), .C(n14691), .D(r_SM_Main[1]), 
         .Z(UartClk_2_enable_36)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i8373_4_lut.init = 16'h3233;
    LUT4 i1_4_lut_adj_235 (.A(r_Bit_Index[2]), .B(r_SM_Main[0]), .C(n18579), 
         .D(r_SM_Main[1]), .Z(n18750)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_235.init = 16'h1200;
    LUT4 i7447_2_lut (.A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .Z(n18579)) /* synthesis lut_function=(A (B)) */ ;
    defparam i7447_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_236 (.A(r_SM_Main[0]), .B(r_SM_Main[2]), .Z(n18560)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_236.init = 16'heeee;
    LUT4 i1_3_lut_adj_237 (.A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .C(r_Bit_Index[2]), 
         .Z(n14667)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_237.init = 16'h8080;
    LUT4 i1_2_lut_adj_238 (.A(r_Bit_Index[0]), .B(r_Bit_Index[2]), .Z(n18566)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(114[17:39])
    defparam i1_2_lut_adj_238.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_278_4_lut (.A(r_SM_Main[1]), .B(n19821), .C(r_SM_Main[2]), 
         .D(r_SM_Main[0]), .Z(n19817)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_278_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_adj_239 (.A(r_Bit_Index[0]), .B(r_SM_Main[1]), .Z(n18523)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_239.init = 16'h4444;
    FD1S3AX UartClk_3039_3066__i0 (.D(n17[0]), .CK(clk_80mhz), .Q(n30[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_3039_3066__i0.GSR = "ENABLED";
    LUT4 i8363_2_lut_4_lut (.A(r_SM_Main[1]), .B(n19821), .C(r_SM_Main[2]), 
         .D(r_SM_Main[0]), .Z(UartClk_2_enable_17)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i8363_2_lut_4_lut.init = 16'h0800;
    LUT4 i1_2_lut_rep_282 (.A(n14691), .B(n18528), .Z(n19821)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_282.init = 16'heeee;
    LUT4 r_SM_Main_2__N_2959_2__bdd_3_lut_8433_4_lut (.A(n14691), .B(n18528), 
         .C(r_SM_Main[0]), .D(n14667), .Z(n19413)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam r_SM_Main_2__N_2959_2__bdd_3_lut_8433_4_lut.init = 16'h1e10;
    LUT4 i1_3_lut_rep_281_4_lut (.A(n14691), .B(n18528), .C(r_SM_Main[2]), 
         .D(r_SM_Main[1]), .Z(n19820)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;
    defparam i1_3_lut_rep_281_4_lut.init = 16'hf1ff;
    LUT4 i8389_3_lut_3_lut_4_lut (.A(n14691), .B(n18528), .C(n18560), 
         .D(r_SM_Main[1]), .Z(UartClk_2_enable_19)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+(D))))) */ ;
    defparam i8389_3_lut_3_lut_4_lut.init = 16'h0e0f;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut (.A(r_SM_Main[0]), 
         .B(n18528), .C(n14691), .Z(n19848)) /* synthesis lut_function=(!(A (B+(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(69[7] 161[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut.init = 16'h5757;
    FD1P3IX r_Clock_Count_3041__i2 (.D(n69[2]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i2.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_3041__i1 (.D(n69[1]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i1.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i2 (.D(n19821), .CK(UartClk[2]), .CD(n18550), .Q(r_SM_Main[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i2.GSR = "ENABLED";
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut (.A(r_SM_Main[0]), 
         .B(r_SM_Main_2__N_2965[0]), .C(r_Rx_Data), .Z(n19847)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(69[7] 161[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut.init = 16'h0202;
    FD1S3AX UartClk_3039_3066__i1 (.D(n17[1]), .CK(clk_80mhz), .Q(n30[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_3039_3066__i1.GSR = "ENABLED";
    FD1S3AX UartClk_3039_3066__i2 (.D(n17[2]), .CK(clk_80mhz), .Q(UartClk[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_3039_3066__i2.GSR = "ENABLED";
    CCU2C r_Clock_Count_3041_add_4_17 (.A0(r_Clock_Count[15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17064), .S0(n69[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041_add_4_17.INIT0 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_17.INIT1 = 16'h0000;
    defparam r_Clock_Count_3041_add_4_17.INJECT1_0 = "NO";
    defparam r_Clock_Count_3041_add_4_17.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_3041_add_4_15 (.A0(r_Clock_Count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17063), .COUT(n17064), .S0(n69[13]), 
          .S1(n69[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041_add_4_15.INIT0 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_15.INIT1 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_15.INJECT1_0 = "NO";
    defparam r_Clock_Count_3041_add_4_15.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_3041_add_4_13 (.A0(r_Clock_Count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17062), .COUT(n17063), .S0(n69[11]), 
          .S1(n69[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041_add_4_13.INIT0 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_13.INIT1 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_13.INJECT1_0 = "NO";
    defparam r_Clock_Count_3041_add_4_13.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_3041_add_4_11 (.A0(r_Clock_Count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17061), .COUT(n17062), .S0(n69[9]), 
          .S1(n69[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041_add_4_11.INIT0 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_11.INIT1 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_11.INJECT1_0 = "NO";
    defparam r_Clock_Count_3041_add_4_11.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_3041_add_4_9 (.A0(r_Clock_Count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17060), .COUT(n17061), .S0(n69[7]), 
          .S1(n69[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041_add_4_9.INIT0 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_9.INIT1 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_9.INJECT1_0 = "NO";
    defparam r_Clock_Count_3041_add_4_9.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_3041_add_4_7 (.A0(r_Clock_Count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17059), .COUT(n17060), .S0(n69[5]), 
          .S1(n69[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041_add_4_7.INIT0 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_7.INIT1 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_7.INJECT1_0 = "NO";
    defparam r_Clock_Count_3041_add_4_7.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_3041_add_4_5 (.A0(r_Clock_Count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17058), .COUT(n17059), .S0(n69[3]), 
          .S1(n69[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041_add_4_5.INIT0 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_5.INIT1 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_5.INJECT1_0 = "NO";
    defparam r_Clock_Count_3041_add_4_5.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_3041_add_4_3 (.A0(r_Clock_Count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n17057), .COUT(n17058), .S0(n69[1]), 
          .S1(n69[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041_add_4_3.INIT0 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_3.INIT1 = 16'haaa0;
    defparam r_Clock_Count_3041_add_4_3.INJECT1_0 = "NO";
    defparam r_Clock_Count_3041_add_4_3.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_3041_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(r_Clock_Count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n17057), .S1(n69[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041_add_4_1.INIT0 = 16'h0000;
    defparam r_Clock_Count_3041_add_4_1.INIT1 = 16'h555f;
    defparam r_Clock_Count_3041_add_4_1.INJECT1_0 = "NO";
    defparam r_Clock_Count_3041_add_4_1.INJECT1_1 = "NO";
    LUT4 i8348_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n19817), .C(r_Bit_Index[2]), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_14)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(114[17:39])
    defparam i8348_2_lut_3_lut_4_lut.init = 16'h1000;
    PFUMX i8434 (.BLUT(n19414), .ALUT(n19413), .C0(r_SM_Main[1]), .Z(n19415));
    LUT4 i1_2_lut_rep_290 (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .Z(n19829)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(69[7] 161[14])
    defparam i1_2_lut_rep_290.init = 16'h2222;
    LUT4 i8366_2_lut_3_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .Z(n18550)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(69[7] 161[14])
    defparam i8366_2_lut_3_lut.init = 16'hdfdf;
    LUT4 i8358_2_lut_3_lut_4_lut (.A(r_Bit_Index[1]), .B(n19817), .C(r_Bit_Index[2]), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_35)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(114[17:39])
    defparam i8358_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i21_4_lut_4_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .D(n19821), .Z(UartClk_2_enable_29)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(69[7] 161[14])
    defparam i21_4_lut_4_lut.init = 16'h2505;
    LUT4 i8361_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n19817), .C(r_Bit_Index[1]), 
         .D(r_Bit_Index[0]), .Z(UartClk_2_enable_28)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(114[17:39])
    defparam i8361_2_lut_3_lut_4_lut.init = 16'h0001;
    FD1P3IX r_Clock_Count_3041__i0 (.D(n69[0]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i0.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_3041__i14 (.D(n69[14]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[14])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i14.GSR = "ENABLED";
    FD1S3IX o_Rx_DV_59 (.D(r_Rx_DV_last_N_3024), .CK(clk_80mhz), .CD(n14269), 
            .Q(rx_data_valid1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(47[11] 52[8])
    defparam o_Rx_DV_59.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i0 (.D(r_Rx_Data), .SP(UartClk_2_enable_28), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i0.GSR = "ENABLED";
    FD1P3AX r_Rx_DV_64 (.D(r_Rx_DV_N_3025), .SP(UartClk_2_enable_29), .CK(UartClk[2]), 
            .Q(r_Rx_DV)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_DV_64.GSR = "ENABLED";
    PFUMX i8757 (.BLUT(n19847), .ALUT(n19848), .C0(r_SM_Main[1]), .Z(n19849));
    FD1P3IX r_Clock_Count_3041__i15 (.D(n69[15]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[15])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i15.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_3041__i12 (.D(n69[12]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[12])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i12.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_3041__i13 (.D(n69[13]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[13])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i13.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_3041__i10 (.D(n69[10]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[10])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i10.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_3041__i11 (.D(n69[11]), .SP(UartClk_2_enable_34), 
            .CD(n14275), .CK(UartClk[2]), .Q(r_Clock_Count[11])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_3041__i11.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n14691), .B(n18528), .C(n19829), .D(r_SM_Main[0]), 
         .Z(r_Rx_DV_N_3025)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'he000;
    FD1P3AX r_Rx_Byte_i1 (.D(r_Rx_Data), .SP(UartClk_2_enable_35), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i1.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i1 (.D(n18623), .SP(UartClk_2_enable_36), .CK(UartClk[2]), 
            .Q(r_Bit_Index[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=5, LSE_LLINE=245, LSE_RLINE=250 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i1.GSR = "ENABLED";
    CCU2C UartClk_3039_3066_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n17892), .S1(n17[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_3039_3066_add_4_1.INIT0 = 16'h0000;
    defparam UartClk_3039_3066_add_4_1.INIT1 = 16'h555f;
    defparam UartClk_3039_3066_add_4_1.INJECT1_0 = "NO";
    defparam UartClk_3039_3066_add_4_1.INJECT1_1 = "NO";
    CCU2C UartClk_3039_3066_add_4_3 (.A0(n30[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(UartClk[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n17892), .S0(n17[1]), .S1(n17[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_3039_3066_add_4_3.INIT0 = 16'haaa0;
    defparam UartClk_3039_3066_add_4_3.INIT1 = 16'haaa0;
    defparam UartClk_3039_3066_add_4_3.INJECT1_0 = "NO";
    defparam UartClk_3039_3066_add_4_3.INJECT1_1 = "NO";
    LUT4 i4706_1_lut (.A(r_Rx_DV), .Z(n14269)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(66[10] 162[8])
    defparam i4706_1_lut.init = 16'h5555;
    LUT4 r_Rx_DV_last_I_0_1_lut (.A(r_Rx_DV_last), .Z(r_Rx_DV_last_N_3024)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/UartRX.v(50[30:43])
    defparam r_Rx_DV_last_I_0_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module PLL
//

module PLL (clk_25mhz_c, clk_80mhz, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk_25mhz_c;
    output clk_80mhz;
    input GND_net;
    
    wire clk_25mhz_c /* synthesis is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(38[22:31])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(61[34:43])
    
    wire CLKFB_t;
    
    EHXPLLL PLLInst_0 (.CLKI(clk_25mhz_c), .CLKFB(CLKFB_t), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .PHASELOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .CLKOP(clk_80mhz), .CLKINTFB(CLKFB_t)) /* synthesis FREQUENCY_PIN_CLKOP="83.333333", FREQUENCY_PIN_CLKI="25.000000", ICP_CURRENT="5", LPF_RESISTOR="16", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=96, LSE_RLINE=99 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(96[8] 99[5])
    defparam PLLInst_0.CLKI_DIV = 3;
    defparam PLLInst_0.CLKFB_DIV = 10;
    defparam PLLInst_0.CLKOP_DIV = 7;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 6;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "INT_OP";
    defparam PLLInst_0.CLKOP_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.PLL_LOCK_DELAY = 200;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.REFIN_RESET = "DISABLED";
    defparam PLLInst_0.SYNC_ENABLE = "DISABLED";
    defparam PLLInst_0.INT_LOCK_STICKY = "ENABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AMDemodulator
//

module AMDemodulator (cic_sine_clk, led_0_2, led_0_1, n51, n51_adj_229, 
            n19813, \amdemod_out_d_11__N_2379[14] , \amdemod_out_d_11__N_2380[14] , 
            n19815, led_0_0, \cic_sine_out[5] , n19816, \cic_sine_out[4] , 
            \cic_sine_out[3] , \cic_sine_out[2] , \cic_sine_out[1] , \data_in_reg_11__N_2898[7] , 
            n46, n46_adj_230, n48, n48_adj_231, n43, n43_adj_232, 
            n45, n45_adj_233, n40, n40_adj_234, n42, n42_adj_235, 
            cic_cosine_out, \data_in_reg_11__N_2898[6] , n76, n76_adj_236, 
            n19811, \data_in_reg_11__N_2898[5] , \data_in_reg_11__N_2898[4] , 
            \data_in_reg_11__N_2898[3] , \data_in_reg_11__N_2898[2] , \data_in_reg_11__N_2898[1] , 
            n78, n78_adj_237, n73, n73_adj_238, n75, n75_adj_239, 
            \cic_sine_out[0] , n70, n70_adj_240, n72, n72_adj_241, 
            n67, n67_adj_242, n69, n69_adj_243, n64, n64_adj_244, 
            n66, n66_adj_245, \data_in_reg_11__N_2898[0] , n61, n61_adj_246, 
            n63, n63_adj_247, led_0_4, led_0_5, n58, n58_adj_248, 
            n36, n36_adj_249, amdemod_out_d_11__N_2363, n60, n60_adj_250, 
            n34, n34_adj_251, n55, n55_adj_252, n57, n57_adj_253, 
            n52, n52_adj_254, n54, n54_adj_255, n36_adj_256, n36_adj_257, 
            n49, n49_adj_258, n34_adj_259, n34_adj_260, n51_adj_261, 
            n51_adj_262, n46_adj_263, n46_adj_264, n48_adj_265, n48_adj_266, 
            n43_adj_267, n43_adj_268, n45_adj_269, n45_adj_270, n40_adj_271, 
            n40_adj_272, n42_adj_273, n42_adj_274, n76_adj_275, n76_adj_276, 
            n36_adj_277, n36_adj_278, n78_adj_279, n78_adj_280, n34_adj_281, 
            n34_adj_282, n36_adj_283, n36_adj_284, n34_adj_285, n34_adj_286, 
            \square_sum[23] , \square_sum[22] , n4, n34_adj_287, n34_adj_288, 
            n19809, \amdemod_out_d_11__N_2369[11] , \amdemod_out_d_11__N_2370[11] , 
            n36_adj_289, n36_adj_290, n13878, n42_adj_291, \square_sum[25] , 
            amdemod_out_d_11__N_2516, n64_adj_292, n64_adj_293, n66_adj_294, 
            n66_adj_295, n67_adj_296, n67_adj_297, n69_adj_298, n69_adj_299, 
            n58_adj_300, n58_adj_301, n60_adj_302, n60_adj_303, n61_adj_304, 
            n61_adj_305, amdemod_out_d_11__N_2594, n63_adj_306, n63_adj_307, 
            n55_adj_308, n55_adj_309, n57_adj_310, n57_adj_311, n52_adj_312, 
            n52_adj_313, n54_adj_314, n54_adj_315, \amdemod_out[9] , 
            \data_in_reg_11__N_2898[8] , n39, \amdemod_out_d_11__N_2365[3] , 
            n39_adj_316, n49_adj_317, n49_adj_318, n51_adj_319, n51_adj_320, 
            n46_adj_321, n46_adj_322, n48_adj_323, n48_adj_324, n19810, 
            n19828, n19827, \amdemod_out_d_11__N_2365[14] , n24, n13890, 
            n43_adj_325, n43_adj_326, n45_adj_327, n45_adj_328, n40_adj_329, 
            n40_adj_330, n30, n76_adj_331, n76_adj_332, n78_adj_333, 
            n78_adj_334, n42_adj_335, n42_adj_336, \amdemod_out_d_11__N_2409[14] , 
            \amdemod_out_d_11__N_2410[14] , n19808, \amdemod_out_d_11__N_2365[1] , 
            n45_adj_337, n13876, \amdemod_out_d_11__N_2365[6] , n30_adj_338, 
            \amdemod_out_d_11__N_2365[2] , n42_adj_339, amdemod_out_d_11__N_2597, 
            n73_adj_340, n73_adj_341, n75_adj_342, n75_adj_343, n70_adj_344, 
            n70_adj_345, n73_adj_346, n73_adj_347, n75_adj_348, n75_adj_349, 
            n70_adj_350, n70_adj_351, n72_adj_352, n72_adj_353, n72_adj_354, 
            n72_adj_355, n67_adj_356, n67_adj_357, \amdemod_out_d_11__N_2358[5] , 
            n33, n69_adj_358, n69_adj_359, n64_adj_360, n64_adj_361, 
            \amdemod_out_d_11__N_2365[4] , n36_adj_362, \amdemod_out_d_11__N_2365[5] , 
            n33_adj_363, n66_adj_364, n66_adj_365, n36_adj_366, n61_adj_367, 
            n61_adj_368, n63_adj_369, n63_adj_370, n58_adj_371, n58_adj_372, 
            n60_adj_373, n60_adj_374, n55_adj_375, n55_adj_376, n57_adj_377, 
            n57_adj_378, n52_adj_379, n52_adj_380, n54_adj_381, n54_adj_382, 
            n49_adj_383, n49_adj_384, n51_adj_385, n51_adj_386, \amdemod_out_d_11__N_2365[7] , 
            n27, amdemod_out_d_11__N_2564, n46_adj_387, n46_adj_388, 
            n48_adj_389, n48_adj_390, amdemod_out_d_11__N_2567, n46_adj_391, 
            n48_adj_392, n13821, n13815, n43_adj_393, n43_adj_394, 
            amdemod_out_d_11__N_2570, \amdemod_out_d_11__N_2399[14] , \amdemod_out_d_11__N_2400[14] , 
            amdemod_out_d_11__N_2573, n45_adj_395, n45_adj_396, n40_adj_397, 
            n40_adj_398, n42_adj_399, n42_adj_400, amdemod_out_d_11__N_2576, 
            n76_adj_401, n76_adj_402, n19812, amdemod_out_d_11__N_2579, 
            n78_adj_403, n78_adj_404, n73_adj_405, n73_adj_406, \amdemod_out_d_11__N_2389[14] , 
            \amdemod_out_d_11__N_2390[14] , n75_adj_407, n75_adj_408, 
            n70_adj_409, n70_adj_410, amdemod_out_d_11__N_2585, n72_adj_411, 
            n72_adj_412, n67_adj_413, n67_adj_414, amdemod_out_d_11__N_2582, 
            n69_adj_415, n69_adj_416, n19824, n64_adj_417, n64_adj_418, 
            n66_adj_419, n66_adj_420, n61_adj_421, n61_adj_422, n63_adj_423, 
            n63_adj_424, n58_adj_425, n58_adj_426, n60_adj_427, n60_adj_428, 
            n19814, n55_adj_429, n55_adj_430, n57_adj_431, n57_adj_432, 
            amdemod_out_d_11__N_2591, n52_adj_433, n52_adj_434, amdemod_out_d_11__N_2588, 
            n54_adj_435, n54_adj_436, n49_adj_437, n49_adj_438, amdemod_out_d_11__N_2600, 
            amdemod_out_d_11__N_2798, amdemod_out_d_11__N_2801, amdemod_out_d_11__N_2804, 
            amdemod_out_d_11__N_2807, amdemod_out_d_11__N_2810, amdemod_out_d_11__N_2813, 
            amdemod_out_d_11__N_2816, amdemod_out_d_11__N_2819, amdemod_out_d_11__N_2822, 
            amdemod_out_d_11__N_2825, amdemod_out_d_11__N_2828, amdemod_out_d_11__N_2831, 
            amdemod_out_d_11__N_2834, amdemod_out_d_11__N_2720, amdemod_out_d_11__N_2723, 
            amdemod_out_d_11__N_2726, amdemod_out_d_11__N_2729, amdemod_out_d_11__N_2732, 
            amdemod_out_d_11__N_2735, amdemod_out_d_11__N_2738, amdemod_out_d_11__N_2741, 
            amdemod_out_d_11__N_2744, amdemod_out_d_11__N_2747, amdemod_out_d_11__N_2750, 
            amdemod_out_d_11__N_2753, amdemod_out_d_11__N_2756, led_0_3, 
            amdemod_out_d_11__N_2642, amdemod_out_d_11__N_2645, amdemod_out_d_11__N_2648, 
            amdemod_out_d_11__N_2501, amdemod_out_d_11__N_2651, amdemod_out_d_11__N_2654, 
            amdemod_out_d_11__N_2657, amdemod_out_d_11__N_2507, amdemod_out_d_11__N_2660, 
            amdemod_out_d_11__N_2663, amdemod_out_d_11__N_2666, amdemod_out_d_11__N_2669, 
            amdemod_out_d_11__N_2504, amdemod_out_d_11__N_2672, amdemod_out_d_11__N_2675, 
            amdemod_out_d_11__N_2678, amdemod_out_d_11__N_2513, amdemod_out_d_11__N_2510, 
            VCC_net, GND_net, q_squared, i_squared) /* synthesis syn_module_defined=1 */ ;
    input cic_sine_clk;
    input led_0_2;
    input led_0_1;
    input n51;
    input n51_adj_229;
    output n19813;
    input \amdemod_out_d_11__N_2379[14] ;
    input \amdemod_out_d_11__N_2380[14] ;
    output n19815;
    input led_0_0;
    input \cic_sine_out[5] ;
    output n19816;
    input \cic_sine_out[4] ;
    input \cic_sine_out[3] ;
    input \cic_sine_out[2] ;
    input \cic_sine_out[1] ;
    output \data_in_reg_11__N_2898[7] ;
    input n46;
    input n46_adj_230;
    input n48;
    input n48_adj_231;
    input n43;
    input n43_adj_232;
    input n45;
    input n45_adj_233;
    input n40;
    input n40_adj_234;
    input n42;
    input n42_adj_235;
    input [11:0]cic_cosine_out;
    output \data_in_reg_11__N_2898[6] ;
    input n76;
    input n76_adj_236;
    output n19811;
    output \data_in_reg_11__N_2898[5] ;
    output \data_in_reg_11__N_2898[4] ;
    output \data_in_reg_11__N_2898[3] ;
    output \data_in_reg_11__N_2898[2] ;
    output \data_in_reg_11__N_2898[1] ;
    input n78;
    input n78_adj_237;
    input n73;
    input n73_adj_238;
    input n75;
    input n75_adj_239;
    input \cic_sine_out[0] ;
    input n70;
    input n70_adj_240;
    input n72;
    input n72_adj_241;
    input n67;
    input n67_adj_242;
    input n69;
    input n69_adj_243;
    input n64;
    input n64_adj_244;
    input n66;
    input n66_adj_245;
    output \data_in_reg_11__N_2898[0] ;
    input n61;
    input n61_adj_246;
    input n63;
    input n63_adj_247;
    input led_0_4;
    input led_0_5;
    input n58;
    input n58_adj_248;
    input n36;
    input n36_adj_249;
    output amdemod_out_d_11__N_2363;
    input n60;
    input n60_adj_250;
    input n34;
    input n34_adj_251;
    input n55;
    input n55_adj_252;
    input n57;
    input n57_adj_253;
    input n52;
    input n52_adj_254;
    input n54;
    input n54_adj_255;
    input n36_adj_256;
    input n36_adj_257;
    input n49;
    input n49_adj_258;
    input n34_adj_259;
    input n34_adj_260;
    input n51_adj_261;
    input n51_adj_262;
    input n46_adj_263;
    input n46_adj_264;
    input n48_adj_265;
    input n48_adj_266;
    input n43_adj_267;
    input n43_adj_268;
    input n45_adj_269;
    input n45_adj_270;
    input n40_adj_271;
    input n40_adj_272;
    input n42_adj_273;
    input n42_adj_274;
    input n76_adj_275;
    input n76_adj_276;
    input n36_adj_277;
    input n36_adj_278;
    input n78_adj_279;
    input n78_adj_280;
    input n34_adj_281;
    input n34_adj_282;
    input n36_adj_283;
    input n36_adj_284;
    input n34_adj_285;
    input n34_adj_286;
    input \square_sum[23] ;
    input \square_sum[22] ;
    output n4;
    input n34_adj_287;
    input n34_adj_288;
    output n19809;
    input \amdemod_out_d_11__N_2369[11] ;
    input \amdemod_out_d_11__N_2370[11] ;
    input n36_adj_289;
    input n36_adj_290;
    output n13878;
    input n42_adj_291;
    input \square_sum[25] ;
    output amdemod_out_d_11__N_2516;
    input n64_adj_292;
    input n64_adj_293;
    input n66_adj_294;
    input n66_adj_295;
    input n67_adj_296;
    input n67_adj_297;
    input n69_adj_298;
    input n69_adj_299;
    input n58_adj_300;
    input n58_adj_301;
    input n60_adj_302;
    input n60_adj_303;
    input n61_adj_304;
    input n61_adj_305;
    output amdemod_out_d_11__N_2594;
    input n63_adj_306;
    input n63_adj_307;
    input n55_adj_308;
    input n55_adj_309;
    input n57_adj_310;
    input n57_adj_311;
    input n52_adj_312;
    input n52_adj_313;
    input n54_adj_314;
    input n54_adj_315;
    output \amdemod_out[9] ;
    output \data_in_reg_11__N_2898[8] ;
    input n39;
    input \amdemod_out_d_11__N_2365[3] ;
    input n39_adj_316;
    input n49_adj_317;
    input n49_adj_318;
    input n51_adj_319;
    input n51_adj_320;
    input n46_adj_321;
    input n46_adj_322;
    input n48_adj_323;
    input n48_adj_324;
    output n19810;
    output n19828;
    output n19827;
    input \amdemod_out_d_11__N_2365[14] ;
    input n24;
    output n13890;
    input n43_adj_325;
    input n43_adj_326;
    input n45_adj_327;
    input n45_adj_328;
    input n40_adj_329;
    input n40_adj_330;
    input n30;
    input n76_adj_331;
    input n76_adj_332;
    input n78_adj_333;
    input n78_adj_334;
    input n42_adj_335;
    input n42_adj_336;
    input \amdemod_out_d_11__N_2409[14] ;
    input \amdemod_out_d_11__N_2410[14] ;
    output n19808;
    input \amdemod_out_d_11__N_2365[1] ;
    input n45_adj_337;
    output n13876;
    input \amdemod_out_d_11__N_2365[6] ;
    input n30_adj_338;
    input \amdemod_out_d_11__N_2365[2] ;
    input n42_adj_339;
    output amdemod_out_d_11__N_2597;
    input n73_adj_340;
    input n73_adj_341;
    input n75_adj_342;
    input n75_adj_343;
    input n70_adj_344;
    input n70_adj_345;
    input n73_adj_346;
    input n73_adj_347;
    input n75_adj_348;
    input n75_adj_349;
    input n70_adj_350;
    input n70_adj_351;
    input n72_adj_352;
    input n72_adj_353;
    input n72_adj_354;
    input n72_adj_355;
    input n67_adj_356;
    input n67_adj_357;
    output \amdemod_out_d_11__N_2358[5] ;
    input n33;
    input n69_adj_358;
    input n69_adj_359;
    input n64_adj_360;
    input n64_adj_361;
    input \amdemod_out_d_11__N_2365[4] ;
    input n36_adj_362;
    input \amdemod_out_d_11__N_2365[5] ;
    input n33_adj_363;
    input n66_adj_364;
    input n66_adj_365;
    input n36_adj_366;
    input n61_adj_367;
    input n61_adj_368;
    input n63_adj_369;
    input n63_adj_370;
    input n58_adj_371;
    input n58_adj_372;
    input n60_adj_373;
    input n60_adj_374;
    input n55_adj_375;
    input n55_adj_376;
    input n57_adj_377;
    input n57_adj_378;
    input n52_adj_379;
    input n52_adj_380;
    input n54_adj_381;
    input n54_adj_382;
    input n49_adj_383;
    input n49_adj_384;
    input n51_adj_385;
    input n51_adj_386;
    input \amdemod_out_d_11__N_2365[7] ;
    input n27;
    output amdemod_out_d_11__N_2564;
    input n46_adj_387;
    input n46_adj_388;
    input n48_adj_389;
    input n48_adj_390;
    output amdemod_out_d_11__N_2567;
    input n46_adj_391;
    input n48_adj_392;
    output n13821;
    output n13815;
    input n43_adj_393;
    input n43_adj_394;
    output amdemod_out_d_11__N_2570;
    input \amdemod_out_d_11__N_2399[14] ;
    input \amdemod_out_d_11__N_2400[14] ;
    output amdemod_out_d_11__N_2573;
    input n45_adj_395;
    input n45_adj_396;
    input n40_adj_397;
    input n40_adj_398;
    input n42_adj_399;
    input n42_adj_400;
    output amdemod_out_d_11__N_2576;
    input n76_adj_401;
    input n76_adj_402;
    output n19812;
    output amdemod_out_d_11__N_2579;
    input n78_adj_403;
    input n78_adj_404;
    input n73_adj_405;
    input n73_adj_406;
    input \amdemod_out_d_11__N_2389[14] ;
    input \amdemod_out_d_11__N_2390[14] ;
    input n75_adj_407;
    input n75_adj_408;
    input n70_adj_409;
    input n70_adj_410;
    output amdemod_out_d_11__N_2585;
    input n72_adj_411;
    input n72_adj_412;
    input n67_adj_413;
    input n67_adj_414;
    output amdemod_out_d_11__N_2582;
    input n69_adj_415;
    input n69_adj_416;
    output n19824;
    input n64_adj_417;
    input n64_adj_418;
    input n66_adj_419;
    input n66_adj_420;
    input n61_adj_421;
    input n61_adj_422;
    input n63_adj_423;
    input n63_adj_424;
    input n58_adj_425;
    input n58_adj_426;
    input n60_adj_427;
    input n60_adj_428;
    output n19814;
    input n55_adj_429;
    input n55_adj_430;
    input n57_adj_431;
    input n57_adj_432;
    output amdemod_out_d_11__N_2591;
    input n52_adj_433;
    input n52_adj_434;
    output amdemod_out_d_11__N_2588;
    input n54_adj_435;
    input n54_adj_436;
    input n49_adj_437;
    input n49_adj_438;
    output amdemod_out_d_11__N_2600;
    output amdemod_out_d_11__N_2798;
    output amdemod_out_d_11__N_2801;
    output amdemod_out_d_11__N_2804;
    output amdemod_out_d_11__N_2807;
    output amdemod_out_d_11__N_2810;
    output amdemod_out_d_11__N_2813;
    output amdemod_out_d_11__N_2816;
    output amdemod_out_d_11__N_2819;
    output amdemod_out_d_11__N_2822;
    output amdemod_out_d_11__N_2825;
    output amdemod_out_d_11__N_2828;
    output amdemod_out_d_11__N_2831;
    output amdemod_out_d_11__N_2834;
    output amdemod_out_d_11__N_2720;
    output amdemod_out_d_11__N_2723;
    output amdemod_out_d_11__N_2726;
    output amdemod_out_d_11__N_2729;
    output amdemod_out_d_11__N_2732;
    output amdemod_out_d_11__N_2735;
    output amdemod_out_d_11__N_2738;
    output amdemod_out_d_11__N_2741;
    output amdemod_out_d_11__N_2744;
    output amdemod_out_d_11__N_2747;
    output amdemod_out_d_11__N_2750;
    output amdemod_out_d_11__N_2753;
    output amdemod_out_d_11__N_2756;
    input led_0_3;
    output amdemod_out_d_11__N_2642;
    output amdemod_out_d_11__N_2645;
    output amdemod_out_d_11__N_2648;
    output amdemod_out_d_11__N_2501;
    output amdemod_out_d_11__N_2651;
    output amdemod_out_d_11__N_2654;
    output amdemod_out_d_11__N_2657;
    output amdemod_out_d_11__N_2507;
    output amdemod_out_d_11__N_2660;
    output amdemod_out_d_11__N_2663;
    output amdemod_out_d_11__N_2666;
    output amdemod_out_d_11__N_2669;
    output amdemod_out_d_11__N_2504;
    output amdemod_out_d_11__N_2672;
    output amdemod_out_d_11__N_2675;
    output amdemod_out_d_11__N_2678;
    output amdemod_out_d_11__N_2513;
    output amdemod_out_d_11__N_2510;
    input VCC_net;
    input GND_net;
    output [23:0]q_squared;
    output [23:0]i_squared;
    
    wire cic_sine_clk /* synthesis SET_AS_NETWORK=cic_sine_clk, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(78[33:45])
    wire [11:0]i_data_b;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(21[34:42])
    
    wire n18938, amdemod_out_d_11__N_2377, n18899, n18900;
    wire [15:0]amdemod_out_d;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(17[21:34])
    
    wire amdemod_out_d_11__N_2372, n18936, n18935, n18933, n18932, 
        n18930, n18929;
    wire [11:0]q_data_a;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(25[34:42])
    
    wire n18924, n18923, n18921, n18920, n18918, n18917, n18915, 
        n18914, n18912, n18911, n18909, n18908, n18906, n18905, 
        n18897, n18896, n18891, n18890, n19016, n18879, n19017, 
        n18878, n18876, n18875, n18873, n18872, n18870, n18869, 
        n18894, n18971, n18893, n18972, n18926, n18927, n19312, 
        n19724, n19725, amdemod_out_d_11__N_2367, n19313, n19314, 
        n19023, n19022, n18882, n18881, n19041, n19303, n19040, 
        n18966, n19304, n18884, n18885, n18965, n19038, n19037, 
        n19035, n19034, n19836, n19835, n19032, n19031, n19029, 
        n19028, amdemod_out_d_11__N_2412, n19026, n19025, n19020, 
        n19839, n19014, n19013, n19019, amdemod_out_d_11__N_2402, 
        n19838, n18887, n18888, n19011, n19010, n19008, n19007, 
        n19005, n19842, n19004, n19002, n19832, n19841, n19001, 
        n19833, n18999, n18998, n18996, n18995, n18993, n18992, 
        n18990, n18989, n18987, n18986, n19845, n19844, n18984, 
        n18983, amdemod_out_d_11__N_2407, amdemod_out_d_11__N_2397, amdemod_out_d_11__N_2392, 
        amdemod_out_d_11__N_2387, amdemod_out_d_11__N_2382, n19305, n18981, 
        n18980, n18975, n18974, n18969, n19306, n18968, n19307, 
        n18963, n19308, n19309, n18962, n19310, n18960, n19311, 
        n18959, n18957, n18956, n18954, n18953, n18951, n18950, 
        n18948, n18947, n18945, n18944, n18942, n18941, n18939;
    
    FD1S3AX i_data_b_i8 (.D(led_0_2), .CK(cic_sine_clk), .Q(i_data_b[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam i_data_b_i8.GSR = "ENABLED";
    FD1S3AX i_data_b_i7 (.D(led_0_1), .CK(cic_sine_clk), .Q(i_data_b[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam i_data_b_i7.GSR = "ENABLED";
    LUT4 i7804_3_lut (.A(n51), .B(n51_adj_229), .C(n19813), .Z(n18938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7804_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_16_1_lut_3_lut (.A(\amdemod_out_d_11__N_2379[14] ), 
         .B(\amdemod_out_d_11__N_2380[14] ), .C(n19815), .Z(amdemod_out_d_11__N_2377)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_16_1_lut_3_lut.init = 16'h3535;
    FD1S3AX i_data_b_i6 (.D(led_0_0), .CK(cic_sine_clk), .Q(i_data_b[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam i_data_b_i6.GSR = "ENABLED";
    FD1S3AX i_data_b_i5 (.D(\cic_sine_out[5] ), .CK(cic_sine_clk), .Q(i_data_b[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam i_data_b_i5.GSR = "ENABLED";
    LUT4 i7767_3_lut_rep_276 (.A(n18899), .B(n18900), .C(n19816), .Z(n19815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7767_3_lut_rep_276.init = 16'hcaca;
    FD1S3AX i_data_b_i4 (.D(\cic_sine_out[4] ), .CK(cic_sine_clk), .Q(i_data_b[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam i_data_b_i4.GSR = "ENABLED";
    FD1S3AX i_data_b_i3 (.D(\cic_sine_out[3] ), .CK(cic_sine_clk), .Q(i_data_b[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam i_data_b_i3.GSR = "ENABLED";
    FD1S3AX i_data_b_i2 (.D(\cic_sine_out[2] ), .CK(cic_sine_clk), .Q(i_data_b[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam i_data_b_i2.GSR = "ENABLED";
    FD1S3AX i_data_b_i1 (.D(\cic_sine_out[1] ), .CK(cic_sine_clk), .Q(i_data_b[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam i_data_b_i1.GSR = "ENABLED";
    FD1S3AX amdemod_out_i8 (.D(amdemod_out_d[7]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2898[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_i8.GSR = "ENABLED";
    LUT4 amdemod_out_d_11__I_14_1_lut_3_lut (.A(n18899), .B(n18900), .C(n19816), 
         .Z(amdemod_out_d_11__N_2372)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam amdemod_out_d_11__I_14_1_lut_3_lut.init = 16'h3535;
    LUT4 i7802_3_lut (.A(n46), .B(n46_adj_230), .C(n19813), .Z(n18936)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7802_3_lut.init = 16'hcaca;
    LUT4 i7801_3_lut (.A(n48), .B(n48_adj_231), .C(n19813), .Z(n18935)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7801_3_lut.init = 16'hcaca;
    LUT4 i7799_3_lut (.A(n43), .B(n43_adj_232), .C(n19813), .Z(n18933)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7799_3_lut.init = 16'hcaca;
    LUT4 i7798_3_lut (.A(n45), .B(n45_adj_233), .C(n19813), .Z(n18932)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7798_3_lut.init = 16'hcaca;
    LUT4 i7796_3_lut (.A(n40), .B(n40_adj_234), .C(n19813), .Z(n18930)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7796_3_lut.init = 16'hcaca;
    LUT4 i7795_3_lut (.A(n42), .B(n42_adj_235), .C(n19813), .Z(n18929)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7795_3_lut.init = 16'hcaca;
    FD1S3AX q_data_a_i1 (.D(cic_cosine_out[1]), .CK(cic_sine_clk), .Q(q_data_a[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam q_data_a_i1.GSR = "ENABLED";
    FD1S3AX amdemod_out_i7 (.D(amdemod_out_d[6]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2898[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_i7.GSR = "ENABLED";
    LUT4 i7790_3_lut (.A(n76), .B(n76_adj_236), .C(n19811), .Z(n18924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7790_3_lut.init = 16'hcaca;
    FD1S3AX amdemod_out_i6 (.D(amdemod_out_d[5]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2898[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_i6.GSR = "ENABLED";
    FD1S3AX amdemod_out_i5 (.D(amdemod_out_d[4]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2898[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_i5.GSR = "ENABLED";
    FD1S3AX amdemod_out_i4 (.D(amdemod_out_d[3]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2898[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_i4.GSR = "ENABLED";
    FD1S3AX amdemod_out_i3 (.D(amdemod_out_d[2]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2898[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_i3.GSR = "ENABLED";
    FD1S3AX amdemod_out_i2 (.D(amdemod_out_d[1]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2898[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_i2.GSR = "ENABLED";
    LUT4 i7789_3_lut (.A(n78), .B(n78_adj_237), .C(n19811), .Z(n18923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7789_3_lut.init = 16'hcaca;
    FD1S3AX q_data_a_i11 (.D(cic_cosine_out[11]), .CK(cic_sine_clk), .Q(q_data_a[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam q_data_a_i11.GSR = "ENABLED";
    FD1S3AX q_data_a_i10 (.D(cic_cosine_out[10]), .CK(cic_sine_clk), .Q(q_data_a[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam q_data_a_i10.GSR = "ENABLED";
    FD1S3AX q_data_a_i9 (.D(cic_cosine_out[9]), .CK(cic_sine_clk), .Q(q_data_a[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam q_data_a_i9.GSR = "ENABLED";
    FD1S3AX q_data_a_i8 (.D(cic_cosine_out[8]), .CK(cic_sine_clk), .Q(q_data_a[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam q_data_a_i8.GSR = "ENABLED";
    FD1S3AX q_data_a_i7 (.D(cic_cosine_out[7]), .CK(cic_sine_clk), .Q(q_data_a[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam q_data_a_i7.GSR = "ENABLED";
    FD1S3AX q_data_a_i6 (.D(cic_cosine_out[6]), .CK(cic_sine_clk), .Q(q_data_a[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam q_data_a_i6.GSR = "ENABLED";
    FD1S3AX q_data_a_i5 (.D(cic_cosine_out[5]), .CK(cic_sine_clk), .Q(q_data_a[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam q_data_a_i5.GSR = "ENABLED";
    FD1S3AX q_data_a_i4 (.D(cic_cosine_out[4]), .CK(cic_sine_clk), .Q(q_data_a[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam q_data_a_i4.GSR = "ENABLED";
    LUT4 i7787_3_lut (.A(n73), .B(n73_adj_238), .C(n19811), .Z(n18921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7787_3_lut.init = 16'hcaca;
    LUT4 i7786_3_lut (.A(n75), .B(n75_adj_239), .C(n19811), .Z(n18920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7786_3_lut.init = 16'hcaca;
    FD1S3AX i_data_b_i0 (.D(\cic_sine_out[0] ), .CK(cic_sine_clk), .Q(i_data_b[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam i_data_b_i0.GSR = "ENABLED";
    LUT4 i7784_3_lut (.A(n70), .B(n70_adj_240), .C(n19811), .Z(n18918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7784_3_lut.init = 16'hcaca;
    LUT4 i7783_3_lut (.A(n72), .B(n72_adj_241), .C(n19811), .Z(n18917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7783_3_lut.init = 16'hcaca;
    LUT4 i7781_3_lut (.A(n67), .B(n67_adj_242), .C(n19811), .Z(n18915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7781_3_lut.init = 16'hcaca;
    LUT4 i7780_3_lut (.A(n69), .B(n69_adj_243), .C(n19811), .Z(n18914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7780_3_lut.init = 16'hcaca;
    LUT4 i7778_3_lut (.A(n64), .B(n64_adj_244), .C(n19811), .Z(n18912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7778_3_lut.init = 16'hcaca;
    LUT4 i7777_3_lut (.A(n66), .B(n66_adj_245), .C(n19811), .Z(n18911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7777_3_lut.init = 16'hcaca;
    FD1S3AX q_data_a_i0 (.D(cic_cosine_out[0]), .CK(cic_sine_clk), .Q(q_data_a[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam q_data_a_i0.GSR = "ENABLED";
    FD1S3AX amdemod_out_i1 (.D(amdemod_out_d[0]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2898[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_i1.GSR = "ENABLED";
    FD1S3AX q_data_a_i3 (.D(cic_cosine_out[3]), .CK(cic_sine_clk), .Q(q_data_a[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam q_data_a_i3.GSR = "ENABLED";
    FD1S3AX q_data_a_i2 (.D(cic_cosine_out[2]), .CK(cic_sine_clk), .Q(q_data_a[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam q_data_a_i2.GSR = "ENABLED";
    LUT4 i7775_3_lut (.A(n61), .B(n61_adj_246), .C(n19811), .Z(n18909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7775_3_lut.init = 16'hcaca;
    LUT4 i7774_3_lut (.A(n63), .B(n63_adj_247), .C(n19811), .Z(n18908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7774_3_lut.init = 16'hcaca;
    FD1S3AX i_data_b_i10 (.D(led_0_4), .CK(cic_sine_clk), .Q(i_data_b[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam i_data_b_i10.GSR = "ENABLED";
    FD1S3AX i_data_b_i11 (.D(led_0_5), .CK(cic_sine_clk), .Q(i_data_b[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam i_data_b_i11.GSR = "ENABLED";
    LUT4 i7772_3_lut (.A(n58), .B(n58_adj_248), .C(n19811), .Z(n18906)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7772_3_lut.init = 16'hcaca;
    LUT4 i7765_3_lut (.A(n36), .B(n36_adj_249), .C(amdemod_out_d_11__N_2363), 
         .Z(n18899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7765_3_lut.init = 16'hcaca;
    LUT4 i7771_3_lut (.A(n60), .B(n60_adj_250), .C(n19811), .Z(n18905)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7771_3_lut.init = 16'hcaca;
    LUT4 i7766_3_lut (.A(n34), .B(n34_adj_251), .C(amdemod_out_d_11__N_2363), 
         .Z(n18900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7766_3_lut.init = 16'hcaca;
    LUT4 i7763_3_lut (.A(n55), .B(n55_adj_252), .C(n19811), .Z(n18897)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7763_3_lut.init = 16'hcaca;
    LUT4 i7762_3_lut (.A(n57), .B(n57_adj_253), .C(n19811), .Z(n18896)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7762_3_lut.init = 16'hcaca;
    LUT4 i7757_3_lut (.A(n52), .B(n52_adj_254), .C(n19811), .Z(n18891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7757_3_lut.init = 16'hcaca;
    LUT4 i7756_3_lut (.A(n54), .B(n54_adj_255), .C(n19811), .Z(n18890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7756_3_lut.init = 16'hcaca;
    LUT4 i7882_3_lut (.A(n36_adj_256), .B(n36_adj_257), .C(n19815), .Z(n19016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7882_3_lut.init = 16'hcaca;
    LUT4 i7745_3_lut (.A(n49), .B(n49_adj_258), .C(n19811), .Z(n18879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7745_3_lut.init = 16'hcaca;
    LUT4 i7883_3_lut (.A(n34_adj_259), .B(n34_adj_260), .C(n19815), .Z(n19017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7883_3_lut.init = 16'hcaca;
    LUT4 i7744_3_lut (.A(n51_adj_261), .B(n51_adj_262), .C(n19811), .Z(n18878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7744_3_lut.init = 16'hcaca;
    LUT4 i7742_3_lut (.A(n46_adj_263), .B(n46_adj_264), .C(n19811), .Z(n18876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7742_3_lut.init = 16'hcaca;
    LUT4 i7741_3_lut (.A(n48_adj_265), .B(n48_adj_266), .C(n19811), .Z(n18875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7741_3_lut.init = 16'hcaca;
    LUT4 i7739_3_lut (.A(n43_adj_267), .B(n43_adj_268), .C(n19811), .Z(n18873)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7739_3_lut.init = 16'hcaca;
    LUT4 i7738_3_lut (.A(n45_adj_269), .B(n45_adj_270), .C(n19811), .Z(n18872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7738_3_lut.init = 16'hcaca;
    LUT4 i7736_3_lut (.A(n40_adj_271), .B(n40_adj_272), .C(n19811), .Z(n18870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7736_3_lut.init = 16'hcaca;
    LUT4 i7735_3_lut (.A(n42_adj_273), .B(n42_adj_274), .C(n19811), .Z(n18869)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7735_3_lut.init = 16'hcaca;
    LUT4 i7760_3_lut (.A(n76_adj_275), .B(n76_adj_276), .C(amdemod_out_d_11__N_2363), 
         .Z(n18894)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7760_3_lut.init = 16'hcaca;
    LUT4 i7837_3_lut (.A(n36_adj_277), .B(n36_adj_278), .C(n19813), .Z(n18971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7837_3_lut.init = 16'hcaca;
    LUT4 i7759_3_lut (.A(n78_adj_279), .B(n78_adj_280), .C(amdemod_out_d_11__N_2363), 
         .Z(n18893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7759_3_lut.init = 16'hcaca;
    LUT4 i7838_3_lut (.A(n34_adj_281), .B(n34_adj_282), .C(n19813), .Z(n18972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7838_3_lut.init = 16'hcaca;
    LUT4 i7792_3_lut (.A(n36_adj_283), .B(n36_adj_284), .C(n19811), .Z(n18926)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7792_3_lut.init = 16'hcaca;
    LUT4 i7793_3_lut (.A(n34_adj_285), .B(n34_adj_286), .C(n19811), .Z(n18927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7793_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), .Z(n4)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut.init = 16'h6666;
    LUT4 amdemod_out_d_11__I_17_rep_208_3_lut (.A(\amdemod_out_d_11__N_2379[14] ), 
         .B(\amdemod_out_d_11__N_2380[14] ), .C(n19815), .Z(n19312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_17_rep_208_3_lut.init = 16'hcaca;
    LUT4 n34_bdd_3_lut_8671 (.A(n34_adj_287), .B(n34_adj_288), .C(n19809), 
         .Z(n19724)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam n34_bdd_3_lut_8671.init = 16'h3535;
    LUT4 amdemod_out_d_11__I_13_rep_277 (.A(\amdemod_out_d_11__N_2369[11] ), 
         .B(\amdemod_out_d_11__N_2370[11] ), .C(amdemod_out_d_11__N_2363), 
         .Z(n19816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_13_rep_277.init = 16'hcaca;
    LUT4 n34_bdd_3_lut (.A(n36_adj_289), .B(n36_adj_290), .C(n19809), 
         .Z(n19725)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam n34_bdd_3_lut.init = 16'h3535;
    LUT4 amdemod_out_d_11__I_12_1_lut_3_lut (.A(\amdemod_out_d_11__N_2369[11] ), 
         .B(\amdemod_out_d_11__N_2370[11] ), .C(amdemod_out_d_11__N_2363), 
         .Z(amdemod_out_d_11__N_2367)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_12_1_lut_3_lut.init = 16'h3535;
    LUT4 i4322_3_lut (.A(n13878), .B(n42_adj_291), .C(\square_sum[25] ), 
         .Z(amdemod_out_d_11__N_2516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4322_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_17_rep_209_3_lut (.A(\amdemod_out_d_11__N_2379[14] ), 
         .B(\amdemod_out_d_11__N_2380[14] ), .C(n19815), .Z(n19313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_17_rep_209_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_17_rep_210_3_lut (.A(\amdemod_out_d_11__N_2379[14] ), 
         .B(\amdemod_out_d_11__N_2380[14] ), .C(n19815), .Z(n19314)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_17_rep_210_3_lut.init = 16'hcaca;
    LUT4 i7889_3_lut (.A(n64_adj_292), .B(n64_adj_293), .C(amdemod_out_d_11__N_2363), 
         .Z(n19023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7889_3_lut.init = 16'hcaca;
    LUT4 i7888_3_lut (.A(n66_adj_294), .B(n66_adj_295), .C(amdemod_out_d_11__N_2363), 
         .Z(n19022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7888_3_lut.init = 16'hcaca;
    LUT4 i7748_3_lut (.A(n67_adj_296), .B(n67_adj_297), .C(amdemod_out_d_11__N_2363), 
         .Z(n18882)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7748_3_lut.init = 16'hcaca;
    LUT4 i7747_3_lut (.A(n69_adj_298), .B(n69_adj_299), .C(amdemod_out_d_11__N_2363), 
         .Z(n18881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7747_3_lut.init = 16'hcaca;
    LUT4 i7907_3_lut (.A(n58_adj_300), .B(n58_adj_301), .C(amdemod_out_d_11__N_2363), 
         .Z(n19041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7907_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_13_rep_199_3_lut (.A(\amdemod_out_d_11__N_2369[11] ), 
         .B(\amdemod_out_d_11__N_2370[11] ), .C(amdemod_out_d_11__N_2363), 
         .Z(n19303)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_13_rep_199_3_lut.init = 16'hcaca;
    LUT4 i7906_3_lut (.A(n60_adj_302), .B(n60_adj_303), .C(amdemod_out_d_11__N_2363), 
         .Z(n19040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7906_3_lut.init = 16'hcaca;
    LUT4 i7832_3_lut (.A(n61_adj_304), .B(n61_adj_305), .C(amdemod_out_d_11__N_2363), 
         .Z(n18966)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7832_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_13_rep_200_3_lut (.A(\amdemod_out_d_11__N_2369[11] ), 
         .B(\amdemod_out_d_11__N_2370[11] ), .C(amdemod_out_d_11__N_2363), 
         .Z(n19304)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_13_rep_200_3_lut.init = 16'hcaca;
    PFUMX i7752 (.BLUT(n18884), .ALUT(n18885), .C0(n19303), .Z(amdemod_out_d_11__N_2594));
    LUT4 i7831_3_lut (.A(n63_adj_306), .B(n63_adj_307), .C(amdemod_out_d_11__N_2363), 
         .Z(n18965)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7831_3_lut.init = 16'hcaca;
    LUT4 i7904_3_lut (.A(n55_adj_308), .B(n55_adj_309), .C(amdemod_out_d_11__N_2363), 
         .Z(n19038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7904_3_lut.init = 16'hcaca;
    LUT4 i7903_3_lut (.A(n57_adj_310), .B(n57_adj_311), .C(amdemod_out_d_11__N_2363), 
         .Z(n19037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7903_3_lut.init = 16'hcaca;
    LUT4 i7901_3_lut (.A(n52_adj_312), .B(n52_adj_313), .C(amdemod_out_d_11__N_2363), 
         .Z(n19035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7901_3_lut.init = 16'hcaca;
    LUT4 i7900_3_lut (.A(n54_adj_314), .B(n54_adj_315), .C(amdemod_out_d_11__N_2363), 
         .Z(n19034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7900_3_lut.init = 16'hcaca;
    FD1S3AX amdemod_out_i10 (.D(amdemod_out_d[9]), .CK(cic_sine_clk), .Q(\amdemod_out[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_i10.GSR = "ENABLED";
    FD1S3AX amdemod_out_i9 (.D(amdemod_out_d[8]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2898[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_i9.GSR = "ENABLED";
    LUT4 i4324_3_lut_then_1_lut (.A(n39), .Z(n19836)) /* synthesis lut_function=(A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4324_3_lut_then_1_lut.init = 16'haaaa;
    LUT4 i4324_3_lut_else_1_lut (.A(\square_sum[22] ), .B(\amdemod_out_d_11__N_2365[3] ), 
         .C(n39_adj_316), .D(\square_sum[23] ), .Z(n19835)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4324_3_lut_else_1_lut.init = 16'hf0e4;
    LUT4 i7898_3_lut (.A(n49_adj_317), .B(n49_adj_318), .C(amdemod_out_d_11__N_2363), 
         .Z(n19032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7898_3_lut.init = 16'hcaca;
    LUT4 i7897_3_lut (.A(n51_adj_319), .B(n51_adj_320), .C(amdemod_out_d_11__N_2363), 
         .Z(n19031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7897_3_lut.init = 16'hcaca;
    LUT4 i7895_3_lut (.A(n46_adj_321), .B(n46_adj_322), .C(amdemod_out_d_11__N_2363), 
         .Z(n19029)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7895_3_lut.init = 16'hcaca;
    LUT4 i7894_3_lut (.A(n48_adj_323), .B(n48_adj_324), .C(amdemod_out_d_11__N_2363), 
         .Z(n19028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7894_3_lut.init = 16'hcaca;
    FD1S3AX amdemod_out_d__0_i1 (.D(amdemod_out_d_11__N_2412), .CK(cic_sine_clk), 
            .Q(amdemod_out_d[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_d__0_i1.GSR = "ENABLED";
    LUT4 i7794_3_lut_rep_270 (.A(n18926), .B(n18927), .C(n19810), .Z(n19809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7794_3_lut_rep_270.init = 16'hcaca;
    LUT4 i4333_3_lut_4_lut (.A(n19828), .B(n19827), .C(\amdemod_out_d_11__N_2365[14] ), 
         .D(n24), .Z(n13890)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4333_3_lut_4_lut.init = 16'hfe10;
    LUT4 i7892_3_lut (.A(n43_adj_325), .B(n43_adj_326), .C(amdemod_out_d_11__N_2363), 
         .Z(n19026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7892_3_lut.init = 16'hcaca;
    LUT4 i7891_3_lut (.A(n45_adj_327), .B(n45_adj_328), .C(amdemod_out_d_11__N_2363), 
         .Z(n19025)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7891_3_lut.init = 16'hcaca;
    LUT4 i7886_3_lut (.A(n40_adj_329), .B(n40_adj_330), .C(amdemod_out_d_11__N_2363), 
         .Z(n19020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7886_3_lut.init = 16'hcaca;
    LUT4 i4330_3_lut_then_1_lut (.A(n30), .Z(n19839)) /* synthesis lut_function=(A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4330_3_lut_then_1_lut.init = 16'haaaa;
    LUT4 i7880_3_lut (.A(n76_adj_331), .B(n76_adj_332), .C(n19815), .Z(n19014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7880_3_lut.init = 16'hcaca;
    LUT4 i7879_3_lut (.A(n78_adj_333), .B(n78_adj_334), .C(n19815), .Z(n19013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7879_3_lut.init = 16'hcaca;
    LUT4 i7885_3_lut (.A(n42_adj_335), .B(n42_adj_336), .C(amdemod_out_d_11__N_2363), 
         .Z(n19019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7885_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_29_rep_269 (.A(\amdemod_out_d_11__N_2409[14] ), 
         .B(\amdemod_out_d_11__N_2410[14] ), .C(n19809), .Z(n19808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_29_rep_269.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_26_1_lut_3_lut (.A(n18926), .B(n18927), .C(n19810), 
         .Z(amdemod_out_d_11__N_2402)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam amdemod_out_d_11__I_26_1_lut_3_lut.init = 16'h3535;
    LUT4 i4319_3_lut_4_lut (.A(n19828), .B(n19827), .C(\amdemod_out_d_11__N_2365[1] ), 
         .D(n45_adj_337), .Z(n13876)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4319_3_lut_4_lut.init = 16'hfe10;
    LUT4 i4330_3_lut_else_1_lut (.A(\square_sum[22] ), .B(\amdemod_out_d_11__N_2365[6] ), 
         .C(n30_adj_338), .D(\square_sum[23] ), .Z(n19838)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4330_3_lut_else_1_lut.init = 16'hf0e4;
    LUT4 i4321_3_lut_4_lut (.A(n19828), .B(n19827), .C(\amdemod_out_d_11__N_2365[2] ), 
         .D(n42_adj_339), .Z(n13878)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4321_3_lut_4_lut.init = 16'hfe10;
    PFUMX i7755 (.BLUT(n18887), .ALUT(n18888), .C0(n19303), .Z(amdemod_out_d_11__N_2597));
    LUT4 i7754_3_lut (.A(n73_adj_340), .B(n73_adj_341), .C(amdemod_out_d_11__N_2363), 
         .Z(n18888)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7754_3_lut.init = 16'hcaca;
    LUT4 i7753_3_lut (.A(n75_adj_342), .B(n75_adj_343), .C(amdemod_out_d_11__N_2363), 
         .Z(n18887)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7753_3_lut.init = 16'hcaca;
    LUT4 i7751_3_lut (.A(n70_adj_344), .B(n70_adj_345), .C(amdemod_out_d_11__N_2363), 
         .Z(n18885)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7751_3_lut.init = 16'hcaca;
    LUT4 i7877_3_lut (.A(n73_adj_346), .B(n73_adj_347), .C(n19815), .Z(n19011)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7877_3_lut.init = 16'hcaca;
    LUT4 i7876_3_lut (.A(n75_adj_348), .B(n75_adj_349), .C(n19815), .Z(n19010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7876_3_lut.init = 16'hcaca;
    LUT4 i7874_3_lut (.A(n70_adj_350), .B(n70_adj_351), .C(n19815), .Z(n19008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7874_3_lut.init = 16'hcaca;
    LUT4 i7873_3_lut (.A(n72_adj_352), .B(n72_adj_353), .C(n19815), .Z(n19007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7873_3_lut.init = 16'hcaca;
    LUT4 i7750_3_lut (.A(n72_adj_354), .B(n72_adj_355), .C(amdemod_out_d_11__N_2363), 
         .Z(n18884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7750_3_lut.init = 16'hcaca;
    LUT4 i7871_3_lut (.A(n67_adj_356), .B(n67_adj_357), .C(n19815), .Z(n19005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7871_3_lut.init = 16'hcaca;
    LUT4 i3390_1_lut (.A(\square_sum[25] ), .Z(\amdemod_out_d_11__N_2358[5] )) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam i3390_1_lut.init = 16'h5555;
    LUT4 i4328_3_lut_then_1_lut (.A(n33), .Z(n19842)) /* synthesis lut_function=(A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4328_3_lut_then_1_lut.init = 16'haaaa;
    LUT4 i7870_3_lut (.A(n69_adj_358), .B(n69_adj_359), .C(n19815), .Z(n19004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7870_3_lut.init = 16'hcaca;
    LUT4 i7868_3_lut (.A(n64_adj_360), .B(n64_adj_361), .C(n19815), .Z(n19002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7868_3_lut.init = 16'hcaca;
    LUT4 i4326_3_lut_else_1_lut (.A(\square_sum[22] ), .B(\amdemod_out_d_11__N_2365[4] ), 
         .C(n36_adj_362), .D(\square_sum[23] ), .Z(n19832)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4326_3_lut_else_1_lut.init = 16'hf0e4;
    LUT4 i4328_3_lut_else_1_lut (.A(\square_sum[22] ), .B(\amdemod_out_d_11__N_2365[5] ), 
         .C(n33_adj_363), .D(\square_sum[23] ), .Z(n19841)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4328_3_lut_else_1_lut.init = 16'hf0e4;
    LUT4 i7867_3_lut (.A(n66_adj_364), .B(n66_adj_365), .C(n19815), .Z(n19001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7867_3_lut.init = 16'hcaca;
    LUT4 i4326_3_lut_then_1_lut (.A(n36_adj_366), .Z(n19833)) /* synthesis lut_function=(A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4326_3_lut_then_1_lut.init = 16'haaaa;
    LUT4 i7865_3_lut (.A(n61_adj_367), .B(n61_adj_368), .C(n19815), .Z(n18999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7865_3_lut.init = 16'hcaca;
    LUT4 i7864_3_lut (.A(n63_adj_369), .B(n63_adj_370), .C(n19815), .Z(n18998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7864_3_lut.init = 16'hcaca;
    LUT4 i7862_3_lut (.A(n58_adj_371), .B(n58_adj_372), .C(n19815), .Z(n18996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7862_3_lut.init = 16'hcaca;
    LUT4 i7861_3_lut (.A(n60_adj_373), .B(n60_adj_374), .C(n19815), .Z(n18995)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7861_3_lut.init = 16'hcaca;
    LUT4 i7859_3_lut (.A(n55_adj_375), .B(n55_adj_376), .C(n19815), .Z(n18993)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7859_3_lut.init = 16'hcaca;
    LUT4 i7858_3_lut (.A(n57_adj_377), .B(n57_adj_378), .C(n19815), .Z(n18992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7858_3_lut.init = 16'hcaca;
    LUT4 i7856_3_lut (.A(n52_adj_379), .B(n52_adj_380), .C(n19815), .Z(n18990)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7856_3_lut.init = 16'hcaca;
    LUT4 i7855_3_lut (.A(n54_adj_381), .B(n54_adj_382), .C(n19815), .Z(n18989)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7855_3_lut.init = 16'hcaca;
    LUT4 i7853_3_lut (.A(n49_adj_383), .B(n49_adj_384), .C(n19815), .Z(n18987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7853_3_lut.init = 16'hcaca;
    LUT4 i7852_3_lut (.A(n51_adj_385), .B(n51_adj_386), .C(n19815), .Z(n18986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7852_3_lut.init = 16'hcaca;
    LUT4 i4332_3_lut_then_1_lut (.A(n30), .Z(n19845)) /* synthesis lut_function=(A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4332_3_lut_then_1_lut.init = 16'haaaa;
    LUT4 i4332_3_lut_else_1_lut (.A(\square_sum[22] ), .B(\amdemod_out_d_11__N_2365[7] ), 
         .C(n27), .D(\square_sum[23] ), .Z(n19844)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4332_3_lut_else_1_lut.init = 16'hf0e4;
    PFUMX i7887 (.BLUT(n19019), .ALUT(n19020), .C0(n19304), .Z(amdemod_out_d_11__N_2564));
    LUT4 i7850_3_lut (.A(n46_adj_387), .B(n46_adj_388), .C(n19815), .Z(n18984)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7850_3_lut.init = 16'hcaca;
    LUT4 i7849_3_lut (.A(n48_adj_389), .B(n48_adj_390), .C(n19815), .Z(n18983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7849_3_lut.init = 16'hcaca;
    PFUMX i7893 (.BLUT(n19025), .ALUT(n19026), .C0(n19304), .Z(amdemod_out_d_11__N_2567));
    LUT4 i4259_4_lut (.A(n46_adj_391), .B(n48_adj_392), .C(n13821), .D(n19828), 
         .Z(n13815)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4259_4_lut.init = 16'hccca;
    FD1S3AX amdemod_out_d__0_i2 (.D(amdemod_out_d_11__N_2407), .CK(cic_sine_clk), 
            .Q(amdemod_out_d[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_d__0_i2.GSR = "ENABLED";
    LUT4 i3357_2_lut (.A(\square_sum[25] ), .B(\square_sum[22] ), .Z(n13821)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(58[20:38])
    defparam i3357_2_lut.init = 16'heeee;
    FD1S3AX amdemod_out_d__0_i3 (.D(amdemod_out_d_11__N_2402), .CK(cic_sine_clk), 
            .Q(amdemod_out_d[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_d__0_i3.GSR = "ENABLED";
    FD1S3AX amdemod_out_d__0_i4 (.D(amdemod_out_d_11__N_2397), .CK(cic_sine_clk), 
            .Q(amdemod_out_d[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_d__0_i4.GSR = "ENABLED";
    FD1S3AX amdemod_out_d__0_i5 (.D(amdemod_out_d_11__N_2392), .CK(cic_sine_clk), 
            .Q(amdemod_out_d[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_d__0_i5.GSR = "ENABLED";
    FD1S3AX amdemod_out_d__0_i6 (.D(amdemod_out_d_11__N_2387), .CK(cic_sine_clk), 
            .Q(amdemod_out_d[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_d__0_i6.GSR = "ENABLED";
    FD1S3AX amdemod_out_d__0_i7 (.D(amdemod_out_d_11__N_2382), .CK(cic_sine_clk), 
            .Q(amdemod_out_d[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_d__0_i7.GSR = "ENABLED";
    FD1S3AX amdemod_out_d__0_i8 (.D(amdemod_out_d_11__N_2377), .CK(cic_sine_clk), 
            .Q(amdemod_out_d[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_d__0_i8.GSR = "ENABLED";
    FD1S3AX amdemod_out_d__0_i9 (.D(amdemod_out_d_11__N_2372), .CK(cic_sine_clk), 
            .Q(amdemod_out_d[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_d__0_i9.GSR = "ENABLED";
    FD1S3AX amdemod_out_d__0_i10 (.D(amdemod_out_d_11__N_2367), .CK(cic_sine_clk), 
            .Q(amdemod_out_d[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam amdemod_out_d__0_i10.GSR = "ENABLED";
    LUT4 amdemod_out_d_11__I_13_rep_201_3_lut (.A(\amdemod_out_d_11__N_2369[11] ), 
         .B(\amdemod_out_d_11__N_2370[11] ), .C(amdemod_out_d_11__N_2363), 
         .Z(n19305)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_13_rep_201_3_lut.init = 16'hcaca;
    LUT4 i7847_3_lut (.A(n43_adj_393), .B(n43_adj_394), .C(n19815), .Z(n18981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7847_3_lut.init = 16'hcaca;
    PFUMX i7896 (.BLUT(n19028), .ALUT(n19029), .C0(n19304), .Z(amdemod_out_d_11__N_2570));
    LUT4 amdemod_out_d_11__I_25_rep_271 (.A(\amdemod_out_d_11__N_2399[14] ), 
         .B(\amdemod_out_d_11__N_2400[14] ), .C(n19811), .Z(n19810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_25_rep_271.init = 16'hcaca;
    PFUMX i7899 (.BLUT(n19031), .ALUT(n19032), .C0(n19305), .Z(amdemod_out_d_11__N_2573));
    LUT4 amdemod_out_d_11__I_24_1_lut_3_lut (.A(\amdemod_out_d_11__N_2399[14] ), 
         .B(\amdemod_out_d_11__N_2400[14] ), .C(n19811), .Z(amdemod_out_d_11__N_2397)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_24_1_lut_3_lut.init = 16'h3535;
    LUT4 i7846_3_lut (.A(n45_adj_395), .B(n45_adj_396), .C(n19815), .Z(n18980)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7846_3_lut.init = 16'hcaca;
    LUT4 i7841_3_lut (.A(n40_adj_397), .B(n40_adj_398), .C(n19815), .Z(n18975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7841_3_lut.init = 16'hcaca;
    LUT4 i7840_3_lut (.A(n42_adj_399), .B(n42_adj_400), .C(n19815), .Z(n18974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7840_3_lut.init = 16'hcaca;
    PFUMX i7902 (.BLUT(n19034), .ALUT(n19035), .C0(n19305), .Z(amdemod_out_d_11__N_2576));
    LUT4 i7835_3_lut (.A(n76_adj_401), .B(n76_adj_402), .C(n19813), .Z(n18969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7835_3_lut.init = 16'hcaca;
    LUT4 i3239_2_lut_rep_288 (.A(\square_sum[25] ), .B(\square_sum[22] ), 
         .Z(n19827)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i3239_2_lut_rep_288.init = 16'h4444;
    LUT4 i7839_3_lut_rep_272 (.A(n18971), .B(n18972), .C(n19812), .Z(n19811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7839_3_lut_rep_272.init = 16'hcaca;
    PFUMX i7905 (.BLUT(n19037), .ALUT(n19038), .C0(n19305), .Z(amdemod_out_d_11__N_2579));
    LUT4 i4198_3_lut_rep_289 (.A(\square_sum[23] ), .B(\square_sum[25] ), 
         .C(\square_sum[22] ), .Z(n19828)) /* synthesis lut_function=(A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4198_3_lut_rep_289.init = 16'ha2a2;
    LUT4 amdemod_out_d_11__I_25_rep_202_3_lut (.A(\amdemod_out_d_11__N_2399[14] ), 
         .B(\amdemod_out_d_11__N_2400[14] ), .C(n19811), .Z(n19306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_25_rep_202_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_22_1_lut_3_lut (.A(n18971), .B(n18972), .C(n19812), 
         .Z(amdemod_out_d_11__N_2392)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam amdemod_out_d_11__I_22_1_lut_3_lut.init = 16'h3535;
    LUT4 i7834_3_lut (.A(n78_adj_403), .B(n78_adj_404), .C(n19813), .Z(n18968)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7834_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_25_rep_203_3_lut (.A(\amdemod_out_d_11__N_2399[14] ), 
         .B(\amdemod_out_d_11__N_2400[14] ), .C(n19811), .Z(n19307)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_25_rep_203_3_lut.init = 16'hcaca;
    LUT4 i7829_3_lut (.A(n73_adj_405), .B(n73_adj_406), .C(n19813), .Z(n18963)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7829_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_25_rep_204_3_lut (.A(\amdemod_out_d_11__N_2399[14] ), 
         .B(\amdemod_out_d_11__N_2400[14] ), .C(n19811), .Z(n19308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_25_rep_204_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_21_rep_205_3_lut (.A(\amdemod_out_d_11__N_2389[14] ), 
         .B(\amdemod_out_d_11__N_2390[14] ), .C(n19813), .Z(n19309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_21_rep_205_3_lut.init = 16'hcaca;
    LUT4 i7828_3_lut (.A(n75_adj_407), .B(n75_adj_408), .C(n19813), .Z(n18962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7828_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_21_rep_206_3_lut (.A(\amdemod_out_d_11__N_2389[14] ), 
         .B(\amdemod_out_d_11__N_2390[14] ), .C(n19813), .Z(n19310)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_21_rep_206_3_lut.init = 16'hcaca;
    LUT4 i7826_3_lut (.A(n70_adj_409), .B(n70_adj_410), .C(n19813), .Z(n18960)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7826_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_21_rep_207_3_lut (.A(\amdemod_out_d_11__N_2389[14] ), 
         .B(\amdemod_out_d_11__N_2390[14] ), .C(n19813), .Z(n19311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_21_rep_207_3_lut.init = 16'hcaca;
    PFUMX i7833 (.BLUT(n18965), .ALUT(n18966), .C0(n19303), .Z(amdemod_out_d_11__N_2585));
    LUT4 i7825_3_lut (.A(n72_adj_411), .B(n72_adj_412), .C(n19813), .Z(n18959)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7825_3_lut.init = 16'hcaca;
    LUT4 i7823_3_lut (.A(n67_adj_413), .B(n67_adj_414), .C(n19813), .Z(n18957)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7823_3_lut.init = 16'hcaca;
    PFUMX i7908 (.BLUT(n19040), .ALUT(n19041), .C0(n19305), .Z(amdemod_out_d_11__N_2582));
    LUT4 i7822_3_lut (.A(n69_adj_415), .B(n69_adj_416), .C(n19813), .Z(n18956)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7822_3_lut.init = 16'hcaca;
    LUT4 i3241_2_lut_rep_285_3_lut_3_lut (.A(\square_sum[23] ), .B(\square_sum[25] ), 
         .C(\square_sum[22] ), .Z(n19824)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i3241_2_lut_rep_285_3_lut_3_lut.init = 16'hb2b2;
    LUT4 i7820_3_lut (.A(n64_adj_417), .B(n64_adj_418), .C(n19813), .Z(n18954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7820_3_lut.init = 16'hcaca;
    LUT4 i7819_3_lut (.A(n66_adj_419), .B(n66_adj_420), .C(n19813), .Z(n18953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7819_3_lut.init = 16'hcaca;
    LUT4 i7817_3_lut (.A(n61_adj_421), .B(n61_adj_422), .C(n19813), .Z(n18951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7817_3_lut.init = 16'hcaca;
    LUT4 i7816_3_lut (.A(n63_adj_423), .B(n63_adj_424), .C(n19813), .Z(n18950)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7816_3_lut.init = 16'hcaca;
    LUT4 i7814_3_lut (.A(n58_adj_425), .B(n58_adj_426), .C(n19813), .Z(n18948)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7814_3_lut.init = 16'hcaca;
    LUT4 i7813_3_lut (.A(n60_adj_427), .B(n60_adj_428), .C(n19813), .Z(n18947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7813_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_21_rep_273 (.A(\amdemod_out_d_11__N_2389[14] ), 
         .B(\amdemod_out_d_11__N_2390[14] ), .C(n19813), .Z(n19812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_21_rep_273.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_20_1_lut_3_lut (.A(\amdemod_out_d_11__N_2389[14] ), 
         .B(\amdemod_out_d_11__N_2390[14] ), .C(n19813), .Z(amdemod_out_d_11__N_2387)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_20_1_lut_3_lut.init = 16'h3535;
    LUT4 i7884_3_lut_rep_274 (.A(n19016), .B(n19017), .C(n19814), .Z(n19813)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7884_3_lut_rep_274.init = 16'hcaca;
    LUT4 i7811_3_lut (.A(n55_adj_429), .B(n55_adj_430), .C(n19813), .Z(n18945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7811_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_18_1_lut_3_lut (.A(n19016), .B(n19017), .C(n19814), 
         .Z(amdemod_out_d_11__N_2382)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam amdemod_out_d_11__I_18_1_lut_3_lut.init = 16'h3535;
    LUT4 i7810_3_lut (.A(n57_adj_431), .B(n57_adj_432), .C(n19813), .Z(n18944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7810_3_lut.init = 16'hcaca;
    PFUMX i7749 (.BLUT(n18881), .ALUT(n18882), .C0(n19816), .Z(amdemod_out_d_11__N_2591));
    LUT4 i7808_3_lut (.A(n52_adj_433), .B(n52_adj_434), .C(n19813), .Z(n18942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7808_3_lut.init = 16'hcaca;
    PFUMX i7890 (.BLUT(n19022), .ALUT(n19023), .C0(n19304), .Z(amdemod_out_d_11__N_2588));
    LUT4 i7807_3_lut (.A(n54_adj_435), .B(n54_adj_436), .C(n19813), .Z(n18941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7807_3_lut.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_17_rep_275 (.A(\amdemod_out_d_11__N_2379[14] ), 
         .B(\amdemod_out_d_11__N_2380[14] ), .C(n19815), .Z(n19814)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_17_rep_275.init = 16'hcaca;
    LUT4 amdemod_out_d_11__I_28_1_lut_3_lut (.A(\amdemod_out_d_11__N_2409[14] ), 
         .B(\amdemod_out_d_11__N_2410[14] ), .C(n19809), .Z(amdemod_out_d_11__N_2407)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(57[18] 59[12])
    defparam amdemod_out_d_11__I_28_1_lut_3_lut.init = 16'h3535;
    LUT4 i7805_3_lut (.A(n49_adj_437), .B(n49_adj_438), .C(n19813), .Z(n18939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7805_3_lut.init = 16'hcaca;
    LUT4 i4334_3_lut (.A(n13890), .B(n30), .C(\square_sum[25] ), .Z(amdemod_out_d_11__N_2363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(56[20:38])
    defparam i4334_3_lut.init = 16'hcaca;
    PFUMX i8672 (.BLUT(n19725), .ALUT(n19724), .C0(n19808), .Z(amdemod_out_d_11__N_2412));
    PFUMX i7761 (.BLUT(n18893), .ALUT(n18894), .C0(n19303), .Z(amdemod_out_d_11__N_2600));
    PFUMX i7737 (.BLUT(n18869), .ALUT(n18870), .C0(n19810), .Z(amdemod_out_d_11__N_2798));
    PFUMX i7740 (.BLUT(n18872), .ALUT(n18873), .C0(n19306), .Z(amdemod_out_d_11__N_2801));
    PFUMX i7743 (.BLUT(n18875), .ALUT(n18876), .C0(n19306), .Z(amdemod_out_d_11__N_2804));
    PFUMX i7746 (.BLUT(n18878), .ALUT(n18879), .C0(n19306), .Z(amdemod_out_d_11__N_2807));
    PFUMX i7758 (.BLUT(n18890), .ALUT(n18891), .C0(n19306), .Z(amdemod_out_d_11__N_2810));
    PFUMX i7764 (.BLUT(n18896), .ALUT(n18897), .C0(n19307), .Z(amdemod_out_d_11__N_2813));
    PFUMX i7773 (.BLUT(n18905), .ALUT(n18906), .C0(n19307), .Z(amdemod_out_d_11__N_2816));
    PFUMX i7776 (.BLUT(n18908), .ALUT(n18909), .C0(n19307), .Z(amdemod_out_d_11__N_2819));
    PFUMX i7779 (.BLUT(n18911), .ALUT(n18912), .C0(n19307), .Z(amdemod_out_d_11__N_2822));
    PFUMX i7782 (.BLUT(n18914), .ALUT(n18915), .C0(n19308), .Z(amdemod_out_d_11__N_2825));
    PFUMX i7785 (.BLUT(n18917), .ALUT(n18918), .C0(n19308), .Z(amdemod_out_d_11__N_2828));
    PFUMX i7788 (.BLUT(n18920), .ALUT(n18921), .C0(n19308), .Z(amdemod_out_d_11__N_2831));
    PFUMX i7791 (.BLUT(n18923), .ALUT(n18924), .C0(n19308), .Z(amdemod_out_d_11__N_2834));
    PFUMX i7797 (.BLUT(n18929), .ALUT(n18930), .C0(n19812), .Z(amdemod_out_d_11__N_2720));
    PFUMX i7800 (.BLUT(n18932), .ALUT(n18933), .C0(n19309), .Z(amdemod_out_d_11__N_2723));
    PFUMX i7803 (.BLUT(n18935), .ALUT(n18936), .C0(n19309), .Z(amdemod_out_d_11__N_2726));
    PFUMX i7806 (.BLUT(n18938), .ALUT(n18939), .C0(n19309), .Z(amdemod_out_d_11__N_2729));
    PFUMX i7809 (.BLUT(n18941), .ALUT(n18942), .C0(n19309), .Z(amdemod_out_d_11__N_2732));
    PFUMX i7812 (.BLUT(n18944), .ALUT(n18945), .C0(n19310), .Z(amdemod_out_d_11__N_2735));
    PFUMX i7815 (.BLUT(n18947), .ALUT(n18948), .C0(n19310), .Z(amdemod_out_d_11__N_2738));
    PFUMX i7818 (.BLUT(n18950), .ALUT(n18951), .C0(n19310), .Z(amdemod_out_d_11__N_2741));
    PFUMX i7821 (.BLUT(n18953), .ALUT(n18954), .C0(n19310), .Z(amdemod_out_d_11__N_2744));
    PFUMX i7824 (.BLUT(n18956), .ALUT(n18957), .C0(n19311), .Z(amdemod_out_d_11__N_2747));
    PFUMX i7827 (.BLUT(n18959), .ALUT(n18960), .C0(n19311), .Z(amdemod_out_d_11__N_2750));
    PFUMX i7830 (.BLUT(n18962), .ALUT(n18963), .C0(n19311), .Z(amdemod_out_d_11__N_2753));
    PFUMX i7836 (.BLUT(n18968), .ALUT(n18969), .C0(n19311), .Z(amdemod_out_d_11__N_2756));
    FD1S3AX i_data_b_i9 (.D(led_0_3), .CK(cic_sine_clk), .Q(i_data_b[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=6, LSE_RCOL=5, LSE_LLINE=219, LSE_RLINE=224 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(91[9] 100[6])
    defparam i_data_b_i9.GSR = "ENABLED";
    PFUMX i7842 (.BLUT(n18974), .ALUT(n18975), .C0(n19814), .Z(amdemod_out_d_11__N_2642));
    PFUMX i7848 (.BLUT(n18980), .ALUT(n18981), .C0(n19312), .Z(amdemod_out_d_11__N_2645));
    PFUMX i7851 (.BLUT(n18983), .ALUT(n18984), .C0(n19312), .Z(amdemod_out_d_11__N_2648));
    PFUMX i8755 (.BLUT(n19844), .ALUT(n19845), .C0(\square_sum[25] ), 
          .Z(amdemod_out_d_11__N_2501));
    PFUMX i7854 (.BLUT(n18986), .ALUT(n18987), .C0(n19312), .Z(amdemod_out_d_11__N_2651));
    PFUMX i7857 (.BLUT(n18989), .ALUT(n18990), .C0(n19312), .Z(amdemod_out_d_11__N_2654));
    PFUMX i7860 (.BLUT(n18992), .ALUT(n18993), .C0(n19313), .Z(amdemod_out_d_11__N_2657));
    PFUMX i8753 (.BLUT(n19841), .ALUT(n19842), .C0(\square_sum[25] ), 
          .Z(amdemod_out_d_11__N_2507));
    PFUMX i7863 (.BLUT(n18995), .ALUT(n18996), .C0(n19313), .Z(amdemod_out_d_11__N_2660));
    PFUMX i7866 (.BLUT(n18998), .ALUT(n18999), .C0(n19313), .Z(amdemod_out_d_11__N_2663));
    PFUMX i7869 (.BLUT(n19001), .ALUT(n19002), .C0(n19313), .Z(amdemod_out_d_11__N_2666));
    PFUMX i7872 (.BLUT(n19004), .ALUT(n19005), .C0(n19314), .Z(amdemod_out_d_11__N_2669));
    PFUMX i8751 (.BLUT(n19838), .ALUT(n19839), .C0(\square_sum[25] ), 
          .Z(amdemod_out_d_11__N_2504));
    PFUMX i7875 (.BLUT(n19007), .ALUT(n19008), .C0(n19314), .Z(amdemod_out_d_11__N_2672));
    PFUMX i7878 (.BLUT(n19010), .ALUT(n19011), .C0(n19314), .Z(amdemod_out_d_11__N_2675));
    PFUMX i7881 (.BLUT(n19013), .ALUT(n19014), .C0(n19314), .Z(amdemod_out_d_11__N_2678));
    PFUMX i8749 (.BLUT(n19835), .ALUT(n19836), .C0(\square_sum[25] ), 
          .Z(amdemod_out_d_11__N_2513));
    PFUMX i8747 (.BLUT(n19832), .ALUT(n19833), .C0(\square_sum[25] ), 
          .Z(amdemod_out_d_11__N_2510));
    Multiplier Multiplier2 (.cic_sine_clk(cic_sine_clk), .VCC_net(VCC_net), 
            .GND_net(GND_net), .q_data_a({q_data_a}), .q_squared({q_squared})) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(79[14] 85[27])
    Multiplier_U1 Multiplier1 (.cic_sine_clk(cic_sine_clk), .VCC_net(VCC_net), 
            .GND_net(GND_net), .i_data_b({i_data_b}), .i_squared({i_squared})) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/AMDemod.v(71[14] 77[27])
    
endmodule
//
// Verilog Description of module Multiplier
//

module Multiplier (cic_sine_clk, VCC_net, GND_net, q_data_a, q_squared) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input cic_sine_clk;
    input VCC_net;
    input GND_net;
    input [11:0]q_data_a;
    output [23:0]q_squared;
    
    wire cic_sine_clk /* synthesis SET_AS_NETWORK=cic_sine_clk, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(78[33:45])
    
    MULT18X18D dsp_mult_0 (.A17(q_data_a[11]), .A16(q_data_a[10]), .A15(q_data_a[9]), 
            .A14(q_data_a[8]), .A13(q_data_a[7]), .A12(q_data_a[6]), .A11(q_data_a[5]), 
            .A10(q_data_a[4]), .A9(q_data_a[3]), .A8(q_data_a[2]), .A7(q_data_a[1]), 
            .A6(q_data_a[0]), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(q_data_a[11]), 
            .B16(q_data_a[10]), .B15(q_data_a[9]), .B14(q_data_a[8]), 
            .B13(q_data_a[7]), .B12(q_data_a[6]), .B11(q_data_a[5]), .B10(q_data_a[4]), 
            .B9(q_data_a[3]), .B8(q_data_a[2]), .B7(q_data_a[1]), .B6(q_data_a[0]), 
            .B5(GND_net), .B4(GND_net), .B3(GND_net), .B2(GND_net), 
            .B1(GND_net), .B0(GND_net), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(cic_sine_clk), 
            .CE3(VCC_net), .CE2(VCC_net), .CE1(VCC_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .P35(q_squared[23]), .P34(q_squared[22]), .P33(q_squared[21]), 
            .P32(q_squared[20]), .P31(q_squared[19]), .P30(q_squared[18]), 
            .P29(q_squared[17]), .P28(q_squared[16]), .P27(q_squared[15]), 
            .P26(q_squared[14]), .P25(q_squared[13]), .P24(q_squared[12]), 
            .P23(q_squared[11]), .P22(q_squared[10]), .P21(q_squared[9]), 
            .P20(q_squared[8]), .P19(q_squared[7]), .P18(q_squared[6]), 
            .P17(q_squared[5]), .P16(q_squared[4]), .P15(q_squared[3]), 
            .P14(q_squared[2]), .P13(q_squared[1]), .P12(q_squared[0])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=79, LSE_RLINE=85 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Multiplier.v(84[16] 140[57])
    defparam dsp_mult_0.REG_INPUTA_CLK = "CLK0";
    defparam dsp_mult_0.REG_INPUTA_CE = "CE0";
    defparam dsp_mult_0.REG_INPUTA_RST = "RST0";
    defparam dsp_mult_0.REG_INPUTB_CLK = "CLK0";
    defparam dsp_mult_0.REG_INPUTB_CE = "CE0";
    defparam dsp_mult_0.REG_INPUTB_RST = "RST0";
    defparam dsp_mult_0.REG_INPUTC_CLK = "NONE";
    defparam dsp_mult_0.REG_INPUTC_CE = "CE0";
    defparam dsp_mult_0.REG_INPUTC_RST = "RST0";
    defparam dsp_mult_0.REG_PIPELINE_CLK = "CLK0";
    defparam dsp_mult_0.REG_PIPELINE_CE = "CE0";
    defparam dsp_mult_0.REG_PIPELINE_RST = "RST0";
    defparam dsp_mult_0.REG_OUTPUT_CLK = "CLK0";
    defparam dsp_mult_0.REG_OUTPUT_CE = "CE0";
    defparam dsp_mult_0.REG_OUTPUT_RST = "RST0";
    defparam dsp_mult_0.CLK0_DIV = "ENABLED";
    defparam dsp_mult_0.CLK1_DIV = "ENABLED";
    defparam dsp_mult_0.CLK2_DIV = "ENABLED";
    defparam dsp_mult_0.CLK3_DIV = "ENABLED";
    defparam dsp_mult_0.HIGHSPEED_CLK = "NONE";
    defparam dsp_mult_0.GSR = "ENABLED";
    defparam dsp_mult_0.CAS_MATCH_REG = "FALSE";
    defparam dsp_mult_0.SOURCEB_MODE = "B_SHIFT";
    defparam dsp_mult_0.MULT_BYPASS = "DISABLED";
    defparam dsp_mult_0.RESETMODE = "ASYNC";
    
endmodule
//
// Verilog Description of module Multiplier_U1
//

module Multiplier_U1 (cic_sine_clk, VCC_net, GND_net, i_data_b, i_squared) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input cic_sine_clk;
    input VCC_net;
    input GND_net;
    input [11:0]i_data_b;
    output [23:0]i_squared;
    
    wire cic_sine_clk /* synthesis SET_AS_NETWORK=cic_sine_clk, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(78[33:45])
    
    MULT18X18D dsp_mult_0 (.A17(i_data_b[11]), .A16(i_data_b[10]), .A15(i_data_b[9]), 
            .A14(i_data_b[8]), .A13(i_data_b[7]), .A12(i_data_b[6]), .A11(i_data_b[5]), 
            .A10(i_data_b[4]), .A9(i_data_b[3]), .A8(i_data_b[2]), .A7(i_data_b[1]), 
            .A6(i_data_b[0]), .A5(GND_net), .A4(GND_net), .A3(GND_net), 
            .A2(GND_net), .A1(GND_net), .A0(GND_net), .B17(i_data_b[11]), 
            .B16(i_data_b[10]), .B15(i_data_b[9]), .B14(i_data_b[8]), 
            .B13(i_data_b[7]), .B12(i_data_b[6]), .B11(i_data_b[5]), .B10(i_data_b[4]), 
            .B9(i_data_b[3]), .B8(i_data_b[2]), .B7(i_data_b[1]), .B6(i_data_b[0]), 
            .B5(GND_net), .B4(GND_net), .B3(GND_net), .B2(GND_net), 
            .B1(GND_net), .B0(GND_net), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(cic_sine_clk), 
            .CE3(VCC_net), .CE2(VCC_net), .CE1(VCC_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .P35(i_squared[23]), .P34(i_squared[22]), .P33(i_squared[21]), 
            .P32(i_squared[20]), .P31(i_squared[19]), .P30(i_squared[18]), 
            .P29(i_squared[17]), .P28(i_squared[16]), .P27(i_squared[15]), 
            .P26(i_squared[14]), .P25(i_squared[13]), .P24(i_squared[12]), 
            .P23(i_squared[11]), .P22(i_squared[10]), .P21(i_squared[9]), 
            .P20(i_squared[8]), .P19(i_squared[7]), .P18(i_squared[6]), 
            .P17(i_squared[5]), .P16(i_squared[4]), .P15(i_squared[3]), 
            .P14(i_squared[2]), .P13(i_squared[1]), .P12(i_squared[0])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=11, LSE_LCOL=14, LSE_RCOL=27, LSE_LLINE=71, LSE_RLINE=77 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/Multiplier.v(84[16] 140[57])
    defparam dsp_mult_0.REG_INPUTA_CLK = "CLK0";
    defparam dsp_mult_0.REG_INPUTA_CE = "CE0";
    defparam dsp_mult_0.REG_INPUTA_RST = "RST0";
    defparam dsp_mult_0.REG_INPUTB_CLK = "CLK0";
    defparam dsp_mult_0.REG_INPUTB_CE = "CE0";
    defparam dsp_mult_0.REG_INPUTB_RST = "RST0";
    defparam dsp_mult_0.REG_INPUTC_CLK = "NONE";
    defparam dsp_mult_0.REG_INPUTC_CE = "CE0";
    defparam dsp_mult_0.REG_INPUTC_RST = "RST0";
    defparam dsp_mult_0.REG_PIPELINE_CLK = "CLK0";
    defparam dsp_mult_0.REG_PIPELINE_CE = "CE0";
    defparam dsp_mult_0.REG_PIPELINE_RST = "RST0";
    defparam dsp_mult_0.REG_OUTPUT_CLK = "CLK0";
    defparam dsp_mult_0.REG_OUTPUT_CE = "CE0";
    defparam dsp_mult_0.REG_OUTPUT_RST = "RST0";
    defparam dsp_mult_0.CLK0_DIV = "ENABLED";
    defparam dsp_mult_0.CLK1_DIV = "ENABLED";
    defparam dsp_mult_0.CLK2_DIV = "ENABLED";
    defparam dsp_mult_0.CLK3_DIV = "ENABLED";
    defparam dsp_mult_0.HIGHSPEED_CLK = "NONE";
    defparam dsp_mult_0.GSR = "ENABLED";
    defparam dsp_mult_0.CAS_MATCH_REG = "FALSE";
    defparam dsp_mult_0.SOURCEB_MODE = "B_SHIFT";
    defparam dsp_mult_0.MULT_BYPASS = "DISABLED";
    defparam dsp_mult_0.RESETMODE = "ASYNC";
    
endmodule
//
// Verilog Description of module \CIC(REGISTER_WIDTH=72,DECIMATION_RATIO=4096) 
//

module \CIC(REGISTER_WIDTH=72,DECIMATION_RATIO=4096)  (comb_d7, n14, comb_d6, 
            n20, integrator_d_tmp, clk_80mhz, integrator_tmp, \cic_gain[0] , 
            integrator2, integrator2_71__N_1032, \cic_gain[1] , integrator3, 
            integrator3_71__N_1104, integrator4, integrator4_71__N_1176, 
            integrator5, integrator5_71__N_1248, comb6, comb6_71__N_1993, 
            cic_sine_clk, n27, comb7, comb7_71__N_2065, comb8, comb8_71__N_2137, 
            comb_d8, comb9, comb9_71__N_2209, comb_d9, integrator1, 
            integrator1_71__N_960, count, n26, n35, n34, n17, n16, 
            n29, n28, n37, n9, \comb10[67] , \comb10[69] , n8, 
            n36, n23, \comb10[68] , \comb10[70] , n22, n31, n30, 
            n25, n24, n33, n32, n21, n20_adj_115, n19, n18, 
            n25_adj_116, n24_adj_117, n23_adj_118, n22_adj_119, n3, 
            n31_adj_120, n30_adj_121, n29_adj_122, n28_adj_123, n27_adj_124, 
            n26_adj_125, n35_adj_126, n34_adj_127, n2, n37_adj_128, 
            n36_adj_129, n5, n7, n4, n6, n5_adj_130, n4_adj_131, 
            n3_adj_132, n2_adj_133, n17_adj_134, n16_adj_135, n15, 
            n14_adj_136, n11, n10, n13, n12, n25_adj_137, n24_adj_138, 
            n62, \comb10[60] , n23_adj_139, n22_adj_140, n21_adj_141, 
            n20_adj_142, n33_adj_143, n32_adj_144, n31_adj_145, n30_adj_146, 
            n29_adj_147, n28_adj_148, n37_adj_149, n36_adj_150, n3_adj_151, 
            n2_adj_152, n5_adj_153, n4_adj_154, n68, \comb10[66] , 
            n67_adj_228, n76, n78, cout, n79, n81, n82, n84, 
            n85, n87, n88, n90, n91, n93, led_0_2, n94, n96, 
            n97, n99, n100, n102, n103, n105, n67, \comb10[65] , 
            n106, n108, n109, n111, n66, \comb10[64] , n112, n114, 
            n115, n117, n118, n120, n64, \comb10[62] , n19_adj_159, 
            n63, \comb10[61] , n65, \comb10[63] , n7_adj_160, n6_adj_161, 
            n13_adj_162, n12_adj_163, n21_adj_164, n20_adj_165, n15_adj_166, 
            n14_adj_167, n23_adj_168, n22_adj_169, n9_adj_170, n8_adj_171, 
            n17_adj_172, n16_adj_173, n25_adj_174, n24_adj_175, n11_adj_176, 
            n10_adj_177, n19_adj_178, n18_adj_179, n27_adj_180, n26_adj_181, 
            n33_adj_182, n32_adj_183, n35_adj_184, n34_adj_185, n29_adj_186, 
            n28_adj_187, n37_adj_188, n36_adj_189, n3_adj_190, n2_adj_191, 
            n31_adj_192, n30_adj_193, n5_adj_194, n4_adj_195, n11_adj_196, 
            n10_adj_197, n17_adj_198, n16_adj_199, n13_adj_200, n12_adj_201, 
            n7_adj_202, n6_adj_203, n15_adj_204, n14_adj_205, n61_adj_206, 
            \comb10[59] , n19_adj_207, n18_adj_208, n9_adj_209, n8_adj_210, 
            n21_adj_211, led_0_1, led_0_0, \cic_sine_out[5] , n7_adj_212, 
            n6_adj_213, n13_adj_214, n12_adj_215, n15_adj_216, \cic_sine_out[4] , 
            \cic_sine_out[3] , \cic_sine_out[2] , \comb10[71] , \cic_cosine_out[11] , 
            n70, \cic_cosine_out[9] , \cic_cosine_out[8] , \cic_cosine_out[7] , 
            \cic_cosine_out[6] , \cic_cosine_out[5] , \cic_cosine_out[4] , 
            \cic_cosine_out[3] , \cic_cosine_out[2] , led_0_5, led_0_3, 
            n18_adj_217, n11_adj_218, n10_adj_219, n33_adj_220, n32_adj_221, 
            n9_adj_222, n8_adj_223, \cic_cosine_out[10] , led_0_4, \cic_sine_out[1] , 
            \cic_sine_out[0] , n27_adj_224, n26_adj_225, n35_adj_226, 
            n34_adj_227) /* synthesis syn_module_defined=1 */ ;
    output [71:0]comb_d7;
    output n14;
    output [71:0]comb_d6;
    output n20;
    output [71:0]integrator_d_tmp;
    input clk_80mhz;
    output [71:0]integrator_tmp;
    input \cic_gain[0] ;
    output [71:0]integrator2;
    input [71:0]integrator2_71__N_1032;
    input \cic_gain[1] ;
    output [71:0]integrator3;
    input [71:0]integrator3_71__N_1104;
    output [71:0]integrator4;
    input [71:0]integrator4_71__N_1176;
    output [71:0]integrator5;
    input [71:0]integrator5_71__N_1248;
    output [71:0]comb6;
    input [71:0]comb6_71__N_1993;
    output cic_sine_clk;
    output n27;
    output [71:0]comb7;
    input [71:0]comb7_71__N_2065;
    output [71:0]comb8;
    input [71:0]comb8_71__N_2137;
    output [71:0]comb_d8;
    output [71:0]comb9;
    input [71:0]comb9_71__N_2209;
    output [71:0]comb_d9;
    output [71:0]integrator1;
    input [71:0]integrator1_71__N_960;
    output [11:0]count;
    output n26;
    output n35;
    output n34;
    output n17;
    output n16;
    output n29;
    output n28;
    output n37;
    output n9;
    input \comb10[67] ;
    input \comb10[69] ;
    output n8;
    output n36;
    output n23;
    input \comb10[68] ;
    input \comb10[70] ;
    output n22;
    output n31;
    output n30;
    output n25;
    output n24;
    output n33;
    output n32;
    output n21;
    output n20_adj_115;
    output n19;
    output n18;
    output n25_adj_116;
    output n24_adj_117;
    output n23_adj_118;
    output n22_adj_119;
    output n3;
    output n31_adj_120;
    output n30_adj_121;
    output n29_adj_122;
    output n28_adj_123;
    output n27_adj_124;
    output n26_adj_125;
    output n35_adj_126;
    output n34_adj_127;
    output n2;
    output n37_adj_128;
    output n36_adj_129;
    output n5;
    output n7;
    output n4;
    output n6;
    output n5_adj_130;
    output n4_adj_131;
    output n3_adj_132;
    output n2_adj_133;
    output n17_adj_134;
    output n16_adj_135;
    output n15;
    output n14_adj_136;
    output n11;
    output n10;
    output n13;
    output n12;
    output n25_adj_137;
    output n24_adj_138;
    input n62;
    input \comb10[60] ;
    output n23_adj_139;
    output n22_adj_140;
    output n21_adj_141;
    output n20_adj_142;
    output n33_adj_143;
    output n32_adj_144;
    output n31_adj_145;
    output n30_adj_146;
    output n29_adj_147;
    output n28_adj_148;
    output n37_adj_149;
    output n36_adj_150;
    output n3_adj_151;
    output n2_adj_152;
    output n5_adj_153;
    output n4_adj_154;
    input n68;
    input \comb10[66] ;
    input [11:0]n67_adj_228;
    input n76;
    input n78;
    input cout;
    input n79;
    input n81;
    input n82;
    input n84;
    input n85;
    input n87;
    input n88;
    input n90;
    input n91;
    input n93;
    output led_0_2;
    input n94;
    input n96;
    input n97;
    input n99;
    input n100;
    input n102;
    input n103;
    input n105;
    input n67;
    input \comb10[65] ;
    input n106;
    input n108;
    input n109;
    input n111;
    input n66;
    input \comb10[64] ;
    input n112;
    input n114;
    input n115;
    input n117;
    input n118;
    input n120;
    input n64;
    input \comb10[62] ;
    output n19_adj_159;
    input n63;
    input \comb10[61] ;
    input n65;
    input \comb10[63] ;
    output n7_adj_160;
    output n6_adj_161;
    output n13_adj_162;
    output n12_adj_163;
    output n21_adj_164;
    output n20_adj_165;
    output n15_adj_166;
    output n14_adj_167;
    output n23_adj_168;
    output n22_adj_169;
    output n9_adj_170;
    output n8_adj_171;
    output n17_adj_172;
    output n16_adj_173;
    output n25_adj_174;
    output n24_adj_175;
    output n11_adj_176;
    output n10_adj_177;
    output n19_adj_178;
    output n18_adj_179;
    output n27_adj_180;
    output n26_adj_181;
    output n33_adj_182;
    output n32_adj_183;
    output n35_adj_184;
    output n34_adj_185;
    output n29_adj_186;
    output n28_adj_187;
    output n37_adj_188;
    output n36_adj_189;
    output n3_adj_190;
    output n2_adj_191;
    output n31_adj_192;
    output n30_adj_193;
    output n5_adj_194;
    output n4_adj_195;
    output n11_adj_196;
    output n10_adj_197;
    output n17_adj_198;
    output n16_adj_199;
    output n13_adj_200;
    output n12_adj_201;
    output n7_adj_202;
    output n6_adj_203;
    output n15_adj_204;
    output n14_adj_205;
    input n61_adj_206;
    input \comb10[59] ;
    output n19_adj_207;
    output n18_adj_208;
    output n9_adj_209;
    output n8_adj_210;
    output n21_adj_211;
    output led_0_1;
    output led_0_0;
    output \cic_sine_out[5] ;
    output n7_adj_212;
    output n6_adj_213;
    output n13_adj_214;
    output n12_adj_215;
    output n15_adj_216;
    output \cic_sine_out[4] ;
    output \cic_sine_out[3] ;
    output \cic_sine_out[2] ;
    input \comb10[71] ;
    output \cic_cosine_out[11] ;
    input n70;
    output \cic_cosine_out[9] ;
    output \cic_cosine_out[8] ;
    output \cic_cosine_out[7] ;
    output \cic_cosine_out[6] ;
    output \cic_cosine_out[5] ;
    output \cic_cosine_out[4] ;
    output \cic_cosine_out[3] ;
    output \cic_cosine_out[2] ;
    output led_0_5;
    output led_0_3;
    output n18_adj_217;
    output n11_adj_218;
    output n10_adj_219;
    output n33_adj_220;
    output n32_adj_221;
    output n9_adj_222;
    output n8_adj_223;
    output \cic_cosine_out[10] ;
    output led_0_4;
    output \cic_sine_out[1] ;
    output \cic_sine_out[0] ;
    output n27_adj_224;
    output n26_adj_225;
    output n35_adj_226;
    output n34_adj_227;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(61[34:43])
    wire cic_sine_clk /* synthesis SET_AS_NETWORK=cic_sine_clk, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(78[33:45])
    
    wire clk_80mhz_enable_291;
    wire [71:0]comb10;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[99:105])
    
    wire n63_c, n19869, n62_c, decimation_clk, clk_80mhz_enable_1456, 
        n14240, valid_comb, n19868;
    wire [11:0]count_11__N_1980;
    
    wire n61, n19872, n19871, n18858, n18842, n20283, n132, n67_c, 
        clk_80mhz_enable_873, n138, n73, n14270, decimation_clk_N_2353, 
        n18854, n18840;
    wire [71:0]comb10_71__N_2281;
    
    wire n131, n18796, n18780, n18788, clk_80mhz_enable_923, clk_80mhz_enable_973, 
        clk_80mhz_enable_1023, clk_80mhz_enable_1073, clk_80mhz_enable_1123, 
        n18792, clk_80mhz_enable_1173, n137, clk_80mhz_enable_1223, 
        clk_80mhz_enable_1273, clk_80mhz_enable_1323, clk_80mhz_enable_1373, 
        clk_80mhz_enable_1423, n137_adj_3194, n136, n68_adj_3196, n65_c, 
        n134, n133, n135, n70_c, n131_adj_3252, n136_adj_3258, n135_adj_3259, 
        n66_adj_3260, n134_adj_3261, n140, n133_adj_3267, n138_adj_3268, 
        n64_adj_3269, n132_adj_3270, n140_adj_3272, n19851, n19850, 
        n19860, n19859;
    
    LUT4 sub_28_inv_0_i60_1_lut (.A(comb_d7[59]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i54_1_lut (.A(comb_d6[53]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i54_1_lut.init = 16'h5555;
    FD1P3AX integrator_d_tmp_i0_i0 (.D(integrator_tmp[0]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i0.GSR = "ENABLED";
    LUT4 comb10_71__I_0_77_i63_3_lut (.A(comb10[62]), .B(comb10[63]), .C(\cic_gain[0] ), 
         .Z(n63_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i63_3_lut.init = 16'hcaca;
    FD1S3AX integrator2_i0 (.D(integrator2_71__N_1032[0]), .CK(clk_80mhz), 
            .Q(integrator2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i0.GSR = "ENABLED";
    LUT4 i11_3_lut_4_lut_then_3_lut (.A(\cic_gain[1] ), .B(comb10[67]), 
         .C(comb10[69]), .Z(n19869)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam i11_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 comb10_71__I_0_77_i62_3_lut (.A(comb10[61]), .B(comb10[62]), .C(\cic_gain[0] ), 
         .Z(n62_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i62_3_lut.init = 16'hcaca;
    FD1S3AX integrator3_i0 (.D(integrator3_71__N_1104[0]), .CK(clk_80mhz), 
            .Q(integrator3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i0.GSR = "ENABLED";
    FD1S3AX integrator4_i0 (.D(integrator4_71__N_1176[0]), .CK(clk_80mhz), 
            .Q(integrator4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i0.GSR = "ENABLED";
    FD1S3AX integrator5_i0 (.D(integrator5_71__N_1248[0]), .CK(clk_80mhz), 
            .Q(integrator5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i0.GSR = "ENABLED";
    FD1P3AX comb6_i0_i0 (.D(comb6_71__N_1993[0]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(comb6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i0 (.D(comb6[0]), .SP(clk_80mhz_enable_291), .CK(clk_80mhz), 
            .Q(comb_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i0.GSR = "ENABLED";
    FD1S3JX decimation_clk_62 (.D(n14240), .CK(clk_80mhz), .PD(clk_80mhz_enable_1456), 
            .Q(decimation_clk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam decimation_clk_62.GSR = "ENABLED";
    FD1S3AX valid_comb_63 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), .Q(valid_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63.GSR = "ENABLED";
    FD1S3AX data_clk_64 (.D(decimation_clk), .CK(clk_80mhz), .Q(cic_sine_clk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam data_clk_64.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i47_1_lut (.A(comb_d6[46]), .Z(n27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i47_1_lut.init = 16'h5555;
    FD1P3AX comb7_i0_i0 (.D(comb7_71__N_2065[0]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(comb7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i0 (.D(comb7[0]), .SP(clk_80mhz_enable_291), .CK(clk_80mhz), 
            .Q(comb_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX comb8_i0_i0 (.D(comb8_71__N_2137[0]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(comb8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i0 (.D(comb8[0]), .SP(clk_80mhz_enable_291), .CK(clk_80mhz), 
            .Q(comb_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX comb9_i0_i0 (.D(comb9_71__N_2209[0]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(comb9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i0 (.D(comb9[0]), .SP(clk_80mhz_enable_291), .CK(clk_80mhz), 
            .Q(comb_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i0.GSR = "ENABLED";
    FD1S3AX integrator1_i0 (.D(integrator1_71__N_960[0]), .CK(clk_80mhz), 
            .Q(integrator1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i0.GSR = "ENABLED";
    LUT4 i11_3_lut_4_lut_else_3_lut (.A(\cic_gain[1] ), .B(comb10[68]), 
         .C(comb10[70]), .Z(n19868)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam i11_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    FD1S3IX count__i0 (.D(count_11__N_1980[0]), .CK(clk_80mhz), .CD(clk_80mhz_enable_1456), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i0.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i48_1_lut (.A(comb_d6[47]), .Z(n26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i39_1_lut (.A(comb_d6[38]), .Z(n35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i40_1_lut (.A(comb_d6[39]), .Z(n34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i57_1_lut (.A(comb_d7[56]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i58_1_lut (.A(comb_d7[57]), .Z(n16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i45_1_lut (.A(comb_d6[44]), .Z(n29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 comb10_71__I_0_77_i61_3_lut (.A(comb10[60]), .B(comb10[61]), .C(\cic_gain[0] ), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i61_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i46_1_lut (.A(comb_d6[45]), .Z(n28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i37_1_lut (.A(comb_d6[36]), .Z(n37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i65_1_lut (.A(comb_d7[64]), .Z(n9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 i11_3_lut_4_lut_then_3_lut_adj_194 (.A(\cic_gain[1] ), .B(\comb10[67] ), 
         .C(\comb10[69] ), .Z(n19872)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam i11_3_lut_4_lut_then_3_lut_adj_194.init = 16'hd8d8;
    LUT4 sub_28_inv_0_i66_1_lut (.A(comb_d7[65]), .Z(n8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i38_1_lut (.A(comb_d6[37]), .Z(n36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i51_1_lut (.A(comb_d6[50]), .Z(n23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 i11_3_lut_4_lut_else_3_lut_adj_195 (.A(\cic_gain[1] ), .B(\comb10[68] ), 
         .C(\comb10[70] ), .Z(n19871)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam i11_3_lut_4_lut_else_3_lut_adj_195.init = 16'hd8d8;
    LUT4 sub_27_inv_0_i52_1_lut (.A(comb_d6[51]), .Z(n22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i43_1_lut (.A(comb_d6[42]), .Z(n31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i44_1_lut (.A(comb_d6[43]), .Z(n30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i49_1_lut (.A(comb_d6[48]), .Z(n25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_rep_325 (.A(n18858), .B(count[0]), .C(n18842), .D(count[11]), 
         .Z(n20283)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam i1_4_lut_rep_325.init = 16'h8000;
    LUT4 i1_4_lut_rep_326 (.A(n18858), .B(count[0]), .C(n18842), .D(count[11]), 
         .Z(clk_80mhz_enable_1456)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam i1_4_lut_rep_326.init = 16'h8000;
    LUT4 sub_27_inv_0_i50_1_lut (.A(comb_d6[49]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i41_1_lut (.A(comb_d6[40]), .Z(n33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i42_1_lut (.A(comb_d6[41]), .Z(n32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i53_1_lut (.A(comb_d7[52]), .Z(n21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i54_1_lut (.A(comb_d7[53]), .Z(n20_adj_115)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i55_1_lut (.A(comb_d7[54]), .Z(n19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i56_1_lut (.A(comb_d7[55]), .Z(n18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i49_1_lut (.A(comb_d7[48]), .Z(n25_adj_116)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i50_1_lut (.A(comb_d7[49]), .Z(n24_adj_117)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i51_1_lut (.A(comb_d7[50]), .Z(n23_adj_118)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i52_1_lut (.A(comb_d7[51]), .Z(n22_adj_119)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i71_1_lut (.A(comb_d7[70]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i43_1_lut (.A(comb_d7[42]), .Z(n31_adj_120)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i44_1_lut (.A(comb_d7[43]), .Z(n30_adj_121)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i45_1_lut (.A(comb_d7[44]), .Z(n29_adj_122)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i46_1_lut (.A(comb_d7[45]), .Z(n28_adj_123)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i47_1_lut (.A(comb_d7[46]), .Z(n27_adj_124)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i48_1_lut (.A(comb_d7[47]), .Z(n26_adj_125)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i39_1_lut (.A(comb_d7[38]), .Z(n35_adj_126)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i40_1_lut (.A(comb_d7[39]), .Z(n34_adj_127)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i72_1_lut (.A(comb_d7[71]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i37_1_lut (.A(comb_d7[36]), .Z(n37_adj_128)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i38_1_lut (.A(comb_d7[37]), .Z(n36_adj_129)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i69_1_lut (.A(comb_d7[68]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i67_1_lut (.A(comb_d8[66]), .Z(n7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i70_1_lut (.A(comb_d7[69]), .Z(n4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i68_1_lut (.A(comb_d8[67]), .Z(n6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i69_1_lut (.A(comb_d8[68]), .Z(n5_adj_130)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i70_1_lut (.A(comb_d8[69]), .Z(n4_adj_131)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i71_1_lut (.A(comb_d8[70]), .Z(n3_adj_132)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i72_1_lut (.A(comb_d8[71]), .Z(n2_adj_133)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i57_1_lut (.A(comb_d8[56]), .Z(n17_adj_134)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i58_1_lut (.A(comb_d8[57]), .Z(n16_adj_135)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i59_1_lut (.A(comb_d8[58]), .Z(n15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i60_1_lut (.A(comb_d8[59]), .Z(n14_adj_136)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i63_1_lut (.A(comb_d8[62]), .Z(n11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i64_1_lut (.A(comb_d8[63]), .Z(n10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i61_1_lut (.A(comb_d8[60]), .Z(n13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i62_1_lut (.A(comb_d8[61]), .Z(n12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i49_1_lut (.A(comb_d8[48]), .Z(n25_adj_137)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i50_1_lut (.A(comb_d8[49]), .Z(n24_adj_138)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 comb10_71__I_0_77_i132_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n62), .D(\comb10[60] ), .Z(n132)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i132_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_29_inv_0_i51_1_lut (.A(comb_d8[50]), .Z(n23_adj_139)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i52_1_lut (.A(comb_d8[51]), .Z(n22_adj_140)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i53_1_lut (.A(comb_d8[52]), .Z(n21_adj_141)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i54_1_lut (.A(comb_d8[53]), .Z(n20_adj_142)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i41_1_lut (.A(comb_d8[40]), .Z(n33_adj_143)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i42_1_lut (.A(comb_d8[41]), .Z(n32_adj_144)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i43_1_lut (.A(comb_d8[42]), .Z(n31_adj_145)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i44_1_lut (.A(comb_d8[43]), .Z(n30_adj_146)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 comb10_71__I_0_77_i67_3_lut (.A(comb10[66]), .B(comb10[67]), .C(\cic_gain[0] ), 
         .Z(n67_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i67_3_lut.init = 16'hcaca;
    LUT4 sub_29_inv_0_i45_1_lut (.A(comb_d8[44]), .Z(n29_adj_147)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i46_1_lut (.A(comb_d8[45]), .Z(n28_adj_148)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i37_1_lut (.A(comb_d8[36]), .Z(n37_adj_149)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i38_1_lut (.A(comb_d8[37]), .Z(n36_adj_150)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i71_1_lut (.A(integrator_d_tmp[70]), .Z(n3_adj_151)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i72_1_lut (.A(integrator_d_tmp[71]), .Z(n2_adj_152)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i69_1_lut (.A(integrator_d_tmp[68]), .Z(n5_adj_153)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i70_1_lut (.A(integrator_d_tmp[69]), .Z(n4_adj_154)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i70_1_lut.init = 16'h5555;
    FD1P3AX integrator_d_tmp_i0_i71 (.D(integrator_tmp[71]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i70 (.D(integrator_tmp[70]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i69 (.D(integrator_tmp[69]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i68 (.D(integrator_tmp[68]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i67 (.D(integrator_tmp[67]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i66 (.D(integrator_tmp[66]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i65 (.D(integrator_tmp[65]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i64 (.D(integrator_tmp[64]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i63 (.D(integrator_tmp[63]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i62 (.D(integrator_tmp[62]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i61 (.D(integrator_tmp[61]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i60 (.D(integrator_tmp[60]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i59 (.D(integrator_tmp[59]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i58 (.D(integrator_tmp[58]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i57 (.D(integrator_tmp[57]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i56 (.D(integrator_tmp[56]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i55 (.D(integrator_tmp[55]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i54 (.D(integrator_tmp[54]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i53 (.D(integrator_tmp[53]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i52 (.D(integrator_tmp[52]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i51 (.D(integrator_tmp[51]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i50 (.D(integrator_tmp[50]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i49 (.D(integrator_tmp[49]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i48 (.D(integrator_tmp[48]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i47 (.D(integrator_tmp[47]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i46 (.D(integrator_tmp[46]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i45 (.D(integrator_tmp[45]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i44 (.D(integrator_tmp[44]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i43 (.D(integrator_tmp[43]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i42 (.D(integrator_tmp[42]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i41 (.D(integrator_tmp[41]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i40 (.D(integrator_tmp[40]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i39 (.D(integrator_tmp[39]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i38 (.D(integrator_tmp[38]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i37 (.D(integrator_tmp[37]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i36 (.D(integrator_tmp[36]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i35 (.D(integrator_tmp[35]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i34 (.D(integrator_tmp[34]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i33 (.D(integrator_tmp[33]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i32 (.D(integrator_tmp[32]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i31 (.D(integrator_tmp[31]), .SP(clk_80mhz_enable_291), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i30 (.D(integrator_tmp[30]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i29 (.D(integrator_tmp[29]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i28 (.D(integrator_tmp[28]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i27 (.D(integrator_tmp[27]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i26 (.D(integrator_tmp[26]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i25 (.D(integrator_tmp[25]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i24 (.D(integrator_tmp[24]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i23 (.D(integrator_tmp[23]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i22 (.D(integrator_tmp[22]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i21 (.D(integrator_tmp[21]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i20 (.D(integrator_tmp[20]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i19 (.D(integrator_tmp[19]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i18 (.D(integrator_tmp[18]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i17 (.D(integrator_tmp[17]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i16 (.D(integrator_tmp[16]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i15 (.D(integrator_tmp[15]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i14 (.D(integrator_tmp[14]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i13 (.D(integrator_tmp[13]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i12 (.D(integrator_tmp[12]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i11 (.D(integrator_tmp[11]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i10 (.D(integrator_tmp[10]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i9 (.D(integrator_tmp[9]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i8 (.D(integrator_tmp[8]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i7 (.D(integrator_tmp[7]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i7.GSR = "ENABLED";
    LUT4 comb10_71__I_0_77_i138_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n68), .D(\comb10[66] ), .Z(n138)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i138_3_lut_4_lut.init = 16'hf960;
    FD1P3AX integrator_d_tmp_i0_i6 (.D(integrator_tmp[6]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i6.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(n67_adj_228[11]), .B(n73), .Z(count_11__N_1980[11])) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    FD1P3AX integrator_d_tmp_i0_i5 (.D(integrator_tmp[5]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i4 (.D(integrator_tmp[4]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i4.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_196 (.A(n20283), .B(n73), .Z(n14270)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_196.init = 16'hbbbb;
    LUT4 i1_4_lut (.A(n18858), .B(count[0]), .C(n18842), .D(count[11]), 
         .Z(decimation_clk_N_2353)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam i1_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_197 (.A(count[9]), .B(n18854), .C(n18840), .D(count[5]), 
         .Z(n18858)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam i1_4_lut_adj_197.init = 16'h8000;
    FD1S3IX count__i11 (.D(count_11__N_1980[11]), .CK(clk_80mhz), .CD(clk_80mhz_enable_1456), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n67_adj_228[9]), .CK(clk_80mhz), .CD(n14270), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n67_adj_228[8]), .CK(clk_80mhz), .CD(n14270), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n67_adj_228[7]), .CK(clk_80mhz), .CD(n14270), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n67_adj_228[6]), .CK(clk_80mhz), .CD(n14270), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n67_adj_228[5]), .CK(clk_80mhz), .CD(n14270), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n67_adj_228[4]), .CK(clk_80mhz), .CD(n14270), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n67_adj_228[3]), .CK(clk_80mhz), .CD(n14270), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(n67_adj_228[2]), .CK(clk_80mhz), .CD(n14270), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(n67_adj_228[1]), .CK(clk_80mhz), .CD(n14270), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i1.GSR = "ENABLED";
    FD1S3AX integrator1_i71 (.D(integrator1_71__N_960[71]), .CK(clk_80mhz), 
            .Q(integrator1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i71.GSR = "ENABLED";
    LUT4 mux_3408_i16_3_lut (.A(n76), .B(n78), .C(cout), .Z(comb10_71__N_2281[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i16_3_lut.init = 16'hcaca;
    FD1S3AX integrator1_i70 (.D(integrator1_71__N_960[70]), .CK(clk_80mhz), 
            .Q(integrator1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i70.GSR = "ENABLED";
    FD1S3AX integrator1_i69 (.D(integrator1_71__N_960[69]), .CK(clk_80mhz), 
            .Q(integrator1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i69.GSR = "ENABLED";
    FD1S3AX integrator1_i68 (.D(integrator1_71__N_960[68]), .CK(clk_80mhz), 
            .Q(integrator1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i68.GSR = "ENABLED";
    FD1S3AX integrator1_i67 (.D(integrator1_71__N_960[67]), .CK(clk_80mhz), 
            .Q(integrator1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i67.GSR = "ENABLED";
    FD1S3AX integrator1_i66 (.D(integrator1_71__N_960[66]), .CK(clk_80mhz), 
            .Q(integrator1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i66.GSR = "ENABLED";
    FD1S3AX integrator1_i65 (.D(integrator1_71__N_960[65]), .CK(clk_80mhz), 
            .Q(integrator1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i65.GSR = "ENABLED";
    FD1S3AX integrator1_i64 (.D(integrator1_71__N_960[64]), .CK(clk_80mhz), 
            .Q(integrator1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i64.GSR = "ENABLED";
    FD1S3AX integrator1_i63 (.D(integrator1_71__N_960[63]), .CK(clk_80mhz), 
            .Q(integrator1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i63.GSR = "ENABLED";
    FD1S3AX integrator1_i62 (.D(integrator1_71__N_960[62]), .CK(clk_80mhz), 
            .Q(integrator1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i62.GSR = "ENABLED";
    FD1S3AX integrator1_i61 (.D(integrator1_71__N_960[61]), .CK(clk_80mhz), 
            .Q(integrator1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i61.GSR = "ENABLED";
    FD1S3AX integrator1_i60 (.D(integrator1_71__N_960[60]), .CK(clk_80mhz), 
            .Q(integrator1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i60.GSR = "ENABLED";
    FD1S3AX integrator1_i59 (.D(integrator1_71__N_960[59]), .CK(clk_80mhz), 
            .Q(integrator1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i59.GSR = "ENABLED";
    FD1S3AX integrator1_i58 (.D(integrator1_71__N_960[58]), .CK(clk_80mhz), 
            .Q(integrator1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i58.GSR = "ENABLED";
    FD1S3AX integrator1_i57 (.D(integrator1_71__N_960[57]), .CK(clk_80mhz), 
            .Q(integrator1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i57.GSR = "ENABLED";
    FD1S3AX integrator1_i56 (.D(integrator1_71__N_960[56]), .CK(clk_80mhz), 
            .Q(integrator1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i56.GSR = "ENABLED";
    FD1S3AX integrator1_i55 (.D(integrator1_71__N_960[55]), .CK(clk_80mhz), 
            .Q(integrator1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i55.GSR = "ENABLED";
    FD1S3AX integrator1_i54 (.D(integrator1_71__N_960[54]), .CK(clk_80mhz), 
            .Q(integrator1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i54.GSR = "ENABLED";
    FD1S3AX integrator1_i53 (.D(integrator1_71__N_960[53]), .CK(clk_80mhz), 
            .Q(integrator1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i53.GSR = "ENABLED";
    FD1S3AX integrator1_i52 (.D(integrator1_71__N_960[52]), .CK(clk_80mhz), 
            .Q(integrator1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i52.GSR = "ENABLED";
    FD1S3AX integrator1_i51 (.D(integrator1_71__N_960[51]), .CK(clk_80mhz), 
            .Q(integrator1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i51.GSR = "ENABLED";
    FD1S3AX integrator1_i50 (.D(integrator1_71__N_960[50]), .CK(clk_80mhz), 
            .Q(integrator1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i50.GSR = "ENABLED";
    FD1S3AX integrator1_i49 (.D(integrator1_71__N_960[49]), .CK(clk_80mhz), 
            .Q(integrator1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i49.GSR = "ENABLED";
    FD1S3AX integrator1_i48 (.D(integrator1_71__N_960[48]), .CK(clk_80mhz), 
            .Q(integrator1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i48.GSR = "ENABLED";
    FD1S3AX integrator1_i47 (.D(integrator1_71__N_960[47]), .CK(clk_80mhz), 
            .Q(integrator1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i47.GSR = "ENABLED";
    FD1S3AX integrator1_i46 (.D(integrator1_71__N_960[46]), .CK(clk_80mhz), 
            .Q(integrator1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i46.GSR = "ENABLED";
    FD1S3AX integrator1_i45 (.D(integrator1_71__N_960[45]), .CK(clk_80mhz), 
            .Q(integrator1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i45.GSR = "ENABLED";
    FD1S3AX integrator1_i44 (.D(integrator1_71__N_960[44]), .CK(clk_80mhz), 
            .Q(integrator1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i44.GSR = "ENABLED";
    FD1S3AX integrator1_i43 (.D(integrator1_71__N_960[43]), .CK(clk_80mhz), 
            .Q(integrator1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i43.GSR = "ENABLED";
    FD1S3AX integrator1_i42 (.D(integrator1_71__N_960[42]), .CK(clk_80mhz), 
            .Q(integrator1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i42.GSR = "ENABLED";
    FD1S3AX integrator1_i41 (.D(integrator1_71__N_960[41]), .CK(clk_80mhz), 
            .Q(integrator1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i41.GSR = "ENABLED";
    FD1S3AX integrator1_i40 (.D(integrator1_71__N_960[40]), .CK(clk_80mhz), 
            .Q(integrator1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i40.GSR = "ENABLED";
    FD1S3AX integrator1_i39 (.D(integrator1_71__N_960[39]), .CK(clk_80mhz), 
            .Q(integrator1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i39.GSR = "ENABLED";
    FD1S3AX integrator1_i38 (.D(integrator1_71__N_960[38]), .CK(clk_80mhz), 
            .Q(integrator1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i38.GSR = "ENABLED";
    FD1S3AX integrator1_i37 (.D(integrator1_71__N_960[37]), .CK(clk_80mhz), 
            .Q(integrator1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i37.GSR = "ENABLED";
    FD1S3AX integrator1_i36 (.D(integrator1_71__N_960[36]), .CK(clk_80mhz), 
            .Q(integrator1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i36.GSR = "ENABLED";
    FD1S3AX integrator1_i35 (.D(integrator1_71__N_960[35]), .CK(clk_80mhz), 
            .Q(integrator1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i35.GSR = "ENABLED";
    FD1S3AX integrator1_i34 (.D(integrator1_71__N_960[34]), .CK(clk_80mhz), 
            .Q(integrator1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i34.GSR = "ENABLED";
    FD1S3AX integrator1_i33 (.D(integrator1_71__N_960[33]), .CK(clk_80mhz), 
            .Q(integrator1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i33.GSR = "ENABLED";
    FD1S3AX integrator1_i32 (.D(integrator1_71__N_960[32]), .CK(clk_80mhz), 
            .Q(integrator1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i32.GSR = "ENABLED";
    FD1S3AX integrator1_i31 (.D(integrator1_71__N_960[31]), .CK(clk_80mhz), 
            .Q(integrator1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i31.GSR = "ENABLED";
    FD1S3AX integrator1_i30 (.D(integrator1_71__N_960[30]), .CK(clk_80mhz), 
            .Q(integrator1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i30.GSR = "ENABLED";
    FD1S3AX integrator1_i29 (.D(integrator1_71__N_960[29]), .CK(clk_80mhz), 
            .Q(integrator1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i29.GSR = "ENABLED";
    FD1S3AX integrator1_i28 (.D(integrator1_71__N_960[28]), .CK(clk_80mhz), 
            .Q(integrator1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i28.GSR = "ENABLED";
    FD1S3AX integrator1_i27 (.D(integrator1_71__N_960[27]), .CK(clk_80mhz), 
            .Q(integrator1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i27.GSR = "ENABLED";
    FD1S3AX integrator1_i26 (.D(integrator1_71__N_960[26]), .CK(clk_80mhz), 
            .Q(integrator1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i26.GSR = "ENABLED";
    FD1S3AX integrator1_i25 (.D(integrator1_71__N_960[25]), .CK(clk_80mhz), 
            .Q(integrator1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i25.GSR = "ENABLED";
    FD1S3AX integrator1_i24 (.D(integrator1_71__N_960[24]), .CK(clk_80mhz), 
            .Q(integrator1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i24.GSR = "ENABLED";
    FD1S3AX integrator1_i23 (.D(integrator1_71__N_960[23]), .CK(clk_80mhz), 
            .Q(integrator1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i23.GSR = "ENABLED";
    FD1S3AX integrator1_i22 (.D(integrator1_71__N_960[22]), .CK(clk_80mhz), 
            .Q(integrator1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i22.GSR = "ENABLED";
    FD1S3AX integrator1_i21 (.D(integrator1_71__N_960[21]), .CK(clk_80mhz), 
            .Q(integrator1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i21.GSR = "ENABLED";
    FD1S3AX integrator1_i20 (.D(integrator1_71__N_960[20]), .CK(clk_80mhz), 
            .Q(integrator1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i20.GSR = "ENABLED";
    FD1S3AX integrator1_i19 (.D(integrator1_71__N_960[19]), .CK(clk_80mhz), 
            .Q(integrator1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i19.GSR = "ENABLED";
    FD1S3AX integrator1_i18 (.D(integrator1_71__N_960[18]), .CK(clk_80mhz), 
            .Q(integrator1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i18.GSR = "ENABLED";
    FD1S3AX integrator1_i17 (.D(integrator1_71__N_960[17]), .CK(clk_80mhz), 
            .Q(integrator1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i17.GSR = "ENABLED";
    FD1S3AX integrator1_i16 (.D(integrator1_71__N_960[16]), .CK(clk_80mhz), 
            .Q(integrator1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i16.GSR = "ENABLED";
    FD1S3AX integrator1_i15 (.D(integrator1_71__N_960[15]), .CK(clk_80mhz), 
            .Q(integrator1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i15.GSR = "ENABLED";
    FD1S3AX integrator1_i14 (.D(integrator1_71__N_960[14]), .CK(clk_80mhz), 
            .Q(integrator1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i14.GSR = "ENABLED";
    FD1S3AX integrator1_i13 (.D(integrator1_71__N_960[13]), .CK(clk_80mhz), 
            .Q(integrator1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i13.GSR = "ENABLED";
    FD1S3AX integrator1_i12 (.D(integrator1_71__N_960[12]), .CK(clk_80mhz), 
            .Q(integrator1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i12.GSR = "ENABLED";
    FD1S3AX integrator1_i11 (.D(integrator1_71__N_960[11]), .CK(clk_80mhz), 
            .Q(integrator1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i11.GSR = "ENABLED";
    FD1S3AX integrator1_i10 (.D(integrator1_71__N_960[10]), .CK(clk_80mhz), 
            .Q(integrator1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i10.GSR = "ENABLED";
    FD1S3AX integrator1_i9 (.D(integrator1_71__N_960[9]), .CK(clk_80mhz), 
            .Q(integrator1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i9.GSR = "ENABLED";
    FD1S3AX integrator1_i8 (.D(integrator1_71__N_960[8]), .CK(clk_80mhz), 
            .Q(integrator1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i8.GSR = "ENABLED";
    FD1S3AX integrator1_i7 (.D(integrator1_71__N_960[7]), .CK(clk_80mhz), 
            .Q(integrator1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i7.GSR = "ENABLED";
    FD1S3AX integrator1_i6 (.D(integrator1_71__N_960[6]), .CK(clk_80mhz), 
            .Q(integrator1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i6.GSR = "ENABLED";
    FD1S3AX integrator1_i5 (.D(integrator1_71__N_960[5]), .CK(clk_80mhz), 
            .Q(integrator1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i5.GSR = "ENABLED";
    FD1S3AX integrator1_i4 (.D(integrator1_71__N_960[4]), .CK(clk_80mhz), 
            .Q(integrator1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i4.GSR = "ENABLED";
    FD1S3AX integrator1_i3 (.D(integrator1_71__N_960[3]), .CK(clk_80mhz), 
            .Q(integrator1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i3.GSR = "ENABLED";
    FD1S3AX integrator1_i2 (.D(integrator1_71__N_960[2]), .CK(clk_80mhz), 
            .Q(integrator1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i2.GSR = "ENABLED";
    FD1S3AX integrator1_i1 (.D(integrator1_71__N_960[1]), .CK(clk_80mhz), 
            .Q(integrator1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i1.GSR = "ENABLED";
    LUT4 mux_3408_i15_3_lut (.A(n79), .B(n81), .C(cout), .Z(comb10_71__N_2281[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i15_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_198 (.A(count[7]), .B(count[4]), .Z(n18842)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam i1_2_lut_adj_198.init = 16'h8888;
    LUT4 comb10_71__I_0_77_i131_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n61), .D(comb10[59]), .Z(n131)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i131_3_lut_4_lut.init = 16'hf960;
    LUT4 i1_4_lut_adj_199 (.A(count[3]), .B(count[2]), .C(count[10]), 
         .D(count[6]), .Z(n18854)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam i1_4_lut_adj_199.init = 16'h8000;
    LUT4 mux_3408_i14_3_lut (.A(n82), .B(n84), .C(cout), .Z(comb10_71__N_2281[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i14_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_200 (.A(count[1]), .B(count[8]), .Z(n18840)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam i1_2_lut_adj_200.init = 16'h8888;
    LUT4 i1_2_lut_adj_201 (.A(n73), .B(decimation_clk), .Z(n14240)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(65[35:40])
    defparam i1_2_lut_adj_201.init = 16'h8888;
    FD1P3AX comb10__i16 (.D(comb10_71__N_2281[71]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i16.GSR = "ENABLED";
    FD1P3AX comb10__i15 (.D(comb10_71__N_2281[70]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i15.GSR = "ENABLED";
    FD1P3AX comb10__i14 (.D(comb10_71__N_2281[69]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i14.GSR = "ENABLED";
    FD1P3AX comb10__i13 (.D(comb10_71__N_2281[68]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i13.GSR = "ENABLED";
    FD1P3AX comb10__i12 (.D(comb10_71__N_2281[67]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i12.GSR = "ENABLED";
    FD1P3AX comb10__i11 (.D(comb10_71__N_2281[66]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i11.GSR = "ENABLED";
    FD1P3AX comb10__i10 (.D(comb10_71__N_2281[65]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i10.GSR = "ENABLED";
    FD1P3AX comb10__i9 (.D(comb10_71__N_2281[64]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i9.GSR = "ENABLED";
    FD1P3AX comb10__i8 (.D(comb10_71__N_2281[63]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i8.GSR = "ENABLED";
    FD1P3AX comb10__i7 (.D(comb10_71__N_2281[62]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i7.GSR = "ENABLED";
    FD1P3AX comb10__i6 (.D(comb10_71__N_2281[61]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i6.GSR = "ENABLED";
    FD1P3AX comb10__i5 (.D(comb10_71__N_2281[60]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i5.GSR = "ENABLED";
    FD1P3AX comb10__i4 (.D(comb10_71__N_2281[59]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i4.GSR = "ENABLED";
    FD1P3AX comb10__i3 (.D(comb10_71__N_2281[58]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i3.GSR = "ENABLED";
    FD1P3AX comb10__i2 (.D(comb10_71__N_2281[57]), .SP(clk_80mhz_enable_873), 
            .CK(clk_80mhz), .Q(comb10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i2.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i71 (.D(comb9[71]), .SP(clk_80mhz_enable_873), .CK(clk_80mhz), 
            .Q(comb_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i70 (.D(comb9[70]), .SP(clk_80mhz_enable_873), .CK(clk_80mhz), 
            .Q(comb_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i69 (.D(comb9[69]), .SP(clk_80mhz_enable_873), .CK(clk_80mhz), 
            .Q(comb_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i68 (.D(comb9[68]), .SP(clk_80mhz_enable_873), .CK(clk_80mhz), 
            .Q(comb_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i67 (.D(comb9[67]), .SP(clk_80mhz_enable_873), .CK(clk_80mhz), 
            .Q(comb_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i66 (.D(comb9[66]), .SP(clk_80mhz_enable_873), .CK(clk_80mhz), 
            .Q(comb_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i66.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_202 (.A(count[11]), .B(n18796), .C(n18780), .D(n18788), 
         .Z(n73)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_202.init = 16'hfffd;
    FD1P3AX comb_d9_i0_i65 (.D(comb9[65]), .SP(clk_80mhz_enable_873), .CK(clk_80mhz), 
            .Q(comb_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i64 (.D(comb9[64]), .SP(clk_80mhz_enable_873), .CK(clk_80mhz), 
            .Q(comb_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i63 (.D(comb9[63]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i62 (.D(comb9[62]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i61 (.D(comb9[61]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i60 (.D(comb9[60]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i59 (.D(comb9[59]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i58 (.D(comb9[58]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i57 (.D(comb9[57]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i56 (.D(comb9[56]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i55 (.D(comb9[55]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i54 (.D(comb9[54]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i53 (.D(comb9[53]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i52 (.D(comb9[52]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i51 (.D(comb9[51]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i50 (.D(comb9[50]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i49 (.D(comb9[49]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i48 (.D(comb9[48]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i47 (.D(comb9[47]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i46 (.D(comb9[46]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i45 (.D(comb9[45]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i44 (.D(comb9[44]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i43 (.D(comb9[43]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i42 (.D(comb9[42]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i41 (.D(comb9[41]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i40 (.D(comb9[40]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i39 (.D(comb9[39]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i38 (.D(comb9[38]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i37 (.D(comb9[37]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i36 (.D(comb9[36]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i35 (.D(comb9[35]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i34 (.D(comb9[34]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i33 (.D(comb9[33]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i32 (.D(comb9[32]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i31 (.D(comb9[31]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i30 (.D(comb9[30]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i29 (.D(comb9[29]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i28 (.D(comb9[28]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i27 (.D(comb9[27]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i26 (.D(comb9[26]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i3 (.D(integrator_tmp[3]), .SP(clk_80mhz_enable_923), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i25 (.D(comb9[25]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i24 (.D(comb9[24]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i24.GSR = "ENABLED";
    LUT4 mux_3408_i13_3_lut (.A(n85), .B(n87), .C(cout), .Z(comb10_71__N_2281[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i13_3_lut.init = 16'hcaca;
    FD1P3AX comb_d9_i0_i23 (.D(comb9[23]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i22 (.D(comb9[22]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i21 (.D(comb9[21]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i20 (.D(comb9[20]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i19 (.D(comb9[19]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i18 (.D(comb9[18]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i17 (.D(comb9[17]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i2 (.D(integrator_tmp[2]), .SP(clk_80mhz_enable_923), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i16 (.D(comb9[16]), .SP(clk_80mhz_enable_923), .CK(clk_80mhz), 
            .Q(comb_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i15 (.D(comb9[15]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i14 (.D(comb9[14]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i13 (.D(comb9[13]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i12 (.D(comb9[12]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i11 (.D(comb9[11]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i10 (.D(comb9[10]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i9 (.D(comb9[9]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i8 (.D(comb9[8]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i7 (.D(comb9[7]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i6 (.D(comb9[6]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i5 (.D(comb9[5]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i4 (.D(comb9[4]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i3 (.D(comb9[3]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i2 (.D(comb9[2]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i1 (.D(comb9[1]), .SP(clk_80mhz_enable_973), .CK(clk_80mhz), 
            .Q(comb_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i1 (.D(integrator_tmp[1]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX comb9_i0_i71 (.D(comb9_71__N_2209[71]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i71.GSR = "ENABLED";
    FD1P3AX comb9_i0_i70 (.D(comb9_71__N_2209[70]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i70.GSR = "ENABLED";
    FD1P3AX comb9_i0_i69 (.D(comb9_71__N_2209[69]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i69.GSR = "ENABLED";
    FD1P3AX comb9_i0_i68 (.D(comb9_71__N_2209[68]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i68.GSR = "ENABLED";
    FD1P3AX comb9_i0_i67 (.D(comb9_71__N_2209[67]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i67.GSR = "ENABLED";
    FD1P3AX comb9_i0_i66 (.D(comb9_71__N_2209[66]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i66.GSR = "ENABLED";
    FD1P3AX comb9_i0_i65 (.D(comb9_71__N_2209[65]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i65.GSR = "ENABLED";
    FD1P3AX comb9_i0_i64 (.D(comb9_71__N_2209[64]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i64.GSR = "ENABLED";
    FD1P3AX comb9_i0_i63 (.D(comb9_71__N_2209[63]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i63.GSR = "ENABLED";
    FD1P3AX comb9_i0_i62 (.D(comb9_71__N_2209[62]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i62.GSR = "ENABLED";
    FD1P3AX comb9_i0_i61 (.D(comb9_71__N_2209[61]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i61.GSR = "ENABLED";
    FD1P3AX comb9_i0_i60 (.D(comb9_71__N_2209[60]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i60.GSR = "ENABLED";
    FD1P3AX comb9_i0_i59 (.D(comb9_71__N_2209[59]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i59.GSR = "ENABLED";
    FD1P3AX comb9_i0_i58 (.D(comb9_71__N_2209[58]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i58.GSR = "ENABLED";
    FD1P3AX comb9_i0_i57 (.D(comb9_71__N_2209[57]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i57.GSR = "ENABLED";
    FD1P3AX comb9_i0_i56 (.D(comb9_71__N_2209[56]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i56.GSR = "ENABLED";
    FD1P3AX comb9_i0_i55 (.D(comb9_71__N_2209[55]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i55.GSR = "ENABLED";
    FD1P3AX comb9_i0_i54 (.D(comb9_71__N_2209[54]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i54.GSR = "ENABLED";
    FD1P3AX comb9_i0_i53 (.D(comb9_71__N_2209[53]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i53.GSR = "ENABLED";
    FD1P3AX comb9_i0_i52 (.D(comb9_71__N_2209[52]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i52.GSR = "ENABLED";
    FD1P3AX comb9_i0_i51 (.D(comb9_71__N_2209[51]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i51.GSR = "ENABLED";
    FD1P3AX comb9_i0_i50 (.D(comb9_71__N_2209[50]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i50.GSR = "ENABLED";
    FD1P3AX comb9_i0_i49 (.D(comb9_71__N_2209[49]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i49.GSR = "ENABLED";
    FD1P3AX comb9_i0_i48 (.D(comb9_71__N_2209[48]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i48.GSR = "ENABLED";
    FD1P3AX comb9_i0_i47 (.D(comb9_71__N_2209[47]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i47.GSR = "ENABLED";
    FD1P3AX comb9_i0_i46 (.D(comb9_71__N_2209[46]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i46.GSR = "ENABLED";
    FD1P3AX comb9_i0_i45 (.D(comb9_71__N_2209[45]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i45.GSR = "ENABLED";
    FD1P3AX comb9_i0_i44 (.D(comb9_71__N_2209[44]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i44.GSR = "ENABLED";
    FD1P3AX comb9_i0_i43 (.D(comb9_71__N_2209[43]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i43.GSR = "ENABLED";
    FD1P3AX comb9_i0_i42 (.D(comb9_71__N_2209[42]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i42.GSR = "ENABLED";
    FD1P3AX comb9_i0_i41 (.D(comb9_71__N_2209[41]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i41.GSR = "ENABLED";
    FD1P3AX comb9_i0_i40 (.D(comb9_71__N_2209[40]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i40.GSR = "ENABLED";
    FD1P3AX comb9_i0_i39 (.D(comb9_71__N_2209[39]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i39.GSR = "ENABLED";
    FD1P3AX comb9_i0_i38 (.D(comb9_71__N_2209[38]), .SP(clk_80mhz_enable_973), 
            .CK(clk_80mhz), .Q(comb9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i38.GSR = "ENABLED";
    FD1P3AX comb9_i0_i37 (.D(comb9_71__N_2209[37]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i37.GSR = "ENABLED";
    FD1P3AX comb9_i0_i36 (.D(comb9_71__N_2209[36]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i36.GSR = "ENABLED";
    FD1P3AX comb9_i0_i35 (.D(comb9_71__N_2209[35]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i35.GSR = "ENABLED";
    FD1P3AX comb9_i0_i34 (.D(comb9_71__N_2209[34]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i34.GSR = "ENABLED";
    FD1P3AX comb9_i0_i33 (.D(comb9_71__N_2209[33]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i33.GSR = "ENABLED";
    FD1P3AX comb9_i0_i32 (.D(comb9_71__N_2209[32]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i32.GSR = "ENABLED";
    FD1P3AX comb9_i0_i31 (.D(comb9_71__N_2209[31]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i31.GSR = "ENABLED";
    FD1P3AX comb9_i0_i30 (.D(comb9_71__N_2209[30]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i30.GSR = "ENABLED";
    FD1P3AX comb9_i0_i29 (.D(comb9_71__N_2209[29]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i29.GSR = "ENABLED";
    FD1P3AX comb9_i0_i28 (.D(comb9_71__N_2209[28]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i28.GSR = "ENABLED";
    FD1P3AX comb9_i0_i27 (.D(comb9_71__N_2209[27]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i27.GSR = "ENABLED";
    FD1P3AX comb9_i0_i26 (.D(comb9_71__N_2209[26]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i26.GSR = "ENABLED";
    FD1P3AX comb9_i0_i25 (.D(comb9_71__N_2209[25]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i25.GSR = "ENABLED";
    FD1P3AX comb9_i0_i24 (.D(comb9_71__N_2209[24]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i24.GSR = "ENABLED";
    FD1P3AX comb9_i0_i23 (.D(comb9_71__N_2209[23]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i23.GSR = "ENABLED";
    FD1P3AX comb9_i0_i22 (.D(comb9_71__N_2209[22]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i22.GSR = "ENABLED";
    FD1P3AX comb9_i0_i21 (.D(comb9_71__N_2209[21]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i21.GSR = "ENABLED";
    FD1P3AX comb9_i0_i20 (.D(comb9_71__N_2209[20]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i20.GSR = "ENABLED";
    FD1P3AX comb9_i0_i19 (.D(comb9_71__N_2209[19]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i19.GSR = "ENABLED";
    FD1P3AX comb9_i0_i18 (.D(comb9_71__N_2209[18]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i18.GSR = "ENABLED";
    FD1P3AX comb9_i0_i17 (.D(comb9_71__N_2209[17]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i17.GSR = "ENABLED";
    FD1P3AX comb9_i0_i16 (.D(comb9_71__N_2209[16]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i16.GSR = "ENABLED";
    FD1P3AX comb9_i0_i15 (.D(comb9_71__N_2209[15]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i15.GSR = "ENABLED";
    FD1P3AX comb9_i0_i14 (.D(comb9_71__N_2209[14]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i14.GSR = "ENABLED";
    FD1P3AX comb9_i0_i13 (.D(comb9_71__N_2209[13]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i13.GSR = "ENABLED";
    FD1P3AX comb9_i0_i12 (.D(comb9_71__N_2209[12]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i12.GSR = "ENABLED";
    FD1P3AX comb9_i0_i11 (.D(comb9_71__N_2209[11]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i11.GSR = "ENABLED";
    FD1P3AX comb9_i0_i10 (.D(comb9_71__N_2209[10]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i10.GSR = "ENABLED";
    FD1P3AX comb9_i0_i9 (.D(comb9_71__N_2209[9]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i9.GSR = "ENABLED";
    FD1P3AX comb9_i0_i8 (.D(comb9_71__N_2209[8]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i8.GSR = "ENABLED";
    FD1P3AX comb9_i0_i7 (.D(comb9_71__N_2209[7]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i7.GSR = "ENABLED";
    FD1P3AX comb9_i0_i6 (.D(comb9_71__N_2209[6]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i6.GSR = "ENABLED";
    FD1P3AX comb9_i0_i5 (.D(comb9_71__N_2209[5]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i5.GSR = "ENABLED";
    FD1P3AX comb9_i0_i4 (.D(comb9_71__N_2209[4]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i4.GSR = "ENABLED";
    FD1P3AX comb9_i0_i3 (.D(comb9_71__N_2209[3]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i3.GSR = "ENABLED";
    FD1P3AX comb9_i0_i2 (.D(comb9_71__N_2209[2]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i2.GSR = "ENABLED";
    FD1P3AX comb9_i0_i1 (.D(comb9_71__N_2209[1]), .SP(clk_80mhz_enable_1023), 
            .CK(clk_80mhz), .Q(comb9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i71 (.D(comb8[71]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i70 (.D(comb8[70]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i69 (.D(comb8[69]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i68 (.D(comb8[68]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i67 (.D(comb8[67]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i66 (.D(comb8[66]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i65 (.D(comb8[65]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i64 (.D(comb8[64]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i63 (.D(comb8[63]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i62 (.D(comb8[62]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i61 (.D(comb8[61]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i60 (.D(comb8[60]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i59 (.D(comb8[59]), .SP(clk_80mhz_enable_1023), .CK(clk_80mhz), 
            .Q(comb_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i58 (.D(comb8[58]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i57 (.D(comb8[57]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i56 (.D(comb8[56]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i55 (.D(comb8[55]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i54 (.D(comb8[54]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i53 (.D(comb8[53]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i52 (.D(comb8[52]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i51 (.D(comb8[51]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i50 (.D(comb8[50]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i49 (.D(comb8[49]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i48 (.D(comb8[48]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i47 (.D(comb8[47]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i46 (.D(comb8[46]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i45 (.D(comb8[45]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i44 (.D(comb8[44]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i43 (.D(comb8[43]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i42 (.D(comb8[42]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i41 (.D(comb8[41]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i40 (.D(comb8[40]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i39 (.D(comb8[39]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i38 (.D(comb8[38]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i37 (.D(comb8[37]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i36 (.D(comb8[36]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i35 (.D(comb8[35]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i34 (.D(comb8[34]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i33 (.D(comb8[33]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i32 (.D(comb8[32]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i31 (.D(comb8[31]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i30 (.D(comb8[30]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i29 (.D(comb8[29]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i28 (.D(comb8[28]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i27 (.D(comb8[27]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i26 (.D(comb8[26]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i25 (.D(comb8[25]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i24 (.D(comb8[24]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i23 (.D(comb8[23]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i22 (.D(comb8[22]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i21 (.D(comb8[21]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i20 (.D(comb8[20]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i19 (.D(comb8[19]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i18 (.D(comb8[18]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i17 (.D(comb8[17]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i16 (.D(comb8[16]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i15 (.D(comb8[15]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i14 (.D(comb8[14]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i13 (.D(comb8[13]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i12 (.D(comb8[12]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i11 (.D(comb8[11]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i10 (.D(comb8[10]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i9 (.D(comb8[9]), .SP(clk_80mhz_enable_1073), .CK(clk_80mhz), 
            .Q(comb_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i8 (.D(comb8[8]), .SP(clk_80mhz_enable_1123), .CK(clk_80mhz), 
            .Q(comb_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i7 (.D(comb8[7]), .SP(clk_80mhz_enable_1123), .CK(clk_80mhz), 
            .Q(comb_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i6 (.D(comb8[6]), .SP(clk_80mhz_enable_1123), .CK(clk_80mhz), 
            .Q(comb_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i5 (.D(comb8[5]), .SP(clk_80mhz_enable_1123), .CK(clk_80mhz), 
            .Q(comb_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i4 (.D(comb8[4]), .SP(clk_80mhz_enable_1123), .CK(clk_80mhz), 
            .Q(comb_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i3 (.D(comb8[3]), .SP(clk_80mhz_enable_1123), .CK(clk_80mhz), 
            .Q(comb_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i2 (.D(comb8[2]), .SP(clk_80mhz_enable_1123), .CK(clk_80mhz), 
            .Q(comb_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i1 (.D(comb8[1]), .SP(clk_80mhz_enable_1123), .CK(clk_80mhz), 
            .Q(comb_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX comb8_i0_i71 (.D(comb8_71__N_2137[71]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i71.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_203 (.A(count[4]), .B(n18792), .C(count[9]), .D(count[1]), 
         .Z(n18796)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_203.init = 16'hfffe;
    LUT4 mux_3408_i12_3_lut (.A(n88), .B(n90), .C(cout), .Z(comb10_71__N_2281[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i12_3_lut.init = 16'hcaca;
    FD1P3AX comb8_i0_i70 (.D(comb8_71__N_2137[70]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i70.GSR = "ENABLED";
    FD1P3AX comb8_i0_i69 (.D(comb8_71__N_2137[69]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i69.GSR = "ENABLED";
    FD1P3AX comb8_i0_i68 (.D(comb8_71__N_2137[68]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i68.GSR = "ENABLED";
    FD1P3AX comb8_i0_i67 (.D(comb8_71__N_2137[67]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i67.GSR = "ENABLED";
    FD1P3AX comb8_i0_i66 (.D(comb8_71__N_2137[66]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i66.GSR = "ENABLED";
    FD1P3AX comb8_i0_i65 (.D(comb8_71__N_2137[65]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i65.GSR = "ENABLED";
    FD1P3AX comb8_i0_i64 (.D(comb8_71__N_2137[64]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i64.GSR = "ENABLED";
    FD1P3AX comb8_i0_i63 (.D(comb8_71__N_2137[63]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i63.GSR = "ENABLED";
    FD1P3AX comb8_i0_i62 (.D(comb8_71__N_2137[62]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i62.GSR = "ENABLED";
    FD1P3AX comb8_i0_i61 (.D(comb8_71__N_2137[61]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i61.GSR = "ENABLED";
    FD1P3AX comb8_i0_i60 (.D(comb8_71__N_2137[60]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i60.GSR = "ENABLED";
    FD1P3AX comb8_i0_i59 (.D(comb8_71__N_2137[59]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i59.GSR = "ENABLED";
    FD1P3AX comb8_i0_i58 (.D(comb8_71__N_2137[58]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i58.GSR = "ENABLED";
    FD1P3AX comb8_i0_i57 (.D(comb8_71__N_2137[57]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i57.GSR = "ENABLED";
    FD1P3AX comb8_i0_i56 (.D(comb8_71__N_2137[56]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i56.GSR = "ENABLED";
    FD1P3AX comb8_i0_i55 (.D(comb8_71__N_2137[55]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i55.GSR = "ENABLED";
    FD1P3AX comb8_i0_i54 (.D(comb8_71__N_2137[54]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i54.GSR = "ENABLED";
    FD1P3AX comb8_i0_i53 (.D(comb8_71__N_2137[53]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i53.GSR = "ENABLED";
    FD1P3AX comb8_i0_i52 (.D(comb8_71__N_2137[52]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i52.GSR = "ENABLED";
    FD1P3AX comb8_i0_i51 (.D(comb8_71__N_2137[51]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i51.GSR = "ENABLED";
    FD1P3AX comb8_i0_i50 (.D(comb8_71__N_2137[50]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i50.GSR = "ENABLED";
    FD1P3AX comb8_i0_i49 (.D(comb8_71__N_2137[49]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i49.GSR = "ENABLED";
    FD1P3AX comb8_i0_i48 (.D(comb8_71__N_2137[48]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i48.GSR = "ENABLED";
    FD1P3AX comb8_i0_i47 (.D(comb8_71__N_2137[47]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i47.GSR = "ENABLED";
    FD1P3AX comb8_i0_i46 (.D(comb8_71__N_2137[46]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i46.GSR = "ENABLED";
    FD1P3AX comb8_i0_i45 (.D(comb8_71__N_2137[45]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i45.GSR = "ENABLED";
    FD1P3AX comb8_i0_i44 (.D(comb8_71__N_2137[44]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i44.GSR = "ENABLED";
    FD1P3AX comb8_i0_i43 (.D(comb8_71__N_2137[43]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i43.GSR = "ENABLED";
    FD1P3AX comb8_i0_i42 (.D(comb8_71__N_2137[42]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i42.GSR = "ENABLED";
    FD1P3AX comb8_i0_i41 (.D(comb8_71__N_2137[41]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i41.GSR = "ENABLED";
    FD1P3AX comb8_i0_i40 (.D(comb8_71__N_2137[40]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i40.GSR = "ENABLED";
    FD1P3AX comb8_i0_i39 (.D(comb8_71__N_2137[39]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i39.GSR = "ENABLED";
    FD1P3AX comb8_i0_i38 (.D(comb8_71__N_2137[38]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i38.GSR = "ENABLED";
    FD1P3AX comb8_i0_i37 (.D(comb8_71__N_2137[37]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i37.GSR = "ENABLED";
    FD1P3AX comb8_i0_i36 (.D(comb8_71__N_2137[36]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i36.GSR = "ENABLED";
    FD1P3AX comb8_i0_i35 (.D(comb8_71__N_2137[35]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i35.GSR = "ENABLED";
    FD1P3AX comb8_i0_i34 (.D(comb8_71__N_2137[34]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i34.GSR = "ENABLED";
    FD1P3AX comb8_i0_i33 (.D(comb8_71__N_2137[33]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i33.GSR = "ENABLED";
    FD1P3AX comb8_i0_i32 (.D(comb8_71__N_2137[32]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i32.GSR = "ENABLED";
    FD1P3AX comb8_i0_i31 (.D(comb8_71__N_2137[31]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i31.GSR = "ENABLED";
    FD1P3AX comb8_i0_i30 (.D(comb8_71__N_2137[30]), .SP(clk_80mhz_enable_1123), 
            .CK(clk_80mhz), .Q(comb8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i30.GSR = "ENABLED";
    FD1P3AX comb8_i0_i29 (.D(comb8_71__N_2137[29]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i29.GSR = "ENABLED";
    FD1P3AX comb8_i0_i28 (.D(comb8_71__N_2137[28]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i28.GSR = "ENABLED";
    FD1P3AX comb8_i0_i27 (.D(comb8_71__N_2137[27]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i27.GSR = "ENABLED";
    FD1P3AX comb8_i0_i26 (.D(comb8_71__N_2137[26]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i26.GSR = "ENABLED";
    FD1P3AX comb8_i0_i25 (.D(comb8_71__N_2137[25]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i25.GSR = "ENABLED";
    FD1P3AX comb8_i0_i24 (.D(comb8_71__N_2137[24]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i24.GSR = "ENABLED";
    FD1P3AX comb8_i0_i23 (.D(comb8_71__N_2137[23]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i23.GSR = "ENABLED";
    FD1P3AX comb8_i0_i22 (.D(comb8_71__N_2137[22]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i22.GSR = "ENABLED";
    FD1P3AX comb8_i0_i21 (.D(comb8_71__N_2137[21]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i21.GSR = "ENABLED";
    FD1P3AX comb8_i0_i20 (.D(comb8_71__N_2137[20]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i20.GSR = "ENABLED";
    FD1P3AX comb8_i0_i19 (.D(comb8_71__N_2137[19]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i19.GSR = "ENABLED";
    FD1P3AX comb8_i0_i18 (.D(comb8_71__N_2137[18]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i18.GSR = "ENABLED";
    FD1P3AX comb8_i0_i17 (.D(comb8_71__N_2137[17]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i17.GSR = "ENABLED";
    FD1P3AX comb8_i0_i16 (.D(comb8_71__N_2137[16]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i16.GSR = "ENABLED";
    FD1P3AX comb8_i0_i15 (.D(comb8_71__N_2137[15]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i15.GSR = "ENABLED";
    FD1P3AX comb8_i0_i14 (.D(comb8_71__N_2137[14]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i14.GSR = "ENABLED";
    FD1P3AX comb8_i0_i13 (.D(comb8_71__N_2137[13]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i13.GSR = "ENABLED";
    FD1P3AX comb8_i0_i12 (.D(comb8_71__N_2137[12]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i12.GSR = "ENABLED";
    FD1P3AX comb8_i0_i11 (.D(comb8_71__N_2137[11]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i11.GSR = "ENABLED";
    FD1P3AX comb8_i0_i10 (.D(comb8_71__N_2137[10]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i10.GSR = "ENABLED";
    FD1P3AX comb8_i0_i9 (.D(comb8_71__N_2137[9]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i9.GSR = "ENABLED";
    FD1P3AX comb8_i0_i8 (.D(comb8_71__N_2137[8]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i8.GSR = "ENABLED";
    FD1P3AX comb8_i0_i7 (.D(comb8_71__N_2137[7]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i7.GSR = "ENABLED";
    FD1P3AX comb8_i0_i6 (.D(comb8_71__N_2137[6]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i6.GSR = "ENABLED";
    FD1P3AX comb8_i0_i5 (.D(comb8_71__N_2137[5]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i5.GSR = "ENABLED";
    FD1P3AX comb8_i0_i4 (.D(comb8_71__N_2137[4]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i4.GSR = "ENABLED";
    FD1P3AX comb8_i0_i3 (.D(comb8_71__N_2137[3]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i3.GSR = "ENABLED";
    FD1P3AX comb8_i0_i2 (.D(comb8_71__N_2137[2]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i2.GSR = "ENABLED";
    FD1P3AX comb8_i0_i1 (.D(comb8_71__N_2137[1]), .SP(clk_80mhz_enable_1173), 
            .CK(clk_80mhz), .Q(comb8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i71 (.D(comb7[71]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i70 (.D(comb7[70]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i69 (.D(comb7[69]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i68 (.D(comb7[68]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i67 (.D(comb7[67]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i66 (.D(comb7[66]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i65 (.D(comb7[65]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i64 (.D(comb7[64]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i63 (.D(comb7[63]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i62 (.D(comb7[62]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i61 (.D(comb7[61]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i60 (.D(comb7[60]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i59 (.D(comb7[59]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i59.GSR = "ENABLED";
    LUT4 mux_3408_i11_3_lut (.A(n91), .B(n93), .C(cout), .Z(comb10_71__N_2281[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i11_3_lut.init = 16'hcaca;
    FD1P3AX comb_d7_i0_i58 (.D(comb7[58]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i58.GSR = "ENABLED";
    LUT4 comb10_71__I_0_77_i209_4_lut_4_lut_4_lut (.A(comb10[68]), .B(n137), 
         .C(\cic_gain[0] ), .D(\cic_gain[1] ), .Z(led_0_2)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i209_4_lut_4_lut_4_lut.init = 16'hccca;
    FD1P3AX comb_d7_i0_i57 (.D(comb7[57]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i56 (.D(comb7[56]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i55 (.D(comb7[55]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i54 (.D(comb7[54]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i53 (.D(comb7[53]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i52 (.D(comb7[52]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i51 (.D(comb7[51]), .SP(clk_80mhz_enable_1173), .CK(clk_80mhz), 
            .Q(comb_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i50 (.D(comb7[50]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i49 (.D(comb7[49]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i48 (.D(comb7[48]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i47 (.D(comb7[47]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i46 (.D(comb7[46]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i45 (.D(comb7[45]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i44 (.D(comb7[44]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i43 (.D(comb7[43]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i42 (.D(comb7[42]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i41 (.D(comb7[41]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i40 (.D(comb7[40]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i39 (.D(comb7[39]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i38 (.D(comb7[38]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i37 (.D(comb7[37]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i36 (.D(comb7[36]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i35 (.D(comb7[35]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i34 (.D(comb7[34]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i33 (.D(comb7[33]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i32 (.D(comb7[32]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i31 (.D(comb7[31]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i30 (.D(comb7[30]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i29 (.D(comb7[29]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i28 (.D(comb7[28]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i27 (.D(comb7[27]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i26 (.D(comb7[26]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i25 (.D(comb7[25]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i24 (.D(comb7[24]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i23 (.D(comb7[23]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i22 (.D(comb7[22]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i21 (.D(comb7[21]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i20 (.D(comb7[20]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i19 (.D(comb7[19]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i18 (.D(comb7[18]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i17 (.D(comb7[17]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i17.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_204 (.A(count[7]), .B(count[2]), .Z(n18780)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_204.init = 16'heeee;
    FD1P3AX comb_d7_i0_i16 (.D(comb7[16]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i15 (.D(comb7[15]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i14 (.D(comb7[14]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i13 (.D(comb7[13]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i12 (.D(comb7[12]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i11 (.D(comb7[11]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i10 (.D(comb7[10]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i9 (.D(comb7[9]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i8 (.D(comb7[8]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i7 (.D(comb7[7]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i6 (.D(comb7[6]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i5 (.D(comb7[5]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i4 (.D(comb7[4]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i3 (.D(comb7[3]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i2 (.D(comb7[2]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i1 (.D(comb7[1]), .SP(clk_80mhz_enable_1223), .CK(clk_80mhz), 
            .Q(comb_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX comb7_i0_i71 (.D(comb7_71__N_2065[71]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i71.GSR = "ENABLED";
    FD1P3AX comb7_i0_i70 (.D(comb7_71__N_2065[70]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i70.GSR = "ENABLED";
    FD1P3AX comb7_i0_i69 (.D(comb7_71__N_2065[69]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i69.GSR = "ENABLED";
    FD1P3AX comb7_i0_i68 (.D(comb7_71__N_2065[68]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i68.GSR = "ENABLED";
    FD1P3AX comb7_i0_i67 (.D(comb7_71__N_2065[67]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i67.GSR = "ENABLED";
    FD1P3AX comb7_i0_i66 (.D(comb7_71__N_2065[66]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i66.GSR = "ENABLED";
    FD1P3AX comb7_i0_i65 (.D(comb7_71__N_2065[65]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i65.GSR = "ENABLED";
    FD1P3AX comb7_i0_i64 (.D(comb7_71__N_2065[64]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i64.GSR = "ENABLED";
    FD1P3AX comb7_i0_i63 (.D(comb7_71__N_2065[63]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i63.GSR = "ENABLED";
    FD1P3AX comb7_i0_i62 (.D(comb7_71__N_2065[62]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i62.GSR = "ENABLED";
    FD1P3AX comb7_i0_i61 (.D(comb7_71__N_2065[61]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i61.GSR = "ENABLED";
    FD1P3AX comb7_i0_i60 (.D(comb7_71__N_2065[60]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i60.GSR = "ENABLED";
    FD1P3AX comb7_i0_i59 (.D(comb7_71__N_2065[59]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i59.GSR = "ENABLED";
    FD1P3AX comb7_i0_i58 (.D(comb7_71__N_2065[58]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i58.GSR = "ENABLED";
    FD1P3AX comb7_i0_i57 (.D(comb7_71__N_2065[57]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i57.GSR = "ENABLED";
    FD1P3AX comb7_i0_i56 (.D(comb7_71__N_2065[56]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i56.GSR = "ENABLED";
    FD1P3AX comb7_i0_i55 (.D(comb7_71__N_2065[55]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i55.GSR = "ENABLED";
    FD1P3AX comb7_i0_i54 (.D(comb7_71__N_2065[54]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i54.GSR = "ENABLED";
    FD1P3AX comb7_i0_i53 (.D(comb7_71__N_2065[53]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i53.GSR = "ENABLED";
    FD1P3AX comb7_i0_i52 (.D(comb7_71__N_2065[52]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i52.GSR = "ENABLED";
    FD1P3AX comb7_i0_i51 (.D(comb7_71__N_2065[51]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i51.GSR = "ENABLED";
    FD1P3AX comb7_i0_i50 (.D(comb7_71__N_2065[50]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i50.GSR = "ENABLED";
    FD1P3AX comb7_i0_i49 (.D(comb7_71__N_2065[49]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i49.GSR = "ENABLED";
    FD1P3AX comb7_i0_i48 (.D(comb7_71__N_2065[48]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i48.GSR = "ENABLED";
    FD1P3AX comb7_i0_i47 (.D(comb7_71__N_2065[47]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i47.GSR = "ENABLED";
    FD1P3AX comb7_i0_i46 (.D(comb7_71__N_2065[46]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i46.GSR = "ENABLED";
    FD1P3AX comb7_i0_i45 (.D(comb7_71__N_2065[45]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i45.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_205 (.A(count[8]), .B(count[5]), .Z(n18788)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_205.init = 16'heeee;
    FD1P3AX comb7_i0_i44 (.D(comb7_71__N_2065[44]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i44.GSR = "ENABLED";
    FD1P3AX comb7_i0_i43 (.D(comb7_71__N_2065[43]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i43.GSR = "ENABLED";
    FD1P3AX comb7_i0_i42 (.D(comb7_71__N_2065[42]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i42.GSR = "ENABLED";
    FD1P3AX comb7_i0_i41 (.D(comb7_71__N_2065[41]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i41.GSR = "ENABLED";
    FD1P3AX comb7_i0_i40 (.D(comb7_71__N_2065[40]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i40.GSR = "ENABLED";
    FD1P3AX comb7_i0_i39 (.D(comb7_71__N_2065[39]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i39.GSR = "ENABLED";
    FD1P3AX comb7_i0_i38 (.D(comb7_71__N_2065[38]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i38.GSR = "ENABLED";
    FD1P3AX comb7_i0_i37 (.D(comb7_71__N_2065[37]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i37.GSR = "ENABLED";
    FD1P3AX comb7_i0_i36 (.D(comb7_71__N_2065[36]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i36.GSR = "ENABLED";
    FD1P3AX comb7_i0_i35 (.D(comb7_71__N_2065[35]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i35.GSR = "ENABLED";
    FD1P3AX comb7_i0_i34 (.D(comb7_71__N_2065[34]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i34.GSR = "ENABLED";
    FD1P3AX comb7_i0_i33 (.D(comb7_71__N_2065[33]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i33.GSR = "ENABLED";
    FD1P3AX comb7_i0_i32 (.D(comb7_71__N_2065[32]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i32.GSR = "ENABLED";
    FD1P3AX comb7_i0_i31 (.D(comb7_71__N_2065[31]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i31.GSR = "ENABLED";
    FD1P3AX comb7_i0_i30 (.D(comb7_71__N_2065[30]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i30.GSR = "ENABLED";
    FD1P3AX comb7_i0_i29 (.D(comb7_71__N_2065[29]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i29.GSR = "ENABLED";
    FD1P3AX comb7_i0_i28 (.D(comb7_71__N_2065[28]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i28.GSR = "ENABLED";
    FD1P3AX comb7_i0_i27 (.D(comb7_71__N_2065[27]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i27.GSR = "ENABLED";
    FD1P3AX comb7_i0_i26 (.D(comb7_71__N_2065[26]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i26.GSR = "ENABLED";
    FD1P3AX comb7_i0_i25 (.D(comb7_71__N_2065[25]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i25.GSR = "ENABLED";
    FD1P3AX comb7_i0_i24 (.D(comb7_71__N_2065[24]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i24.GSR = "ENABLED";
    FD1P3AX comb7_i0_i23 (.D(comb7_71__N_2065[23]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i23.GSR = "ENABLED";
    FD1P3AX comb7_i0_i22 (.D(comb7_71__N_2065[22]), .SP(clk_80mhz_enable_1273), 
            .CK(clk_80mhz), .Q(comb7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i22.GSR = "ENABLED";
    FD1P3AX comb7_i0_i21 (.D(comb7_71__N_2065[21]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i21.GSR = "ENABLED";
    FD1P3AX comb7_i0_i20 (.D(comb7_71__N_2065[20]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i20.GSR = "ENABLED";
    FD1P3AX comb7_i0_i19 (.D(comb7_71__N_2065[19]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i19.GSR = "ENABLED";
    FD1P3AX comb7_i0_i18 (.D(comb7_71__N_2065[18]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i18.GSR = "ENABLED";
    FD1P3AX comb7_i0_i17 (.D(comb7_71__N_2065[17]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i17.GSR = "ENABLED";
    FD1P3AX comb7_i0_i16 (.D(comb7_71__N_2065[16]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i16.GSR = "ENABLED";
    FD1P3AX comb7_i0_i15 (.D(comb7_71__N_2065[15]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i15.GSR = "ENABLED";
    FD1P3AX comb7_i0_i14 (.D(comb7_71__N_2065[14]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i14.GSR = "ENABLED";
    FD1P3AX comb7_i0_i13 (.D(comb7_71__N_2065[13]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i13.GSR = "ENABLED";
    FD1P3AX comb7_i0_i12 (.D(comb7_71__N_2065[12]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i12.GSR = "ENABLED";
    FD1P3AX comb7_i0_i11 (.D(comb7_71__N_2065[11]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i11.GSR = "ENABLED";
    FD1P3AX comb7_i0_i10 (.D(comb7_71__N_2065[10]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i10.GSR = "ENABLED";
    FD1P3AX comb7_i0_i9 (.D(comb7_71__N_2065[9]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i9.GSR = "ENABLED";
    FD1P3AX comb7_i0_i8 (.D(comb7_71__N_2065[8]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i8.GSR = "ENABLED";
    FD1P3AX comb7_i0_i7 (.D(comb7_71__N_2065[7]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i7.GSR = "ENABLED";
    FD1P3AX comb7_i0_i6 (.D(comb7_71__N_2065[6]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i6.GSR = "ENABLED";
    FD1P3AX comb7_i0_i5 (.D(comb7_71__N_2065[5]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i5.GSR = "ENABLED";
    FD1P3AX comb7_i0_i4 (.D(comb7_71__N_2065[4]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i4.GSR = "ENABLED";
    FD1P3AX comb7_i0_i3 (.D(comb7_71__N_2065[3]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i3.GSR = "ENABLED";
    FD1P3AX comb7_i0_i2 (.D(comb7_71__N_2065[2]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i2.GSR = "ENABLED";
    FD1P3AX comb7_i0_i1 (.D(comb7_71__N_2065[1]), .SP(clk_80mhz_enable_1323), 
            .CK(clk_80mhz), .Q(comb7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i1.GSR = "ENABLED";
    LUT4 mux_3408_i10_3_lut (.A(n94), .B(n96), .C(cout), .Z(comb10_71__N_2281[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i10_3_lut.init = 16'hcaca;
    FD1P3AX comb_d6_i0_i71 (.D(comb6[71]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i70 (.D(comb6[70]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i69 (.D(comb6[69]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i68 (.D(comb6[68]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i67 (.D(comb6[67]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i66 (.D(comb6[66]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i65 (.D(comb6[65]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i64 (.D(comb6[64]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i63 (.D(comb6[63]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i62 (.D(comb6[62]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i61 (.D(comb6[61]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i60 (.D(comb6[60]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i59 (.D(comb6[59]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i58 (.D(comb6[58]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i57 (.D(comb6[57]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i56 (.D(comb6[56]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i55 (.D(comb6[55]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i54 (.D(comb6[54]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i53 (.D(comb6[53]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i52 (.D(comb6[52]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i51 (.D(comb6[51]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i50 (.D(comb6[50]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i49 (.D(comb6[49]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i48 (.D(comb6[48]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i47 (.D(comb6[47]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i46 (.D(comb6[46]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i45 (.D(comb6[45]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i44 (.D(comb6[44]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i43 (.D(comb6[43]), .SP(clk_80mhz_enable_1323), .CK(clk_80mhz), 
            .Q(comb_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i42 (.D(comb6[42]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i41 (.D(comb6[41]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i40 (.D(comb6[40]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i39 (.D(comb6[39]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i38 (.D(comb6[38]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i37 (.D(comb6[37]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i36 (.D(comb6[36]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i35 (.D(comb6[35]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i34 (.D(comb6[34]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i33 (.D(comb6[33]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i32 (.D(comb6[32]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i31 (.D(comb6[31]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i30 (.D(comb6[30]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i29 (.D(comb6[29]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i28 (.D(comb6[28]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i27 (.D(comb6[27]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i26 (.D(comb6[26]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i25 (.D(comb6[25]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i24 (.D(comb6[24]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i23 (.D(comb6[23]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i22 (.D(comb6[22]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i22.GSR = "ENABLED";
    LUT4 mux_3408_i9_3_lut (.A(n97), .B(n99), .C(cout), .Z(comb10_71__N_2281[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i9_3_lut.init = 16'hcaca;
    FD1P3AX comb_d6_i0_i21 (.D(comb6[21]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i20 (.D(comb6[20]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i19 (.D(comb6[19]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i18 (.D(comb6[18]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i17 (.D(comb6[17]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i16 (.D(comb6[16]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i15 (.D(comb6[15]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i14 (.D(comb6[14]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i13 (.D(comb6[13]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i12 (.D(comb6[12]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i11 (.D(comb6[11]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i10 (.D(comb6[10]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i9 (.D(comb6[9]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i8 (.D(comb6[8]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i7 (.D(comb6[7]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i6 (.D(comb6[6]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i5 (.D(comb6[5]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i4 (.D(comb6[4]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i3 (.D(comb6[3]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i2 (.D(comb6[2]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i1 (.D(comb6[1]), .SP(clk_80mhz_enable_1373), .CK(clk_80mhz), 
            .Q(comb_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX comb6_i0_i71 (.D(comb6_71__N_1993[71]), .SP(clk_80mhz_enable_1373), 
            .CK(clk_80mhz), .Q(comb6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i71.GSR = "ENABLED";
    FD1P3AX comb6_i0_i70 (.D(comb6_71__N_1993[70]), .SP(clk_80mhz_enable_1373), 
            .CK(clk_80mhz), .Q(comb6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i70.GSR = "ENABLED";
    FD1P3AX comb6_i0_i69 (.D(comb6_71__N_1993[69]), .SP(clk_80mhz_enable_1373), 
            .CK(clk_80mhz), .Q(comb6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i69.GSR = "ENABLED";
    FD1P3AX comb6_i0_i68 (.D(comb6_71__N_1993[68]), .SP(clk_80mhz_enable_1373), 
            .CK(clk_80mhz), .Q(comb6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i68.GSR = "ENABLED";
    FD1P3AX comb6_i0_i67 (.D(comb6_71__N_1993[67]), .SP(clk_80mhz_enable_1373), 
            .CK(clk_80mhz), .Q(comb6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i67.GSR = "ENABLED";
    FD1P3AX comb6_i0_i66 (.D(comb6_71__N_1993[66]), .SP(clk_80mhz_enable_1373), 
            .CK(clk_80mhz), .Q(comb6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i66.GSR = "ENABLED";
    FD1P3AX comb6_i0_i65 (.D(comb6_71__N_1993[65]), .SP(clk_80mhz_enable_1373), 
            .CK(clk_80mhz), .Q(comb6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i65.GSR = "ENABLED";
    FD1P3AX comb6_i0_i64 (.D(comb6_71__N_1993[64]), .SP(clk_80mhz_enable_1373), 
            .CK(clk_80mhz), .Q(comb6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i64.GSR = "ENABLED";
    FD1P3AX comb6_i0_i63 (.D(comb6_71__N_1993[63]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i63.GSR = "ENABLED";
    FD1P3AX comb6_i0_i62 (.D(comb6_71__N_1993[62]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i62.GSR = "ENABLED";
    FD1P3AX comb6_i0_i61 (.D(comb6_71__N_1993[61]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i61.GSR = "ENABLED";
    FD1P3AX comb6_i0_i60 (.D(comb6_71__N_1993[60]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i60.GSR = "ENABLED";
    FD1P3AX comb6_i0_i59 (.D(comb6_71__N_1993[59]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i59.GSR = "ENABLED";
    FD1P3AX comb6_i0_i58 (.D(comb6_71__N_1993[58]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i58.GSR = "ENABLED";
    FD1P3AX comb6_i0_i57 (.D(comb6_71__N_1993[57]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i57.GSR = "ENABLED";
    FD1P3AX comb6_i0_i56 (.D(comb6_71__N_1993[56]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i56.GSR = "ENABLED";
    FD1P3AX comb6_i0_i55 (.D(comb6_71__N_1993[55]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i55.GSR = "ENABLED";
    FD1P3AX comb6_i0_i54 (.D(comb6_71__N_1993[54]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i54.GSR = "ENABLED";
    FD1P3AX comb6_i0_i53 (.D(comb6_71__N_1993[53]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i53.GSR = "ENABLED";
    FD1P3AX comb6_i0_i52 (.D(comb6_71__N_1993[52]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i52.GSR = "ENABLED";
    FD1P3AX comb6_i0_i51 (.D(comb6_71__N_1993[51]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i51.GSR = "ENABLED";
    FD1P3AX comb6_i0_i50 (.D(comb6_71__N_1993[50]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i50.GSR = "ENABLED";
    FD1P3AX comb6_i0_i49 (.D(comb6_71__N_1993[49]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i49.GSR = "ENABLED";
    FD1P3AX comb6_i0_i48 (.D(comb6_71__N_1993[48]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i48.GSR = "ENABLED";
    FD1P3AX comb6_i0_i47 (.D(comb6_71__N_1993[47]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i47.GSR = "ENABLED";
    FD1P3AX comb6_i0_i46 (.D(comb6_71__N_1993[46]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i46.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_206 (.A(count[6]), .B(count[3]), .C(count[10]), 
         .D(count[0]), .Z(n18792)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_206.init = 16'hfffe;
    FD1P3AX comb6_i0_i45 (.D(comb6_71__N_1993[45]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i45.GSR = "ENABLED";
    FD1P3AX comb6_i0_i44 (.D(comb6_71__N_1993[44]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i44.GSR = "ENABLED";
    FD1P3AX comb6_i0_i43 (.D(comb6_71__N_1993[43]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i43.GSR = "ENABLED";
    FD1P3AX comb6_i0_i42 (.D(comb6_71__N_1993[42]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i42.GSR = "ENABLED";
    FD1P3AX comb6_i0_i41 (.D(comb6_71__N_1993[41]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i41.GSR = "ENABLED";
    FD1P3AX comb6_i0_i40 (.D(comb6_71__N_1993[40]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i40.GSR = "ENABLED";
    FD1P3AX comb6_i0_i39 (.D(comb6_71__N_1993[39]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i39.GSR = "ENABLED";
    FD1P3AX comb6_i0_i38 (.D(comb6_71__N_1993[38]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i38.GSR = "ENABLED";
    FD1P3AX comb6_i0_i37 (.D(comb6_71__N_1993[37]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i37.GSR = "ENABLED";
    FD1P3AX comb6_i0_i36 (.D(comb6_71__N_1993[36]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i36.GSR = "ENABLED";
    FD1P3AX comb6_i0_i35 (.D(comb6_71__N_1993[35]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i35.GSR = "ENABLED";
    FD1P3AX comb6_i0_i34 (.D(comb6_71__N_1993[34]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i34.GSR = "ENABLED";
    FD1P3AX comb6_i0_i33 (.D(comb6_71__N_1993[33]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i33.GSR = "ENABLED";
    FD1P3AX comb6_i0_i32 (.D(comb6_71__N_1993[32]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i32.GSR = "ENABLED";
    FD1P3AX comb6_i0_i31 (.D(comb6_71__N_1993[31]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i31.GSR = "ENABLED";
    FD1P3AX comb6_i0_i30 (.D(comb6_71__N_1993[30]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i30.GSR = "ENABLED";
    FD1P3AX comb6_i0_i29 (.D(comb6_71__N_1993[29]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i29.GSR = "ENABLED";
    FD1P3AX comb6_i0_i28 (.D(comb6_71__N_1993[28]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i28.GSR = "ENABLED";
    FD1P3AX comb6_i0_i27 (.D(comb6_71__N_1993[27]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i27.GSR = "ENABLED";
    FD1P3AX comb6_i0_i26 (.D(comb6_71__N_1993[26]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i26.GSR = "ENABLED";
    FD1P3AX comb6_i0_i25 (.D(comb6_71__N_1993[25]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i25.GSR = "ENABLED";
    FD1P3AX comb6_i0_i24 (.D(comb6_71__N_1993[24]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i24.GSR = "ENABLED";
    FD1P3AX comb6_i0_i23 (.D(comb6_71__N_1993[23]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i23.GSR = "ENABLED";
    FD1P3AX comb6_i0_i22 (.D(comb6_71__N_1993[22]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i22.GSR = "ENABLED";
    FD1P3AX comb6_i0_i21 (.D(comb6_71__N_1993[21]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i21.GSR = "ENABLED";
    FD1P3AX comb6_i0_i20 (.D(comb6_71__N_1993[20]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i20.GSR = "ENABLED";
    FD1P3AX comb6_i0_i19 (.D(comb6_71__N_1993[19]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i19.GSR = "ENABLED";
    FD1P3AX comb6_i0_i18 (.D(comb6_71__N_1993[18]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i18.GSR = "ENABLED";
    FD1P3AX comb6_i0_i17 (.D(comb6_71__N_1993[17]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i17.GSR = "ENABLED";
    FD1P3AX comb6_i0_i16 (.D(comb6_71__N_1993[16]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i16.GSR = "ENABLED";
    FD1P3AX comb6_i0_i15 (.D(comb6_71__N_1993[15]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i15.GSR = "ENABLED";
    FD1P3AX comb6_i0_i14 (.D(comb6_71__N_1993[14]), .SP(clk_80mhz_enable_1423), 
            .CK(clk_80mhz), .Q(comb6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i14.GSR = "ENABLED";
    FD1P3AX comb6_i0_i13 (.D(comb6_71__N_1993[13]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i13.GSR = "ENABLED";
    FD1P3AX comb6_i0_i12 (.D(comb6_71__N_1993[12]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i12.GSR = "ENABLED";
    FD1P3AX comb6_i0_i11 (.D(comb6_71__N_1993[11]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i11.GSR = "ENABLED";
    FD1P3AX comb6_i0_i10 (.D(comb6_71__N_1993[10]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i10.GSR = "ENABLED";
    FD1P3AX comb6_i0_i9 (.D(comb6_71__N_1993[9]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i9.GSR = "ENABLED";
    FD1P3AX comb6_i0_i8 (.D(comb6_71__N_1993[8]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i8.GSR = "ENABLED";
    FD1P3AX comb6_i0_i7 (.D(comb6_71__N_1993[7]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i7.GSR = "ENABLED";
    FD1P3AX comb6_i0_i6 (.D(comb6_71__N_1993[6]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i6.GSR = "ENABLED";
    FD1P3AX comb6_i0_i5 (.D(comb6_71__N_1993[5]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i5.GSR = "ENABLED";
    LUT4 mux_3408_i8_3_lut (.A(n100), .B(n102), .C(cout), .Z(comb10_71__N_2281[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i8_3_lut.init = 16'hcaca;
    FD1P3AX comb6_i0_i4 (.D(comb6_71__N_1993[4]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i4.GSR = "ENABLED";
    FD1P3AX comb6_i0_i3 (.D(comb6_71__N_1993[3]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i3.GSR = "ENABLED";
    FD1P3AX comb6_i0_i2 (.D(comb6_71__N_1993[2]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i2.GSR = "ENABLED";
    FD1P3AX comb6_i0_i1 (.D(comb6_71__N_1993[1]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i1.GSR = "ENABLED";
    FD1S3AX integrator5_i71 (.D(integrator5_71__N_1248[71]), .CK(clk_80mhz), 
            .Q(integrator5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i71.GSR = "ENABLED";
    FD1S3AX integrator5_i70 (.D(integrator5_71__N_1248[70]), .CK(clk_80mhz), 
            .Q(integrator5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i70.GSR = "ENABLED";
    FD1S3AX integrator5_i69 (.D(integrator5_71__N_1248[69]), .CK(clk_80mhz), 
            .Q(integrator5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i69.GSR = "ENABLED";
    FD1S3AX integrator5_i68 (.D(integrator5_71__N_1248[68]), .CK(clk_80mhz), 
            .Q(integrator5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i68.GSR = "ENABLED";
    FD1S3AX integrator5_i67 (.D(integrator5_71__N_1248[67]), .CK(clk_80mhz), 
            .Q(integrator5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i67.GSR = "ENABLED";
    FD1S3AX integrator5_i66 (.D(integrator5_71__N_1248[66]), .CK(clk_80mhz), 
            .Q(integrator5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i66.GSR = "ENABLED";
    FD1S3AX integrator5_i65 (.D(integrator5_71__N_1248[65]), .CK(clk_80mhz), 
            .Q(integrator5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i65.GSR = "ENABLED";
    FD1S3AX integrator5_i64 (.D(integrator5_71__N_1248[64]), .CK(clk_80mhz), 
            .Q(integrator5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i64.GSR = "ENABLED";
    FD1S3AX integrator5_i63 (.D(integrator5_71__N_1248[63]), .CK(clk_80mhz), 
            .Q(integrator5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i63.GSR = "ENABLED";
    FD1S3AX integrator5_i62 (.D(integrator5_71__N_1248[62]), .CK(clk_80mhz), 
            .Q(integrator5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i62.GSR = "ENABLED";
    FD1S3AX integrator5_i61 (.D(integrator5_71__N_1248[61]), .CK(clk_80mhz), 
            .Q(integrator5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i61.GSR = "ENABLED";
    FD1S3AX integrator5_i60 (.D(integrator5_71__N_1248[60]), .CK(clk_80mhz), 
            .Q(integrator5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i60.GSR = "ENABLED";
    FD1S3AX integrator5_i59 (.D(integrator5_71__N_1248[59]), .CK(clk_80mhz), 
            .Q(integrator5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i59.GSR = "ENABLED";
    FD1S3AX integrator5_i58 (.D(integrator5_71__N_1248[58]), .CK(clk_80mhz), 
            .Q(integrator5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i58.GSR = "ENABLED";
    FD1S3AX integrator5_i57 (.D(integrator5_71__N_1248[57]), .CK(clk_80mhz), 
            .Q(integrator5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i57.GSR = "ENABLED";
    FD1S3AX integrator5_i56 (.D(integrator5_71__N_1248[56]), .CK(clk_80mhz), 
            .Q(integrator5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i56.GSR = "ENABLED";
    FD1S3AX integrator5_i55 (.D(integrator5_71__N_1248[55]), .CK(clk_80mhz), 
            .Q(integrator5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i55.GSR = "ENABLED";
    FD1S3AX integrator5_i54 (.D(integrator5_71__N_1248[54]), .CK(clk_80mhz), 
            .Q(integrator5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i54.GSR = "ENABLED";
    FD1S3AX integrator5_i53 (.D(integrator5_71__N_1248[53]), .CK(clk_80mhz), 
            .Q(integrator5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i53.GSR = "ENABLED";
    FD1S3AX integrator5_i52 (.D(integrator5_71__N_1248[52]), .CK(clk_80mhz), 
            .Q(integrator5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i52.GSR = "ENABLED";
    FD1S3AX integrator5_i51 (.D(integrator5_71__N_1248[51]), .CK(clk_80mhz), 
            .Q(integrator5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i51.GSR = "ENABLED";
    FD1S3AX integrator5_i50 (.D(integrator5_71__N_1248[50]), .CK(clk_80mhz), 
            .Q(integrator5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i50.GSR = "ENABLED";
    FD1S3AX integrator5_i49 (.D(integrator5_71__N_1248[49]), .CK(clk_80mhz), 
            .Q(integrator5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i49.GSR = "ENABLED";
    FD1S3AX integrator5_i48 (.D(integrator5_71__N_1248[48]), .CK(clk_80mhz), 
            .Q(integrator5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i48.GSR = "ENABLED";
    FD1S3AX integrator5_i47 (.D(integrator5_71__N_1248[47]), .CK(clk_80mhz), 
            .Q(integrator5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i47.GSR = "ENABLED";
    FD1S3AX integrator5_i46 (.D(integrator5_71__N_1248[46]), .CK(clk_80mhz), 
            .Q(integrator5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i46.GSR = "ENABLED";
    FD1S3AX integrator5_i45 (.D(integrator5_71__N_1248[45]), .CK(clk_80mhz), 
            .Q(integrator5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i45.GSR = "ENABLED";
    FD1S3AX integrator5_i44 (.D(integrator5_71__N_1248[44]), .CK(clk_80mhz), 
            .Q(integrator5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i44.GSR = "ENABLED";
    FD1S3AX integrator5_i43 (.D(integrator5_71__N_1248[43]), .CK(clk_80mhz), 
            .Q(integrator5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i43.GSR = "ENABLED";
    FD1S3AX integrator5_i42 (.D(integrator5_71__N_1248[42]), .CK(clk_80mhz), 
            .Q(integrator5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i42.GSR = "ENABLED";
    FD1S3AX integrator5_i41 (.D(integrator5_71__N_1248[41]), .CK(clk_80mhz), 
            .Q(integrator5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i41.GSR = "ENABLED";
    FD1S3AX integrator5_i40 (.D(integrator5_71__N_1248[40]), .CK(clk_80mhz), 
            .Q(integrator5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i40.GSR = "ENABLED";
    FD1S3AX integrator5_i39 (.D(integrator5_71__N_1248[39]), .CK(clk_80mhz), 
            .Q(integrator5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i39.GSR = "ENABLED";
    FD1S3AX integrator5_i38 (.D(integrator5_71__N_1248[38]), .CK(clk_80mhz), 
            .Q(integrator5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i38.GSR = "ENABLED";
    FD1S3AX integrator5_i37 (.D(integrator5_71__N_1248[37]), .CK(clk_80mhz), 
            .Q(integrator5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i37.GSR = "ENABLED";
    FD1S3AX integrator5_i36 (.D(integrator5_71__N_1248[36]), .CK(clk_80mhz), 
            .Q(integrator5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i36.GSR = "ENABLED";
    FD1S3AX integrator5_i35 (.D(integrator5_71__N_1248[35]), .CK(clk_80mhz), 
            .Q(integrator5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i35.GSR = "ENABLED";
    FD1S3AX integrator5_i34 (.D(integrator5_71__N_1248[34]), .CK(clk_80mhz), 
            .Q(integrator5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i34.GSR = "ENABLED";
    FD1S3AX integrator5_i33 (.D(integrator5_71__N_1248[33]), .CK(clk_80mhz), 
            .Q(integrator5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i33.GSR = "ENABLED";
    FD1S3AX integrator5_i32 (.D(integrator5_71__N_1248[32]), .CK(clk_80mhz), 
            .Q(integrator5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i32.GSR = "ENABLED";
    FD1S3AX integrator5_i31 (.D(integrator5_71__N_1248[31]), .CK(clk_80mhz), 
            .Q(integrator5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i31.GSR = "ENABLED";
    FD1S3AX integrator5_i30 (.D(integrator5_71__N_1248[30]), .CK(clk_80mhz), 
            .Q(integrator5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i30.GSR = "ENABLED";
    FD1S3AX integrator5_i29 (.D(integrator5_71__N_1248[29]), .CK(clk_80mhz), 
            .Q(integrator5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i29.GSR = "ENABLED";
    FD1S3AX integrator5_i28 (.D(integrator5_71__N_1248[28]), .CK(clk_80mhz), 
            .Q(integrator5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i28.GSR = "ENABLED";
    FD1S3AX integrator5_i27 (.D(integrator5_71__N_1248[27]), .CK(clk_80mhz), 
            .Q(integrator5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i27.GSR = "ENABLED";
    FD1S3AX integrator5_i26 (.D(integrator5_71__N_1248[26]), .CK(clk_80mhz), 
            .Q(integrator5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i26.GSR = "ENABLED";
    FD1S3AX integrator5_i25 (.D(integrator5_71__N_1248[25]), .CK(clk_80mhz), 
            .Q(integrator5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i25.GSR = "ENABLED";
    FD1S3AX integrator5_i24 (.D(integrator5_71__N_1248[24]), .CK(clk_80mhz), 
            .Q(integrator5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i24.GSR = "ENABLED";
    FD1S3AX integrator5_i23 (.D(integrator5_71__N_1248[23]), .CK(clk_80mhz), 
            .Q(integrator5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i23.GSR = "ENABLED";
    FD1S3AX integrator5_i22 (.D(integrator5_71__N_1248[22]), .CK(clk_80mhz), 
            .Q(integrator5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i22.GSR = "ENABLED";
    FD1S3AX integrator5_i21 (.D(integrator5_71__N_1248[21]), .CK(clk_80mhz), 
            .Q(integrator5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i21.GSR = "ENABLED";
    FD1S3AX integrator5_i20 (.D(integrator5_71__N_1248[20]), .CK(clk_80mhz), 
            .Q(integrator5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i20.GSR = "ENABLED";
    FD1S3AX integrator5_i19 (.D(integrator5_71__N_1248[19]), .CK(clk_80mhz), 
            .Q(integrator5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i19.GSR = "ENABLED";
    FD1S3AX integrator5_i18 (.D(integrator5_71__N_1248[18]), .CK(clk_80mhz), 
            .Q(integrator5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i18.GSR = "ENABLED";
    FD1S3AX integrator5_i17 (.D(integrator5_71__N_1248[17]), .CK(clk_80mhz), 
            .Q(integrator5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i17.GSR = "ENABLED";
    FD1S3AX integrator5_i16 (.D(integrator5_71__N_1248[16]), .CK(clk_80mhz), 
            .Q(integrator5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i16.GSR = "ENABLED";
    FD1S3AX integrator5_i15 (.D(integrator5_71__N_1248[15]), .CK(clk_80mhz), 
            .Q(integrator5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i15.GSR = "ENABLED";
    FD1S3AX integrator5_i14 (.D(integrator5_71__N_1248[14]), .CK(clk_80mhz), 
            .Q(integrator5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i14.GSR = "ENABLED";
    FD1S3AX integrator5_i13 (.D(integrator5_71__N_1248[13]), .CK(clk_80mhz), 
            .Q(integrator5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i13.GSR = "ENABLED";
    FD1S3AX integrator5_i12 (.D(integrator5_71__N_1248[12]), .CK(clk_80mhz), 
            .Q(integrator5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i12.GSR = "ENABLED";
    FD1S3AX integrator5_i11 (.D(integrator5_71__N_1248[11]), .CK(clk_80mhz), 
            .Q(integrator5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i11.GSR = "ENABLED";
    FD1S3AX integrator5_i10 (.D(integrator5_71__N_1248[10]), .CK(clk_80mhz), 
            .Q(integrator5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i10.GSR = "ENABLED";
    FD1S3AX integrator5_i9 (.D(integrator5_71__N_1248[9]), .CK(clk_80mhz), 
            .Q(integrator5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i9.GSR = "ENABLED";
    FD1S3AX integrator5_i8 (.D(integrator5_71__N_1248[8]), .CK(clk_80mhz), 
            .Q(integrator5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i8.GSR = "ENABLED";
    FD1S3AX integrator5_i7 (.D(integrator5_71__N_1248[7]), .CK(clk_80mhz), 
            .Q(integrator5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i7.GSR = "ENABLED";
    FD1S3AX integrator5_i6 (.D(integrator5_71__N_1248[6]), .CK(clk_80mhz), 
            .Q(integrator5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i6.GSR = "ENABLED";
    FD1S3AX integrator5_i5 (.D(integrator5_71__N_1248[5]), .CK(clk_80mhz), 
            .Q(integrator5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i5.GSR = "ENABLED";
    FD1S3AX integrator5_i4 (.D(integrator5_71__N_1248[4]), .CK(clk_80mhz), 
            .Q(integrator5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i4.GSR = "ENABLED";
    FD1S3AX integrator5_i3 (.D(integrator5_71__N_1248[3]), .CK(clk_80mhz), 
            .Q(integrator5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i3.GSR = "ENABLED";
    FD1S3AX integrator5_i2 (.D(integrator5_71__N_1248[2]), .CK(clk_80mhz), 
            .Q(integrator5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i2.GSR = "ENABLED";
    FD1S3AX integrator5_i1 (.D(integrator5_71__N_1248[1]), .CK(clk_80mhz), 
            .Q(integrator5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i1.GSR = "ENABLED";
    FD1S3AX integrator4_i71 (.D(integrator4_71__N_1176[71]), .CK(clk_80mhz), 
            .Q(integrator4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i71.GSR = "ENABLED";
    FD1S3AX integrator4_i70 (.D(integrator4_71__N_1176[70]), .CK(clk_80mhz), 
            .Q(integrator4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i70.GSR = "ENABLED";
    FD1S3AX integrator4_i69 (.D(integrator4_71__N_1176[69]), .CK(clk_80mhz), 
            .Q(integrator4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i69.GSR = "ENABLED";
    FD1S3AX integrator4_i68 (.D(integrator4_71__N_1176[68]), .CK(clk_80mhz), 
            .Q(integrator4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i68.GSR = "ENABLED";
    FD1S3AX integrator4_i67 (.D(integrator4_71__N_1176[67]), .CK(clk_80mhz), 
            .Q(integrator4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i67.GSR = "ENABLED";
    FD1S3AX integrator4_i66 (.D(integrator4_71__N_1176[66]), .CK(clk_80mhz), 
            .Q(integrator4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i66.GSR = "ENABLED";
    FD1S3AX integrator4_i65 (.D(integrator4_71__N_1176[65]), .CK(clk_80mhz), 
            .Q(integrator4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i65.GSR = "ENABLED";
    FD1S3AX integrator4_i64 (.D(integrator4_71__N_1176[64]), .CK(clk_80mhz), 
            .Q(integrator4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i64.GSR = "ENABLED";
    FD1S3AX integrator4_i63 (.D(integrator4_71__N_1176[63]), .CK(clk_80mhz), 
            .Q(integrator4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i63.GSR = "ENABLED";
    FD1S3AX integrator4_i62 (.D(integrator4_71__N_1176[62]), .CK(clk_80mhz), 
            .Q(integrator4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i62.GSR = "ENABLED";
    FD1S3AX integrator4_i61 (.D(integrator4_71__N_1176[61]), .CK(clk_80mhz), 
            .Q(integrator4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i61.GSR = "ENABLED";
    FD1S3AX integrator4_i60 (.D(integrator4_71__N_1176[60]), .CK(clk_80mhz), 
            .Q(integrator4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i60.GSR = "ENABLED";
    FD1S3AX integrator4_i59 (.D(integrator4_71__N_1176[59]), .CK(clk_80mhz), 
            .Q(integrator4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i59.GSR = "ENABLED";
    FD1S3AX integrator4_i58 (.D(integrator4_71__N_1176[58]), .CK(clk_80mhz), 
            .Q(integrator4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i58.GSR = "ENABLED";
    FD1S3AX integrator4_i57 (.D(integrator4_71__N_1176[57]), .CK(clk_80mhz), 
            .Q(integrator4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i57.GSR = "ENABLED";
    FD1S3AX integrator4_i56 (.D(integrator4_71__N_1176[56]), .CK(clk_80mhz), 
            .Q(integrator4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i56.GSR = "ENABLED";
    FD1S3AX integrator4_i55 (.D(integrator4_71__N_1176[55]), .CK(clk_80mhz), 
            .Q(integrator4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i55.GSR = "ENABLED";
    FD1S3AX integrator4_i54 (.D(integrator4_71__N_1176[54]), .CK(clk_80mhz), 
            .Q(integrator4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i54.GSR = "ENABLED";
    FD1S3AX integrator4_i53 (.D(integrator4_71__N_1176[53]), .CK(clk_80mhz), 
            .Q(integrator4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i53.GSR = "ENABLED";
    FD1S3AX integrator4_i52 (.D(integrator4_71__N_1176[52]), .CK(clk_80mhz), 
            .Q(integrator4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i52.GSR = "ENABLED";
    FD1S3AX integrator4_i51 (.D(integrator4_71__N_1176[51]), .CK(clk_80mhz), 
            .Q(integrator4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i51.GSR = "ENABLED";
    FD1S3AX integrator4_i50 (.D(integrator4_71__N_1176[50]), .CK(clk_80mhz), 
            .Q(integrator4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i50.GSR = "ENABLED";
    FD1S3AX integrator4_i49 (.D(integrator4_71__N_1176[49]), .CK(clk_80mhz), 
            .Q(integrator4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i49.GSR = "ENABLED";
    FD1S3AX integrator4_i48 (.D(integrator4_71__N_1176[48]), .CK(clk_80mhz), 
            .Q(integrator4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i48.GSR = "ENABLED";
    FD1S3AX integrator4_i47 (.D(integrator4_71__N_1176[47]), .CK(clk_80mhz), 
            .Q(integrator4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i47.GSR = "ENABLED";
    FD1S3AX integrator4_i46 (.D(integrator4_71__N_1176[46]), .CK(clk_80mhz), 
            .Q(integrator4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i46.GSR = "ENABLED";
    FD1S3AX integrator4_i45 (.D(integrator4_71__N_1176[45]), .CK(clk_80mhz), 
            .Q(integrator4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i45.GSR = "ENABLED";
    FD1S3AX integrator4_i44 (.D(integrator4_71__N_1176[44]), .CK(clk_80mhz), 
            .Q(integrator4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i44.GSR = "ENABLED";
    FD1S3AX integrator4_i43 (.D(integrator4_71__N_1176[43]), .CK(clk_80mhz), 
            .Q(integrator4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i43.GSR = "ENABLED";
    FD1S3AX integrator4_i42 (.D(integrator4_71__N_1176[42]), .CK(clk_80mhz), 
            .Q(integrator4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i42.GSR = "ENABLED";
    FD1S3AX integrator4_i41 (.D(integrator4_71__N_1176[41]), .CK(clk_80mhz), 
            .Q(integrator4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i41.GSR = "ENABLED";
    FD1S3AX integrator4_i40 (.D(integrator4_71__N_1176[40]), .CK(clk_80mhz), 
            .Q(integrator4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i40.GSR = "ENABLED";
    FD1S3AX integrator4_i39 (.D(integrator4_71__N_1176[39]), .CK(clk_80mhz), 
            .Q(integrator4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i39.GSR = "ENABLED";
    FD1S3AX integrator4_i38 (.D(integrator4_71__N_1176[38]), .CK(clk_80mhz), 
            .Q(integrator4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i38.GSR = "ENABLED";
    FD1S3AX integrator4_i37 (.D(integrator4_71__N_1176[37]), .CK(clk_80mhz), 
            .Q(integrator4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i37.GSR = "ENABLED";
    FD1S3AX integrator4_i36 (.D(integrator4_71__N_1176[36]), .CK(clk_80mhz), 
            .Q(integrator4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i36.GSR = "ENABLED";
    FD1S3AX integrator4_i35 (.D(integrator4_71__N_1176[35]), .CK(clk_80mhz), 
            .Q(integrator4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i35.GSR = "ENABLED";
    FD1S3AX integrator4_i34 (.D(integrator4_71__N_1176[34]), .CK(clk_80mhz), 
            .Q(integrator4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i34.GSR = "ENABLED";
    FD1S3AX integrator4_i33 (.D(integrator4_71__N_1176[33]), .CK(clk_80mhz), 
            .Q(integrator4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i33.GSR = "ENABLED";
    FD1S3AX integrator4_i32 (.D(integrator4_71__N_1176[32]), .CK(clk_80mhz), 
            .Q(integrator4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i32.GSR = "ENABLED";
    FD1S3AX integrator4_i31 (.D(integrator4_71__N_1176[31]), .CK(clk_80mhz), 
            .Q(integrator4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i31.GSR = "ENABLED";
    FD1S3AX integrator4_i30 (.D(integrator4_71__N_1176[30]), .CK(clk_80mhz), 
            .Q(integrator4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i30.GSR = "ENABLED";
    FD1S3AX integrator4_i29 (.D(integrator4_71__N_1176[29]), .CK(clk_80mhz), 
            .Q(integrator4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i29.GSR = "ENABLED";
    FD1S3AX integrator4_i28 (.D(integrator4_71__N_1176[28]), .CK(clk_80mhz), 
            .Q(integrator4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i28.GSR = "ENABLED";
    FD1S3AX integrator4_i27 (.D(integrator4_71__N_1176[27]), .CK(clk_80mhz), 
            .Q(integrator4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i27.GSR = "ENABLED";
    FD1S3AX integrator4_i26 (.D(integrator4_71__N_1176[26]), .CK(clk_80mhz), 
            .Q(integrator4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i26.GSR = "ENABLED";
    FD1S3AX integrator4_i25 (.D(integrator4_71__N_1176[25]), .CK(clk_80mhz), 
            .Q(integrator4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i25.GSR = "ENABLED";
    FD1S3AX integrator4_i24 (.D(integrator4_71__N_1176[24]), .CK(clk_80mhz), 
            .Q(integrator4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i24.GSR = "ENABLED";
    FD1S3AX integrator4_i23 (.D(integrator4_71__N_1176[23]), .CK(clk_80mhz), 
            .Q(integrator4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i23.GSR = "ENABLED";
    FD1S3AX integrator4_i22 (.D(integrator4_71__N_1176[22]), .CK(clk_80mhz), 
            .Q(integrator4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i22.GSR = "ENABLED";
    FD1S3AX integrator4_i21 (.D(integrator4_71__N_1176[21]), .CK(clk_80mhz), 
            .Q(integrator4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i21.GSR = "ENABLED";
    FD1S3AX integrator4_i20 (.D(integrator4_71__N_1176[20]), .CK(clk_80mhz), 
            .Q(integrator4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i20.GSR = "ENABLED";
    FD1S3AX integrator4_i19 (.D(integrator4_71__N_1176[19]), .CK(clk_80mhz), 
            .Q(integrator4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i19.GSR = "ENABLED";
    FD1S3AX integrator4_i18 (.D(integrator4_71__N_1176[18]), .CK(clk_80mhz), 
            .Q(integrator4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i18.GSR = "ENABLED";
    FD1S3AX integrator4_i17 (.D(integrator4_71__N_1176[17]), .CK(clk_80mhz), 
            .Q(integrator4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i17.GSR = "ENABLED";
    FD1S3AX integrator4_i16 (.D(integrator4_71__N_1176[16]), .CK(clk_80mhz), 
            .Q(integrator4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i16.GSR = "ENABLED";
    FD1S3AX integrator4_i15 (.D(integrator4_71__N_1176[15]), .CK(clk_80mhz), 
            .Q(integrator4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i15.GSR = "ENABLED";
    FD1S3AX integrator4_i14 (.D(integrator4_71__N_1176[14]), .CK(clk_80mhz), 
            .Q(integrator4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i14.GSR = "ENABLED";
    FD1S3AX integrator4_i13 (.D(integrator4_71__N_1176[13]), .CK(clk_80mhz), 
            .Q(integrator4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i13.GSR = "ENABLED";
    FD1S3AX integrator4_i12 (.D(integrator4_71__N_1176[12]), .CK(clk_80mhz), 
            .Q(integrator4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i12.GSR = "ENABLED";
    FD1S3AX integrator4_i11 (.D(integrator4_71__N_1176[11]), .CK(clk_80mhz), 
            .Q(integrator4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i11.GSR = "ENABLED";
    FD1S3AX integrator4_i10 (.D(integrator4_71__N_1176[10]), .CK(clk_80mhz), 
            .Q(integrator4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i10.GSR = "ENABLED";
    FD1S3AX integrator4_i9 (.D(integrator4_71__N_1176[9]), .CK(clk_80mhz), 
            .Q(integrator4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i9.GSR = "ENABLED";
    FD1S3AX integrator4_i8 (.D(integrator4_71__N_1176[8]), .CK(clk_80mhz), 
            .Q(integrator4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i8.GSR = "ENABLED";
    FD1S3AX integrator4_i7 (.D(integrator4_71__N_1176[7]), .CK(clk_80mhz), 
            .Q(integrator4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i7.GSR = "ENABLED";
    FD1S3AX integrator4_i6 (.D(integrator4_71__N_1176[6]), .CK(clk_80mhz), 
            .Q(integrator4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i6.GSR = "ENABLED";
    FD1S3AX integrator4_i5 (.D(integrator4_71__N_1176[5]), .CK(clk_80mhz), 
            .Q(integrator4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i5.GSR = "ENABLED";
    FD1S3AX integrator4_i4 (.D(integrator4_71__N_1176[4]), .CK(clk_80mhz), 
            .Q(integrator4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i4.GSR = "ENABLED";
    FD1S3AX integrator4_i3 (.D(integrator4_71__N_1176[3]), .CK(clk_80mhz), 
            .Q(integrator4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i3.GSR = "ENABLED";
    FD1S3AX integrator4_i2 (.D(integrator4_71__N_1176[2]), .CK(clk_80mhz), 
            .Q(integrator4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i2.GSR = "ENABLED";
    FD1S3AX integrator4_i1 (.D(integrator4_71__N_1176[1]), .CK(clk_80mhz), 
            .Q(integrator4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i1.GSR = "ENABLED";
    FD1S3AX integrator3_i71 (.D(integrator3_71__N_1104[71]), .CK(clk_80mhz), 
            .Q(integrator3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i71.GSR = "ENABLED";
    FD1S3AX integrator3_i70 (.D(integrator3_71__N_1104[70]), .CK(clk_80mhz), 
            .Q(integrator3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i70.GSR = "ENABLED";
    FD1S3AX integrator3_i69 (.D(integrator3_71__N_1104[69]), .CK(clk_80mhz), 
            .Q(integrator3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i69.GSR = "ENABLED";
    FD1S3AX integrator3_i68 (.D(integrator3_71__N_1104[68]), .CK(clk_80mhz), 
            .Q(integrator3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i68.GSR = "ENABLED";
    FD1S3AX integrator3_i67 (.D(integrator3_71__N_1104[67]), .CK(clk_80mhz), 
            .Q(integrator3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i67.GSR = "ENABLED";
    FD1S3AX integrator3_i66 (.D(integrator3_71__N_1104[66]), .CK(clk_80mhz), 
            .Q(integrator3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i66.GSR = "ENABLED";
    FD1S3AX integrator3_i65 (.D(integrator3_71__N_1104[65]), .CK(clk_80mhz), 
            .Q(integrator3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i65.GSR = "ENABLED";
    FD1S3AX integrator3_i64 (.D(integrator3_71__N_1104[64]), .CK(clk_80mhz), 
            .Q(integrator3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i64.GSR = "ENABLED";
    FD1S3AX integrator3_i63 (.D(integrator3_71__N_1104[63]), .CK(clk_80mhz), 
            .Q(integrator3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i63.GSR = "ENABLED";
    FD1S3AX integrator3_i62 (.D(integrator3_71__N_1104[62]), .CK(clk_80mhz), 
            .Q(integrator3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i62.GSR = "ENABLED";
    FD1S3AX integrator3_i61 (.D(integrator3_71__N_1104[61]), .CK(clk_80mhz), 
            .Q(integrator3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i61.GSR = "ENABLED";
    FD1S3AX integrator3_i60 (.D(integrator3_71__N_1104[60]), .CK(clk_80mhz), 
            .Q(integrator3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i60.GSR = "ENABLED";
    FD1S3AX integrator3_i59 (.D(integrator3_71__N_1104[59]), .CK(clk_80mhz), 
            .Q(integrator3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i59.GSR = "ENABLED";
    FD1S3AX integrator3_i58 (.D(integrator3_71__N_1104[58]), .CK(clk_80mhz), 
            .Q(integrator3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i58.GSR = "ENABLED";
    FD1S3AX integrator3_i57 (.D(integrator3_71__N_1104[57]), .CK(clk_80mhz), 
            .Q(integrator3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i57.GSR = "ENABLED";
    FD1S3AX integrator3_i56 (.D(integrator3_71__N_1104[56]), .CK(clk_80mhz), 
            .Q(integrator3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i56.GSR = "ENABLED";
    FD1S3AX integrator3_i55 (.D(integrator3_71__N_1104[55]), .CK(clk_80mhz), 
            .Q(integrator3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i55.GSR = "ENABLED";
    FD1S3AX integrator3_i54 (.D(integrator3_71__N_1104[54]), .CK(clk_80mhz), 
            .Q(integrator3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i54.GSR = "ENABLED";
    FD1S3AX integrator3_i53 (.D(integrator3_71__N_1104[53]), .CK(clk_80mhz), 
            .Q(integrator3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i53.GSR = "ENABLED";
    FD1S3AX integrator3_i52 (.D(integrator3_71__N_1104[52]), .CK(clk_80mhz), 
            .Q(integrator3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i52.GSR = "ENABLED";
    FD1S3AX integrator3_i51 (.D(integrator3_71__N_1104[51]), .CK(clk_80mhz), 
            .Q(integrator3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i51.GSR = "ENABLED";
    FD1S3AX integrator3_i50 (.D(integrator3_71__N_1104[50]), .CK(clk_80mhz), 
            .Q(integrator3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i50.GSR = "ENABLED";
    FD1S3AX integrator3_i49 (.D(integrator3_71__N_1104[49]), .CK(clk_80mhz), 
            .Q(integrator3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i49.GSR = "ENABLED";
    FD1S3AX integrator3_i48 (.D(integrator3_71__N_1104[48]), .CK(clk_80mhz), 
            .Q(integrator3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i48.GSR = "ENABLED";
    FD1S3AX integrator3_i47 (.D(integrator3_71__N_1104[47]), .CK(clk_80mhz), 
            .Q(integrator3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i47.GSR = "ENABLED";
    FD1S3AX integrator3_i46 (.D(integrator3_71__N_1104[46]), .CK(clk_80mhz), 
            .Q(integrator3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i46.GSR = "ENABLED";
    FD1S3AX integrator3_i45 (.D(integrator3_71__N_1104[45]), .CK(clk_80mhz), 
            .Q(integrator3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i45.GSR = "ENABLED";
    FD1S3AX integrator3_i44 (.D(integrator3_71__N_1104[44]), .CK(clk_80mhz), 
            .Q(integrator3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i44.GSR = "ENABLED";
    FD1S3AX integrator3_i43 (.D(integrator3_71__N_1104[43]), .CK(clk_80mhz), 
            .Q(integrator3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i43.GSR = "ENABLED";
    LUT4 mux_3408_i7_3_lut (.A(n103), .B(n105), .C(cout), .Z(comb10_71__N_2281[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i7_3_lut.init = 16'hcaca;
    FD1S3AX integrator3_i42 (.D(integrator3_71__N_1104[42]), .CK(clk_80mhz), 
            .Q(integrator3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i42.GSR = "ENABLED";
    FD1S3AX integrator3_i41 (.D(integrator3_71__N_1104[41]), .CK(clk_80mhz), 
            .Q(integrator3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i41.GSR = "ENABLED";
    FD1S3AX integrator3_i40 (.D(integrator3_71__N_1104[40]), .CK(clk_80mhz), 
            .Q(integrator3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i40.GSR = "ENABLED";
    FD1S3AX integrator3_i39 (.D(integrator3_71__N_1104[39]), .CK(clk_80mhz), 
            .Q(integrator3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i39.GSR = "ENABLED";
    FD1S3AX integrator3_i38 (.D(integrator3_71__N_1104[38]), .CK(clk_80mhz), 
            .Q(integrator3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i38.GSR = "ENABLED";
    FD1S3AX integrator3_i37 (.D(integrator3_71__N_1104[37]), .CK(clk_80mhz), 
            .Q(integrator3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i37.GSR = "ENABLED";
    FD1S3AX integrator3_i36 (.D(integrator3_71__N_1104[36]), .CK(clk_80mhz), 
            .Q(integrator3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i36.GSR = "ENABLED";
    FD1S3AX integrator3_i35 (.D(integrator3_71__N_1104[35]), .CK(clk_80mhz), 
            .Q(integrator3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i35.GSR = "ENABLED";
    FD1S3AX integrator3_i34 (.D(integrator3_71__N_1104[34]), .CK(clk_80mhz), 
            .Q(integrator3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i34.GSR = "ENABLED";
    FD1S3AX integrator3_i33 (.D(integrator3_71__N_1104[33]), .CK(clk_80mhz), 
            .Q(integrator3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i33.GSR = "ENABLED";
    FD1S3AX integrator3_i32 (.D(integrator3_71__N_1104[32]), .CK(clk_80mhz), 
            .Q(integrator3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i32.GSR = "ENABLED";
    FD1S3AX integrator3_i31 (.D(integrator3_71__N_1104[31]), .CK(clk_80mhz), 
            .Q(integrator3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i31.GSR = "ENABLED";
    FD1S3AX integrator3_i30 (.D(integrator3_71__N_1104[30]), .CK(clk_80mhz), 
            .Q(integrator3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i30.GSR = "ENABLED";
    FD1S3AX integrator3_i29 (.D(integrator3_71__N_1104[29]), .CK(clk_80mhz), 
            .Q(integrator3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i29.GSR = "ENABLED";
    FD1S3AX integrator3_i28 (.D(integrator3_71__N_1104[28]), .CK(clk_80mhz), 
            .Q(integrator3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i28.GSR = "ENABLED";
    FD1S3AX integrator3_i27 (.D(integrator3_71__N_1104[27]), .CK(clk_80mhz), 
            .Q(integrator3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i27.GSR = "ENABLED";
    FD1S3AX integrator3_i26 (.D(integrator3_71__N_1104[26]), .CK(clk_80mhz), 
            .Q(integrator3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i26.GSR = "ENABLED";
    FD1S3AX integrator3_i25 (.D(integrator3_71__N_1104[25]), .CK(clk_80mhz), 
            .Q(integrator3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i25.GSR = "ENABLED";
    FD1S3AX integrator3_i24 (.D(integrator3_71__N_1104[24]), .CK(clk_80mhz), 
            .Q(integrator3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i24.GSR = "ENABLED";
    FD1S3AX integrator3_i23 (.D(integrator3_71__N_1104[23]), .CK(clk_80mhz), 
            .Q(integrator3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i23.GSR = "ENABLED";
    FD1S3AX integrator3_i22 (.D(integrator3_71__N_1104[22]), .CK(clk_80mhz), 
            .Q(integrator3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i22.GSR = "ENABLED";
    FD1S3AX integrator3_i21 (.D(integrator3_71__N_1104[21]), .CK(clk_80mhz), 
            .Q(integrator3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i21.GSR = "ENABLED";
    FD1S3AX integrator3_i20 (.D(integrator3_71__N_1104[20]), .CK(clk_80mhz), 
            .Q(integrator3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i20.GSR = "ENABLED";
    FD1S3AX integrator3_i19 (.D(integrator3_71__N_1104[19]), .CK(clk_80mhz), 
            .Q(integrator3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i19.GSR = "ENABLED";
    FD1S3AX integrator3_i18 (.D(integrator3_71__N_1104[18]), .CK(clk_80mhz), 
            .Q(integrator3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i18.GSR = "ENABLED";
    FD1S3AX integrator3_i17 (.D(integrator3_71__N_1104[17]), .CK(clk_80mhz), 
            .Q(integrator3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i17.GSR = "ENABLED";
    FD1S3AX integrator3_i16 (.D(integrator3_71__N_1104[16]), .CK(clk_80mhz), 
            .Q(integrator3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i16.GSR = "ENABLED";
    FD1S3AX integrator3_i15 (.D(integrator3_71__N_1104[15]), .CK(clk_80mhz), 
            .Q(integrator3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i15.GSR = "ENABLED";
    FD1S3AX integrator3_i14 (.D(integrator3_71__N_1104[14]), .CK(clk_80mhz), 
            .Q(integrator3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i14.GSR = "ENABLED";
    FD1S3AX integrator3_i13 (.D(integrator3_71__N_1104[13]), .CK(clk_80mhz), 
            .Q(integrator3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i13.GSR = "ENABLED";
    FD1S3AX integrator3_i12 (.D(integrator3_71__N_1104[12]), .CK(clk_80mhz), 
            .Q(integrator3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i12.GSR = "ENABLED";
    FD1S3AX integrator3_i11 (.D(integrator3_71__N_1104[11]), .CK(clk_80mhz), 
            .Q(integrator3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i11.GSR = "ENABLED";
    FD1S3AX integrator3_i10 (.D(integrator3_71__N_1104[10]), .CK(clk_80mhz), 
            .Q(integrator3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i10.GSR = "ENABLED";
    FD1S3AX integrator3_i9 (.D(integrator3_71__N_1104[9]), .CK(clk_80mhz), 
            .Q(integrator3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i9.GSR = "ENABLED";
    FD1S3AX integrator3_i8 (.D(integrator3_71__N_1104[8]), .CK(clk_80mhz), 
            .Q(integrator3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i8.GSR = "ENABLED";
    FD1S3AX integrator3_i7 (.D(integrator3_71__N_1104[7]), .CK(clk_80mhz), 
            .Q(integrator3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i7.GSR = "ENABLED";
    FD1S3AX integrator3_i6 (.D(integrator3_71__N_1104[6]), .CK(clk_80mhz), 
            .Q(integrator3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i6.GSR = "ENABLED";
    FD1S3AX integrator3_i5 (.D(integrator3_71__N_1104[5]), .CK(clk_80mhz), 
            .Q(integrator3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i5.GSR = "ENABLED";
    FD1S3AX integrator3_i4 (.D(integrator3_71__N_1104[4]), .CK(clk_80mhz), 
            .Q(integrator3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i4.GSR = "ENABLED";
    FD1S3AX integrator3_i3 (.D(integrator3_71__N_1104[3]), .CK(clk_80mhz), 
            .Q(integrator3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i3.GSR = "ENABLED";
    FD1S3AX integrator3_i2 (.D(integrator3_71__N_1104[2]), .CK(clk_80mhz), 
            .Q(integrator3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i2.GSR = "ENABLED";
    FD1S3AX integrator3_i1 (.D(integrator3_71__N_1104[1]), .CK(clk_80mhz), 
            .Q(integrator3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i1.GSR = "ENABLED";
    FD1S3AX integrator2_i71 (.D(integrator2_71__N_1032[71]), .CK(clk_80mhz), 
            .Q(integrator2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i71.GSR = "ENABLED";
    FD1S3AX integrator2_i70 (.D(integrator2_71__N_1032[70]), .CK(clk_80mhz), 
            .Q(integrator2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i70.GSR = "ENABLED";
    FD1S3AX integrator2_i69 (.D(integrator2_71__N_1032[69]), .CK(clk_80mhz), 
            .Q(integrator2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i69.GSR = "ENABLED";
    FD1S3AX integrator2_i68 (.D(integrator2_71__N_1032[68]), .CK(clk_80mhz), 
            .Q(integrator2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i68.GSR = "ENABLED";
    FD1S3AX integrator2_i67 (.D(integrator2_71__N_1032[67]), .CK(clk_80mhz), 
            .Q(integrator2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i67.GSR = "ENABLED";
    FD1S3AX integrator2_i66 (.D(integrator2_71__N_1032[66]), .CK(clk_80mhz), 
            .Q(integrator2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i66.GSR = "ENABLED";
    FD1S3AX integrator2_i65 (.D(integrator2_71__N_1032[65]), .CK(clk_80mhz), 
            .Q(integrator2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i65.GSR = "ENABLED";
    LUT4 comb10_71__I_0_77_i137_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n67), .D(\comb10[65] ), .Z(n137_adj_3194)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i137_3_lut_4_lut.init = 16'hf960;
    FD1S3AX integrator2_i64 (.D(integrator2_71__N_1032[64]), .CK(clk_80mhz), 
            .Q(integrator2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i64.GSR = "ENABLED";
    FD1S3AX integrator2_i63 (.D(integrator2_71__N_1032[63]), .CK(clk_80mhz), 
            .Q(integrator2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i63.GSR = "ENABLED";
    FD1S3AX integrator2_i62 (.D(integrator2_71__N_1032[62]), .CK(clk_80mhz), 
            .Q(integrator2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i62.GSR = "ENABLED";
    FD1S3AX integrator2_i61 (.D(integrator2_71__N_1032[61]), .CK(clk_80mhz), 
            .Q(integrator2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i61.GSR = "ENABLED";
    FD1S3AX integrator2_i60 (.D(integrator2_71__N_1032[60]), .CK(clk_80mhz), 
            .Q(integrator2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i60.GSR = "ENABLED";
    FD1S3AX integrator2_i59 (.D(integrator2_71__N_1032[59]), .CK(clk_80mhz), 
            .Q(integrator2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i59.GSR = "ENABLED";
    FD1S3AX integrator2_i58 (.D(integrator2_71__N_1032[58]), .CK(clk_80mhz), 
            .Q(integrator2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i58.GSR = "ENABLED";
    FD1S3AX integrator2_i57 (.D(integrator2_71__N_1032[57]), .CK(clk_80mhz), 
            .Q(integrator2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i57.GSR = "ENABLED";
    FD1S3AX integrator2_i56 (.D(integrator2_71__N_1032[56]), .CK(clk_80mhz), 
            .Q(integrator2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i56.GSR = "ENABLED";
    FD1S3AX integrator2_i55 (.D(integrator2_71__N_1032[55]), .CK(clk_80mhz), 
            .Q(integrator2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i55.GSR = "ENABLED";
    FD1S3AX integrator2_i54 (.D(integrator2_71__N_1032[54]), .CK(clk_80mhz), 
            .Q(integrator2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i54.GSR = "ENABLED";
    FD1S3AX integrator2_i53 (.D(integrator2_71__N_1032[53]), .CK(clk_80mhz), 
            .Q(integrator2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i53.GSR = "ENABLED";
    FD1S3AX integrator2_i52 (.D(integrator2_71__N_1032[52]), .CK(clk_80mhz), 
            .Q(integrator2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i52.GSR = "ENABLED";
    FD1S3AX integrator2_i51 (.D(integrator2_71__N_1032[51]), .CK(clk_80mhz), 
            .Q(integrator2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i51.GSR = "ENABLED";
    FD1S3AX integrator2_i50 (.D(integrator2_71__N_1032[50]), .CK(clk_80mhz), 
            .Q(integrator2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i50.GSR = "ENABLED";
    FD1S3AX integrator2_i49 (.D(integrator2_71__N_1032[49]), .CK(clk_80mhz), 
            .Q(integrator2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i49.GSR = "ENABLED";
    FD1S3AX integrator2_i48 (.D(integrator2_71__N_1032[48]), .CK(clk_80mhz), 
            .Q(integrator2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i48.GSR = "ENABLED";
    FD1S3AX integrator2_i47 (.D(integrator2_71__N_1032[47]), .CK(clk_80mhz), 
            .Q(integrator2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i47.GSR = "ENABLED";
    FD1S3AX integrator2_i46 (.D(integrator2_71__N_1032[46]), .CK(clk_80mhz), 
            .Q(integrator2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i46.GSR = "ENABLED";
    FD1S3AX integrator2_i45 (.D(integrator2_71__N_1032[45]), .CK(clk_80mhz), 
            .Q(integrator2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i45.GSR = "ENABLED";
    FD1S3AX integrator2_i44 (.D(integrator2_71__N_1032[44]), .CK(clk_80mhz), 
            .Q(integrator2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i44.GSR = "ENABLED";
    FD1S3AX integrator2_i43 (.D(integrator2_71__N_1032[43]), .CK(clk_80mhz), 
            .Q(integrator2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i43.GSR = "ENABLED";
    FD1S3AX integrator2_i42 (.D(integrator2_71__N_1032[42]), .CK(clk_80mhz), 
            .Q(integrator2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i42.GSR = "ENABLED";
    FD1S3AX integrator2_i41 (.D(integrator2_71__N_1032[41]), .CK(clk_80mhz), 
            .Q(integrator2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i41.GSR = "ENABLED";
    FD1S3AX integrator2_i40 (.D(integrator2_71__N_1032[40]), .CK(clk_80mhz), 
            .Q(integrator2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i40.GSR = "ENABLED";
    FD1S3AX integrator2_i39 (.D(integrator2_71__N_1032[39]), .CK(clk_80mhz), 
            .Q(integrator2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i39.GSR = "ENABLED";
    FD1S3AX integrator2_i38 (.D(integrator2_71__N_1032[38]), .CK(clk_80mhz), 
            .Q(integrator2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i38.GSR = "ENABLED";
    FD1S3AX integrator2_i37 (.D(integrator2_71__N_1032[37]), .CK(clk_80mhz), 
            .Q(integrator2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i37.GSR = "ENABLED";
    FD1S3AX integrator2_i36 (.D(integrator2_71__N_1032[36]), .CK(clk_80mhz), 
            .Q(integrator2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i36.GSR = "ENABLED";
    FD1S3AX integrator2_i35 (.D(integrator2_71__N_1032[35]), .CK(clk_80mhz), 
            .Q(integrator2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i35.GSR = "ENABLED";
    FD1S3AX integrator2_i34 (.D(integrator2_71__N_1032[34]), .CK(clk_80mhz), 
            .Q(integrator2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i34.GSR = "ENABLED";
    FD1S3AX integrator2_i33 (.D(integrator2_71__N_1032[33]), .CK(clk_80mhz), 
            .Q(integrator2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i33.GSR = "ENABLED";
    FD1S3AX integrator2_i32 (.D(integrator2_71__N_1032[32]), .CK(clk_80mhz), 
            .Q(integrator2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i32.GSR = "ENABLED";
    FD1S3AX integrator2_i31 (.D(integrator2_71__N_1032[31]), .CK(clk_80mhz), 
            .Q(integrator2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i31.GSR = "ENABLED";
    FD1S3AX integrator2_i30 (.D(integrator2_71__N_1032[30]), .CK(clk_80mhz), 
            .Q(integrator2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i30.GSR = "ENABLED";
    FD1S3AX integrator2_i29 (.D(integrator2_71__N_1032[29]), .CK(clk_80mhz), 
            .Q(integrator2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i29.GSR = "ENABLED";
    FD1S3AX integrator2_i28 (.D(integrator2_71__N_1032[28]), .CK(clk_80mhz), 
            .Q(integrator2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i28.GSR = "ENABLED";
    FD1S3AX integrator2_i27 (.D(integrator2_71__N_1032[27]), .CK(clk_80mhz), 
            .Q(integrator2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i27.GSR = "ENABLED";
    FD1S3AX integrator2_i26 (.D(integrator2_71__N_1032[26]), .CK(clk_80mhz), 
            .Q(integrator2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i26.GSR = "ENABLED";
    FD1S3AX integrator2_i25 (.D(integrator2_71__N_1032[25]), .CK(clk_80mhz), 
            .Q(integrator2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i25.GSR = "ENABLED";
    FD1S3AX integrator2_i24 (.D(integrator2_71__N_1032[24]), .CK(clk_80mhz), 
            .Q(integrator2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i24.GSR = "ENABLED";
    FD1S3AX integrator2_i23 (.D(integrator2_71__N_1032[23]), .CK(clk_80mhz), 
            .Q(integrator2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i23.GSR = "ENABLED";
    FD1S3AX integrator2_i22 (.D(integrator2_71__N_1032[22]), .CK(clk_80mhz), 
            .Q(integrator2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i22.GSR = "ENABLED";
    FD1S3AX integrator2_i21 (.D(integrator2_71__N_1032[21]), .CK(clk_80mhz), 
            .Q(integrator2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i21.GSR = "ENABLED";
    FD1S3AX integrator2_i20 (.D(integrator2_71__N_1032[20]), .CK(clk_80mhz), 
            .Q(integrator2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i20.GSR = "ENABLED";
    FD1S3AX integrator2_i19 (.D(integrator2_71__N_1032[19]), .CK(clk_80mhz), 
            .Q(integrator2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i19.GSR = "ENABLED";
    FD1S3AX integrator2_i18 (.D(integrator2_71__N_1032[18]), .CK(clk_80mhz), 
            .Q(integrator2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i18.GSR = "ENABLED";
    FD1S3AX integrator2_i17 (.D(integrator2_71__N_1032[17]), .CK(clk_80mhz), 
            .Q(integrator2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i17.GSR = "ENABLED";
    FD1S3AX integrator2_i16 (.D(integrator2_71__N_1032[16]), .CK(clk_80mhz), 
            .Q(integrator2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i16.GSR = "ENABLED";
    FD1S3AX integrator2_i15 (.D(integrator2_71__N_1032[15]), .CK(clk_80mhz), 
            .Q(integrator2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i15.GSR = "ENABLED";
    FD1S3AX integrator2_i14 (.D(integrator2_71__N_1032[14]), .CK(clk_80mhz), 
            .Q(integrator2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i14.GSR = "ENABLED";
    FD1S3AX integrator2_i13 (.D(integrator2_71__N_1032[13]), .CK(clk_80mhz), 
            .Q(integrator2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i13.GSR = "ENABLED";
    FD1S3AX integrator2_i12 (.D(integrator2_71__N_1032[12]), .CK(clk_80mhz), 
            .Q(integrator2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i12.GSR = "ENABLED";
    FD1S3AX integrator2_i11 (.D(integrator2_71__N_1032[11]), .CK(clk_80mhz), 
            .Q(integrator2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i11.GSR = "ENABLED";
    FD1S3AX integrator2_i10 (.D(integrator2_71__N_1032[10]), .CK(clk_80mhz), 
            .Q(integrator2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i10.GSR = "ENABLED";
    FD1S3AX integrator2_i9 (.D(integrator2_71__N_1032[9]), .CK(clk_80mhz), 
            .Q(integrator2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i9.GSR = "ENABLED";
    FD1S3AX integrator2_i8 (.D(integrator2_71__N_1032[8]), .CK(clk_80mhz), 
            .Q(integrator2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i8.GSR = "ENABLED";
    FD1S3AX integrator2_i7 (.D(integrator2_71__N_1032[7]), .CK(clk_80mhz), 
            .Q(integrator2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i7.GSR = "ENABLED";
    FD1S3AX integrator2_i6 (.D(integrator2_71__N_1032[6]), .CK(clk_80mhz), 
            .Q(integrator2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i6.GSR = "ENABLED";
    FD1S3AX integrator2_i5 (.D(integrator2_71__N_1032[5]), .CK(clk_80mhz), 
            .Q(integrator2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i5.GSR = "ENABLED";
    FD1S3AX integrator2_i4 (.D(integrator2_71__N_1032[4]), .CK(clk_80mhz), 
            .Q(integrator2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i4.GSR = "ENABLED";
    FD1S3AX integrator2_i3 (.D(integrator2_71__N_1032[3]), .CK(clk_80mhz), 
            .Q(integrator2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i3.GSR = "ENABLED";
    FD1S3AX integrator2_i2 (.D(integrator2_71__N_1032[2]), .CK(clk_80mhz), 
            .Q(integrator2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i2.GSR = "ENABLED";
    FD1S3AX integrator2_i1 (.D(integrator2_71__N_1032[1]), .CK(clk_80mhz), 
            .Q(integrator2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i1.GSR = "ENABLED";
    LUT4 mux_3408_i6_3_lut (.A(n106), .B(n108), .C(cout), .Z(comb10_71__N_2281[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i6_3_lut.init = 16'hcaca;
    LUT4 mux_3408_i5_3_lut (.A(n109), .B(n111), .C(cout), .Z(comb10_71__N_2281[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i5_3_lut.init = 16'hcaca;
    LUT4 comb10_71__I_0_77_i136_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n66), .D(\comb10[64] ), .Z(n136)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i136_3_lut_4_lut.init = 16'hf960;
    LUT4 mux_3408_i4_3_lut (.A(n112), .B(n114), .C(cout), .Z(comb10_71__N_2281[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3408_i3_3_lut (.A(n115), .B(n117), .C(cout), .Z(comb10_71__N_2281[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i3_3_lut.init = 16'hcaca;
    LUT4 mux_3408_i2_3_lut (.A(n118), .B(n120), .C(cout), .Z(comb10_71__N_2281[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3408_i2_3_lut.init = 16'hcaca;
    LUT4 comb10_71__I_0_77_i68_3_lut (.A(comb10[67]), .B(comb10[68]), .C(\cic_gain[0] ), 
         .Z(n68_adj_3196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i68_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_207 (.A(n67_adj_228[0]), .B(n73), .Z(count_11__N_1980[0])) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_207.init = 16'hbbbb;
    LUT4 comb10_71__I_0_77_i65_3_lut (.A(comb10[64]), .B(comb10[65]), .C(\cic_gain[0] ), 
         .Z(n65_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i65_3_lut.init = 16'hcaca;
    LUT4 comb10_71__I_0_77_i134_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n64), .D(\comb10[62] ), .Z(n134)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i134_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_29_inv_0_i55_1_lut (.A(comb_d8[54]), .Z(n19_adj_159)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 comb10_71__I_0_77_i133_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n63), .D(\comb10[61] ), .Z(n133)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i133_3_lut_4_lut.init = 16'hf960;
    LUT4 comb10_71__I_0_77_i135_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n65), .D(\comb10[63] ), .Z(n135)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i135_3_lut_4_lut.init = 16'hf960;
    LUT4 comb10_71__I_0_77_i70_3_lut (.A(comb10[69]), .B(comb10[70]), .C(\cic_gain[0] ), 
         .Z(n70_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i70_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i67_1_lut (.A(integrator_d_tmp[66]), .Z(n7_adj_160)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i68_1_lut (.A(integrator_d_tmp[67]), .Z(n6_adj_161)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i61_1_lut (.A(integrator_d_tmp[60]), .Z(n13_adj_162)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i62_1_lut (.A(integrator_d_tmp[61]), .Z(n12_adj_163)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i53_1_lut (.A(integrator_d_tmp[52]), .Z(n21_adj_164)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i54_1_lut (.A(integrator_d_tmp[53]), .Z(n20_adj_165)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i59_1_lut (.A(integrator_d_tmp[58]), .Z(n15_adj_166)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i60_1_lut (.A(integrator_d_tmp[59]), .Z(n14_adj_167)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i51_1_lut (.A(integrator_d_tmp[50]), .Z(n23_adj_168)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i52_1_lut (.A(integrator_d_tmp[51]), .Z(n22_adj_169)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i65_1_lut (.A(integrator_d_tmp[64]), .Z(n9_adj_170)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i66_1_lut (.A(integrator_d_tmp[65]), .Z(n8_adj_171)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i57_1_lut (.A(integrator_d_tmp[56]), .Z(n17_adj_172)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i58_1_lut (.A(integrator_d_tmp[57]), .Z(n16_adj_173)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i49_1_lut (.A(integrator_d_tmp[48]), .Z(n25_adj_174)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i50_1_lut (.A(integrator_d_tmp[49]), .Z(n24_adj_175)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i63_1_lut (.A(integrator_d_tmp[62]), .Z(n11_adj_176)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i64_1_lut (.A(integrator_d_tmp[63]), .Z(n10_adj_177)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i55_1_lut (.A(integrator_d_tmp[54]), .Z(n19_adj_178)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i56_1_lut (.A(integrator_d_tmp[55]), .Z(n18_adj_179)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i47_1_lut (.A(integrator_d_tmp[46]), .Z(n27_adj_180)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i48_1_lut (.A(integrator_d_tmp[47]), .Z(n26_adj_181)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i41_1_lut (.A(integrator_d_tmp[40]), .Z(n33_adj_182)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i42_1_lut (.A(integrator_d_tmp[41]), .Z(n32_adj_183)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i39_1_lut (.A(integrator_d_tmp[38]), .Z(n35_adj_184)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i40_1_lut (.A(integrator_d_tmp[39]), .Z(n34_adj_185)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i45_1_lut (.A(integrator_d_tmp[44]), .Z(n29_adj_186)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i46_1_lut (.A(integrator_d_tmp[45]), .Z(n28_adj_187)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i37_1_lut (.A(integrator_d_tmp[36]), .Z(n37_adj_188)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i38_1_lut (.A(integrator_d_tmp[37]), .Z(n36_adj_189)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i71_1_lut (.A(comb_d6[70]), .Z(n3_adj_190)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i72_1_lut (.A(comb_d6[71]), .Z(n2_adj_191)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i43_1_lut (.A(integrator_d_tmp[42]), .Z(n31_adj_192)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i44_1_lut (.A(integrator_d_tmp[43]), .Z(n30_adj_193)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i69_1_lut (.A(comb_d6[68]), .Z(n5_adj_194)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i70_1_lut (.A(comb_d6[69]), .Z(n4_adj_195)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i63_1_lut (.A(comb_d6[62]), .Z(n11_adj_196)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i64_1_lut (.A(comb_d6[63]), .Z(n10_adj_197)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i57_1_lut (.A(comb_d6[56]), .Z(n17_adj_198)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i58_1_lut (.A(comb_d6[57]), .Z(n16_adj_199)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i61_1_lut (.A(comb_d6[60]), .Z(n13_adj_200)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i62_1_lut (.A(comb_d6[61]), .Z(n12_adj_201)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i67_1_lut (.A(comb_d6[66]), .Z(n7_adj_202)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i67_1_lut.init = 16'h5555;
    FD1P3AX integrator_tmp_i0_i0 (.D(integrator5[0]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i0.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i68_1_lut (.A(comb_d6[67]), .Z(n6_adj_203)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i59_1_lut (.A(comb_d6[58]), .Z(n15_adj_204)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i60_1_lut (.A(comb_d6[59]), .Z(n14_adj_205)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 comb10_71__I_0_77_i131_3_lut_4_lut_adj_208 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n61_adj_206), .D(\comb10[59] ), .Z(n131_adj_3252)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i131_3_lut_4_lut_adj_208.init = 16'hf960;
    LUT4 sub_27_inv_0_i55_1_lut (.A(comb_d6[54]), .Z(n19_adj_207)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i56_1_lut (.A(comb_d6[55]), .Z(n18_adj_208)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i65_1_lut (.A(comb_d6[64]), .Z(n9_adj_209)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i66_1_lut (.A(comb_d6[65]), .Z(n8_adj_210)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i53_1_lut (.A(comb_d6[52]), .Z(n21_adj_211)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 comb10_71__I_0_77_i208_3_lut_4_lut (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n68_adj_3196), .D(n136_adj_3258), .Z(led_0_1)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i208_3_lut_4_lut.init = 16'hfe10;
    LUT4 comb10_71__I_0_77_i207_3_lut_4_lut (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n67_c), .D(n135_adj_3259), .Z(led_0_0)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i207_3_lut_4_lut.init = 16'hfe10;
    LUT4 comb10_71__I_0_77_i206_3_lut_4_lut (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n66_adj_3260), .D(n134_adj_3261), .Z(\cic_sine_out[5] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i206_3_lut_4_lut.init = 16'hfe10;
    LUT4 sub_28_inv_0_i67_1_lut (.A(comb_d7[66]), .Z(n7_adj_212)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i68_1_lut (.A(comb_d7[67]), .Z(n6_adj_213)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i61_1_lut (.A(comb_d7[60]), .Z(n13_adj_214)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 comb10_71__I_0_77_i140_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n70_c), .D(comb10[68]), .Z(n140)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i140_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_28_inv_0_i62_1_lut (.A(comb_d7[61]), .Z(n12_adj_215)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i59_1_lut (.A(comb_d7[58]), .Z(n15_adj_216)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 comb10_71__I_0_77_i205_3_lut_4_lut (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n65_c), .D(n133_adj_3267), .Z(\cic_sine_out[4] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i205_3_lut_4_lut.init = 16'hfe10;
    LUT4 comb10_71__I_0_77_i138_3_lut_4_lut_adj_209 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n68_adj_3196), .D(comb10[66]), .Z(n138_adj_3268)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i138_3_lut_4_lut_adj_209.init = 16'hf960;
    LUT4 comb10_71__I_0_77_i204_3_lut_4_lut (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n64_adj_3269), .D(n132_adj_3270), .Z(\cic_sine_out[3] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i204_3_lut_4_lut.init = 16'hfe10;
    LUT4 comb10_71__I_0_77_i203_3_lut_4_lut (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n63_c), .D(n131), .Z(\cic_sine_out[2] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i203_3_lut_4_lut.init = 16'hfe10;
    LUT4 comb10_71__I_0_77_i132_3_lut_4_lut_adj_210 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n62_c), .D(comb10[60]), .Z(n132_adj_3270)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i132_3_lut_4_lut_adj_210.init = 16'hf960;
    LUT4 comb10_71__I_0_77_i212_3_lut_4_lut (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(\comb10[71] ), .D(n140_adj_3272), .Z(\cic_cosine_out[11] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i212_3_lut_4_lut.init = 16'hfe10;
    LUT4 comb10_71__I_0_77_i136_3_lut_4_lut_adj_211 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n66_adj_3260), .D(comb10[64]), .Z(n136_adj_3258)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i136_3_lut_4_lut_adj_211.init = 16'hf960;
    FD1P3AX integrator_tmp_i0_i1 (.D(integrator5[1]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i1.GSR = "ENABLED";
    LUT4 comb10_71__I_0_77_i210_3_lut_4_lut (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n70), .D(n138), .Z(\cic_cosine_out[9] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i210_3_lut_4_lut.init = 16'hfe10;
    LUT4 comb10_71__I_0_77_i141_3_lut_4_lut (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n137_adj_3194), .D(\comb10[68] ), .Z(\cic_cosine_out[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i141_3_lut_4_lut.init = 16'hf1e0;
    LUT4 comb10_71__I_0_77_i208_3_lut_4_lut_adj_212 (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n68), .D(n136), .Z(\cic_cosine_out[7] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i208_3_lut_4_lut_adj_212.init = 16'hfe10;
    LUT4 comb10_71__I_0_77_i133_3_lut_4_lut_adj_213 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n63_c), .D(comb10[61]), .Z(n133_adj_3267)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i133_3_lut_4_lut_adj_213.init = 16'hf960;
    LUT4 comb10_71__I_0_77_i207_3_lut_4_lut_adj_214 (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n67), .D(n135), .Z(\cic_cosine_out[6] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i207_3_lut_4_lut_adj_214.init = 16'hfe10;
    FD1S3AX valid_comb_63_rep_294 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_291)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_294.GSR = "ENABLED";
    LUT4 comb10_71__I_0_77_i137_3_lut_4_lut_adj_215 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n67_c), .D(comb10[65]), .Z(n137)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i137_3_lut_4_lut_adj_215.init = 16'hf960;
    LUT4 comb10_71__I_0_77_i140_3_lut_4_lut_adj_216 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n70), .D(\comb10[68] ), .Z(n140_adj_3272)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i140_3_lut_4_lut_adj_216.init = 16'hf960;
    LUT4 comb10_71__I_0_77_i206_3_lut_4_lut_adj_217 (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n66), .D(n134), .Z(\cic_cosine_out[5] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i206_3_lut_4_lut_adj_217.init = 16'hfe10;
    LUT4 comb10_71__I_0_77_i134_3_lut_4_lut_adj_218 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n64_adj_3269), .D(comb10[62]), .Z(n134_adj_3261)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i134_3_lut_4_lut_adj_218.init = 16'hf960;
    LUT4 comb10_71__I_0_77_i205_3_lut_4_lut_adj_219 (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n65), .D(n133), .Z(\cic_cosine_out[4] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i205_3_lut_4_lut_adj_219.init = 16'hfe10;
    LUT4 comb10_71__I_0_77_i204_3_lut_4_lut_adj_220 (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n64), .D(n132), .Z(\cic_cosine_out[3] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i204_3_lut_4_lut_adj_220.init = 16'hfe10;
    LUT4 comb10_71__I_0_77_i203_3_lut_4_lut_adj_221 (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n63), .D(n131_adj_3252), .Z(\cic_cosine_out[2] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i203_3_lut_4_lut_adj_221.init = 16'hfe10;
    LUT4 i8526_then_3_lut (.A(\cic_gain[1] ), .B(comb10[59]), .C(comb10[57]), 
         .Z(n19851)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i8526_then_3_lut.init = 16'he4e4;
    LUT4 comb10_71__I_0_77_i212_3_lut_4_lut_adj_222 (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(comb10[71]), .D(n140), .Z(led_0_5)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i212_3_lut_4_lut_adj_222.init = 16'hfe10;
    LUT4 comb10_71__I_0_77_i210_3_lut_4_lut_adj_223 (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(n70_c), .D(n138_adj_3268), .Z(led_0_3)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i210_3_lut_4_lut_adj_223.init = 16'hfe10;
    LUT4 i8526_else_3_lut (.A(n61), .B(\cic_gain[1] ), .C(comb10[58]), 
         .Z(n19850)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i8526_else_3_lut.init = 16'he2e2;
    LUT4 comb10_71__I_0_77_i135_3_lut_4_lut_adj_224 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n65_c), .D(comb10[63]), .Z(n135_adj_3259)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam comb10_71__I_0_77_i135_3_lut_4_lut_adj_224.init = 16'hf960;
    LUT4 comb10_71__I_0_77_i66_3_lut (.A(comb10[65]), .B(comb10[66]), .C(\cic_gain[0] ), 
         .Z(n66_adj_3260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i66_3_lut.init = 16'hcaca;
    LUT4 comb10_71__I_0_77_i64_3_lut (.A(comb10[63]), .B(comb10[64]), .C(\cic_gain[0] ), 
         .Z(n64_adj_3269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i64_3_lut.init = 16'hcaca;
    LUT4 sub_29_inv_0_i56_1_lut (.A(comb_d8[55]), .Z(n18_adj_217)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i63_1_lut (.A(comb_d7[62]), .Z(n11_adj_218)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i64_1_lut (.A(comb_d7[63]), .Z(n10_adj_219)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i41_1_lut (.A(comb_d7[40]), .Z(n33_adj_220)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i42_1_lut (.A(comb_d7[41]), .Z(n32_adj_221)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i65_1_lut (.A(comb_d8[64]), .Z(n9_adj_222)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 i8697_then_3_lut (.A(\cic_gain[1] ), .B(comb10[60]), .C(comb10[58]), 
         .Z(n19860)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i8697_then_3_lut.init = 16'he4e4;
    LUT4 i8697_else_3_lut (.A(n62_c), .B(\cic_gain[1] ), .C(comb10[59]), 
         .Z(n19859)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i8697_else_3_lut.init = 16'he2e2;
    LUT4 sub_29_inv_0_i66_1_lut (.A(comb_d8[65]), .Z(n8_adj_223)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i66_1_lut.init = 16'h5555;
    PFUMX i8773 (.BLUT(n19871), .ALUT(n19872), .C0(\cic_gain[0] ), .Z(\cic_cosine_out[10] ));
    PFUMX i8771 (.BLUT(n19868), .ALUT(n19869), .C0(\cic_gain[0] ), .Z(led_0_4));
    PFUMX i8765 (.BLUT(n19859), .ALUT(n19860), .C0(\cic_gain[0] ), .Z(\cic_sine_out[1] ));
    FD1P3AX integrator_tmp_i0_i2 (.D(integrator5[2]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i3 (.D(integrator5[3]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i4 (.D(integrator5[4]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i5 (.D(integrator5[5]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i6 (.D(integrator5[6]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i7 (.D(integrator5[7]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i8 (.D(integrator5[8]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i9 (.D(integrator5[9]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i10 (.D(integrator5[10]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i11 (.D(integrator5[11]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i12 (.D(integrator5[12]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i13 (.D(integrator5[13]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i14 (.D(integrator5[14]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i15 (.D(integrator5[15]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i16 (.D(integrator5[16]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i17 (.D(integrator5[17]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i18 (.D(integrator5[18]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i19 (.D(integrator5[19]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i20 (.D(integrator5[20]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i21 (.D(integrator5[21]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i22 (.D(integrator5[22]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i23 (.D(integrator5[23]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i24 (.D(integrator5[24]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i25 (.D(integrator5[25]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i26 (.D(integrator5[26]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i27 (.D(integrator5[27]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i28 (.D(integrator5[28]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i29 (.D(integrator5[29]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i30 (.D(integrator5[30]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i31 (.D(integrator5[31]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i32 (.D(integrator5[32]), .SP(clk_80mhz_enable_1456), 
            .CK(clk_80mhz), .Q(integrator_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i33 (.D(integrator5[33]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i34 (.D(integrator5[34]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i35 (.D(integrator5[35]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i36 (.D(integrator5[36]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i37 (.D(integrator5[37]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i38 (.D(integrator5[38]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i39 (.D(integrator5[39]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i40 (.D(integrator5[40]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i41 (.D(integrator5[41]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i42 (.D(integrator5[42]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i43 (.D(integrator5[43]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i44 (.D(integrator5[44]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i45 (.D(integrator5[45]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i46 (.D(integrator5[46]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i47 (.D(integrator5[47]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i48 (.D(integrator5[48]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i49 (.D(integrator5[49]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i50 (.D(integrator5[50]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i51 (.D(integrator5[51]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i52 (.D(integrator5[52]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i53 (.D(integrator5[53]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i54 (.D(integrator5[54]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i55 (.D(integrator5[55]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i56 (.D(integrator5[56]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i57 (.D(integrator5[57]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i58 (.D(integrator5[58]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i59 (.D(integrator5[59]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i60 (.D(integrator5[60]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i61 (.D(integrator5[61]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i62 (.D(integrator5[62]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i63 (.D(integrator5[63]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i64 (.D(integrator5[64]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i65 (.D(integrator5[65]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i66 (.D(integrator5[66]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i67 (.D(integrator5[67]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i68 (.D(integrator5[68]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i69 (.D(integrator5[69]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i70 (.D(integrator5[70]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i71 (.D(integrator5[71]), .SP(decimation_clk_N_2353), 
            .CK(clk_80mhz), .Q(integrator_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i71.GSR = "ENABLED";
    PFUMX i8759 (.BLUT(n19850), .ALUT(n19851), .C0(\cic_gain[0] ), .Z(\cic_sine_out[0] ));
    FD1S3IX count__i10 (.D(n67_adj_228[10]), .CK(clk_80mhz), .CD(n14270), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i10.GSR = "ENABLED";
    LUT4 sub_29_inv_0_i47_1_lut (.A(comb_d8[46]), .Z(n27_adj_224)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i48_1_lut (.A(comb_d8[47]), .Z(n26_adj_225)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i48_1_lut.init = 16'h5555;
    FD1S3AX valid_comb_63_rep_306 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1423)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_306.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_305 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1373)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_305.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_304 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1323)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_304.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_303 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1273)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_303.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_302 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1223)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_302.GSR = "ENABLED";
    LUT4 sub_29_inv_0_i39_1_lut (.A(comb_d8[38]), .Z(n35_adj_226)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i39_1_lut.init = 16'h5555;
    FD1S3AX valid_comb_63_rep_301 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1173)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_301.GSR = "ENABLED";
    LUT4 sub_29_inv_0_i40_1_lut (.A(comb_d8[39]), .Z(n34_adj_227)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i40_1_lut.init = 16'h5555;
    FD1S3AX valid_comb_63_rep_300 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1123)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_300.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_299 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1073)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_299.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_298 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1023)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_298.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_297 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_973)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_297.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_296 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_923)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_296.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_295 (.D(clk_80mhz_enable_1456), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_873)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=190, LSE_RLINE=196 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_295.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module PWM
//

module PWM (\data_in_reg[0] , clk_80mhz, \data_in_reg_11__N_2898[0] , 
            \data_in_reg[9] , \data_in_reg[8] , \data_in_reg_11__N_2898[8] , 
            \data_in_reg[7] , \data_in_reg_11__N_2898[7] , \data_in_reg[6] , 
            \data_in_reg_11__N_2898[6] , \data_in_reg[5] , \data_in_reg_11__N_2898[5] , 
            \data_in_reg[4] , \data_in_reg_11__N_2898[4] , \data_in_reg[3] , 
            \data_in_reg_11__N_2898[3] , \data_in_reg[2] , \data_in_reg_11__N_2898[2] , 
            \data_in_reg[1] , \data_in_reg_11__N_2898[1] , count, \amdemod_out[9] , 
            GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    output \data_in_reg[0] ;
    input clk_80mhz;
    input \data_in_reg_11__N_2898[0] ;
    output \data_in_reg[9] ;
    output \data_in_reg[8] ;
    input \data_in_reg_11__N_2898[8] ;
    output \data_in_reg[7] ;
    input \data_in_reg_11__N_2898[7] ;
    output \data_in_reg[6] ;
    input \data_in_reg_11__N_2898[6] ;
    output \data_in_reg[5] ;
    input \data_in_reg_11__N_2898[5] ;
    output \data_in_reg[4] ;
    input \data_in_reg_11__N_2898[4] ;
    output \data_in_reg[3] ;
    input \data_in_reg_11__N_2898[3] ;
    output \data_in_reg[2] ;
    input \data_in_reg_11__N_2898[2] ;
    output \data_in_reg[1] ;
    input \data_in_reg_11__N_2898[1] ;
    output [9:0]count;
    input \amdemod_out[9] ;
    input GND_net;
    input VCC_net;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(61[34:43])
    
    wire clk_80mhz_enable_30;
    wire [11:0]n4469;
    
    wire n17, n15, n11, n12;
    wire [9:0]n45;
    
    wire n17667, n17666, n17665, n17664, n17663;
    
    FD1P3AX data_in_reg__i1 (.D(\data_in_reg_11__N_2898[0] ), .SP(clk_80mhz_enable_30), 
            .CK(clk_80mhz), .Q(\data_in_reg[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=5, LSE_LLINE=233, LSE_RLINE=237 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(46[10] 61[6])
    defparam data_in_reg__i1.GSR = "ENABLED";
    FD1P3AX data_in_reg__i10 (.D(n4469[9]), .SP(clk_80mhz_enable_30), .CK(clk_80mhz), 
            .Q(\data_in_reg[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=5, LSE_LLINE=233, LSE_RLINE=237 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(46[10] 61[6])
    defparam data_in_reg__i10.GSR = "ENABLED";
    FD1P3AX data_in_reg__i9 (.D(\data_in_reg_11__N_2898[8] ), .SP(clk_80mhz_enable_30), 
            .CK(clk_80mhz), .Q(\data_in_reg[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=5, LSE_LLINE=233, LSE_RLINE=237 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(46[10] 61[6])
    defparam data_in_reg__i9.GSR = "ENABLED";
    FD1P3AX data_in_reg__i8 (.D(\data_in_reg_11__N_2898[7] ), .SP(clk_80mhz_enable_30), 
            .CK(clk_80mhz), .Q(\data_in_reg[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=5, LSE_LLINE=233, LSE_RLINE=237 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(46[10] 61[6])
    defparam data_in_reg__i8.GSR = "ENABLED";
    FD1P3AX data_in_reg__i7 (.D(\data_in_reg_11__N_2898[6] ), .SP(clk_80mhz_enable_30), 
            .CK(clk_80mhz), .Q(\data_in_reg[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=5, LSE_LLINE=233, LSE_RLINE=237 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(46[10] 61[6])
    defparam data_in_reg__i7.GSR = "ENABLED";
    FD1P3AX data_in_reg__i6 (.D(\data_in_reg_11__N_2898[5] ), .SP(clk_80mhz_enable_30), 
            .CK(clk_80mhz), .Q(\data_in_reg[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=5, LSE_LLINE=233, LSE_RLINE=237 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(46[10] 61[6])
    defparam data_in_reg__i6.GSR = "ENABLED";
    FD1P3AX data_in_reg__i5 (.D(\data_in_reg_11__N_2898[4] ), .SP(clk_80mhz_enable_30), 
            .CK(clk_80mhz), .Q(\data_in_reg[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=5, LSE_LLINE=233, LSE_RLINE=237 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(46[10] 61[6])
    defparam data_in_reg__i5.GSR = "ENABLED";
    FD1P3AX data_in_reg__i4 (.D(\data_in_reg_11__N_2898[3] ), .SP(clk_80mhz_enable_30), 
            .CK(clk_80mhz), .Q(\data_in_reg[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=5, LSE_LLINE=233, LSE_RLINE=237 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(46[10] 61[6])
    defparam data_in_reg__i4.GSR = "ENABLED";
    FD1P3AX data_in_reg__i3 (.D(\data_in_reg_11__N_2898[2] ), .SP(clk_80mhz_enable_30), 
            .CK(clk_80mhz), .Q(\data_in_reg[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=5, LSE_LLINE=233, LSE_RLINE=237 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(46[10] 61[6])
    defparam data_in_reg__i3.GSR = "ENABLED";
    FD1P3AX data_in_reg__i2 (.D(\data_in_reg_11__N_2898[1] ), .SP(clk_80mhz_enable_30), 
            .CK(clk_80mhz), .Q(\data_in_reg[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=5, LSE_LLINE=233, LSE_RLINE=237 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(46[10] 61[6])
    defparam data_in_reg__i2.GSR = "ENABLED";
    LUT4 i8383_4_lut (.A(n17), .B(n15), .C(n11), .D(n12), .Z(clk_80mhz_enable_30)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(51[9:37])
    defparam i8383_4_lut.init = 16'h0001;
    LUT4 i7_4_lut (.A(count[3]), .B(count[2]), .C(count[1]), .D(count[9]), 
         .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(51[9:37])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(count[6]), .B(count[4]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(51[9:37])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(count[0]), .B(count[5]), .Z(n11)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(51[9:37])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2_2_lut (.A(count[7]), .B(count[8]), .Z(n12)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(51[9:37])
    defparam i2_2_lut.init = 16'heeee;
    FD1S3AX count_3038__i0 (.D(n45[0]), .CK(clk_80mhz), .Q(count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038__i0.GSR = "ENABLED";
    LUT4 i3343_1_lut (.A(\amdemod_out[9] ), .Z(n4469[9])) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(51[5] 53[8])
    defparam i3343_1_lut.init = 16'h5555;
    CCU2C count_3038_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17667), .S0(n45[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038_add_4_11.INIT0 = 16'haaa0;
    defparam count_3038_add_4_11.INIT1 = 16'h0000;
    defparam count_3038_add_4_11.INJECT1_0 = "NO";
    defparam count_3038_add_4_11.INJECT1_1 = "NO";
    CCU2C count_3038_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17666), .COUT(n17667), .S0(n45[7]), .S1(n45[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038_add_4_9.INIT0 = 16'haaa0;
    defparam count_3038_add_4_9.INIT1 = 16'haaa0;
    defparam count_3038_add_4_9.INJECT1_0 = "NO";
    defparam count_3038_add_4_9.INJECT1_1 = "NO";
    CCU2C count_3038_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17665), .COUT(n17666), .S0(n45[5]), .S1(n45[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038_add_4_7.INIT0 = 16'haaa0;
    defparam count_3038_add_4_7.INIT1 = 16'haaa0;
    defparam count_3038_add_4_7.INJECT1_0 = "NO";
    defparam count_3038_add_4_7.INJECT1_1 = "NO";
    CCU2C count_3038_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17664), .COUT(n17665), .S0(n45[3]), .S1(n45[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038_add_4_5.INIT0 = 16'haaa0;
    defparam count_3038_add_4_5.INIT1 = 16'haaa0;
    defparam count_3038_add_4_5.INJECT1_0 = "NO";
    defparam count_3038_add_4_5.INJECT1_1 = "NO";
    CCU2C count_3038_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n17663), .COUT(n17664), .S0(n45[1]), .S1(n45[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038_add_4_3.INIT0 = 16'haaa0;
    defparam count_3038_add_4_3.INIT1 = 16'haaa0;
    defparam count_3038_add_4_3.INJECT1_0 = "NO";
    defparam count_3038_add_4_3.INJECT1_1 = "NO";
    CCU2C count_3038_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n17663), .S1(n45[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038_add_4_1.INIT0 = 16'h0000;
    defparam count_3038_add_4_1.INIT1 = 16'h555f;
    defparam count_3038_add_4_1.INJECT1_0 = "NO";
    defparam count_3038_add_4_1.INJECT1_1 = "NO";
    FD1S3AX count_3038__i1 (.D(n45[1]), .CK(clk_80mhz), .Q(count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038__i1.GSR = "ENABLED";
    FD1S3AX count_3038__i2 (.D(n45[2]), .CK(clk_80mhz), .Q(count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038__i2.GSR = "ENABLED";
    FD1S3AX count_3038__i3 (.D(n45[3]), .CK(clk_80mhz), .Q(count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038__i3.GSR = "ENABLED";
    FD1S3AX count_3038__i4 (.D(n45[4]), .CK(clk_80mhz), .Q(count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038__i4.GSR = "ENABLED";
    FD1S3AX count_3038__i5 (.D(n45[5]), .CK(clk_80mhz), .Q(count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038__i5.GSR = "ENABLED";
    FD1S3AX count_3038__i6 (.D(n45[6]), .CK(clk_80mhz), .Q(count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038__i6.GSR = "ENABLED";
    FD1S3AX count_3038__i7 (.D(n45[7]), .CK(clk_80mhz), .Q(count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038__i7.GSR = "ENABLED";
    FD1S3AX count_3038__i8 (.D(n45[8]), .CK(clk_80mhz), .Q(count[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038__i8.GSR = "ENABLED";
    FD1S3AX count_3038__i9 (.D(n45[9]), .CK(clk_80mhz), .Q(count[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/PWM.v(48[14:26])
    defparam count_3038__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \CIC(REGISTER_WIDTH=72,DECIMATION_RATIO=4096)_U2 
//

module \CIC(REGISTER_WIDTH=72,DECIMATION_RATIO=4096)_U2  (n67_adj_114, \cic_gain[1] , 
            \comb10[60] , n62, \comb10[59] , integrator_tmp, clk_80mhz, 
            integrator5, integrator_d_tmp, integrator2, integrator2_71__N_1032, 
            integrator3, integrator3_71__N_1104, integrator4, integrator4_71__N_1176, 
            integrator5_71__N_1248, comb6, comb6_71__N_1993, comb_d6, 
            comb7, comb7_71__N_2065, comb_d7, comb8, comb8_71__N_2137, 
            comb_d8, comb9, comb9_71__N_2209, comb_d9, integrator1, 
            integrator1_71__N_960, n19, n18, n21, n20, n23, n22, 
            n25, n24, n27, n3, n2, n26, n5, n29, n28_adj_1, 
            n31_adj_2, \comb10[71] , \comb10[70] , \comb10[69] , \comb10[68] , 
            \comb10[67] , \comb10[66] , \comb10[65] , \comb10[64] , 
            \comb10[63] , \comb10[62] , \comb10[61] , n30, n33, n32, 
            n35, n4, n34_adj_3, n37_adj_4, n36, n7, n3_adj_5, 
            n6, n2_adj_6, n5_adj_7, n4_adj_8, n7_adj_9, n6_adj_10, 
            n9, n8, n5_adj_11, n11, \cic_gain[0] , n4_adj_12, n10, 
            n13, n12, n15, n14, n17, n16, n19_adj_13, n18_adj_14, 
            n21_adj_15, n20_adj_16, n23_adj_17, n22_adj_18, n25_adj_19, 
            n24_adj_20, n27_adj_21, n26_adj_22, n29_adj_23, n28_adj_24, 
            n7_adj_25, n31_adj_26, n6_adj_27, n30_adj_28, n33_adj_29, 
            n32_adj_30, n35_adj_31, n9_adj_32, n8_adj_33, n34_adj_34, 
            n37_adj_35, n36_adj_36, n3_adj_37, n2_adj_38, n11_adj_39, 
            n5_adj_40, n4_adj_41, n7_adj_42, n6_adj_43, n10_adj_44, 
            n9_adj_45, n8_adj_46, n11_adj_47, n10_adj_48, n13_adj_49, 
            n12_adj_50, n15_adj_51, n13_adj_52, n14_adj_53, n17_adj_54, 
            n16_adj_55, n19_adj_56, n12_adj_57, n18_adj_58, n15_adj_59, 
            n21_adj_60, count, n20_adj_61, n23_adj_62, n22_adj_63, 
            n25_adj_64, n24_adj_65, n27_adj_66, n26_adj_67, n29_adj_68, 
            n28_adj_69, n31_adj_70, n30_adj_71, n9_adj_72, n8_adj_73, 
            n33_adj_74, n11_adj_75, n10_adj_76, n32_adj_77, n35_adj_78, 
            n70, n68, n67, n66, n65, n64, n63, n34_adj_79, n37_adj_80, 
            n36_adj_81, n13_adj_82, n12_adj_83, n14_adj_84, n15_adj_85, 
            n17_adj_86, n16_adj_87, n14_adj_88, n19_adj_89, n18_adj_90, 
            n21_adj_91, n20_adj_92, n61_adj_93, n23_adj_94, n22_adj_95, 
            n25_adj_96, n17_adj_97, n16_adj_98, n24_adj_99, n27_adj_100, 
            n26_adj_101, n76, n78, cout, n79, n81, n82, n84, 
            n85, n87, n88, n90, n91, n93, n94, n96, n97, n99, 
            n100, n102, n103, n105, n106, n108, n109, n111, 
            n112, n114, n115, n117, n118, n120, n29_adj_102, n28_adj_103, 
            n2_adj_104, n3_adj_105, n31_adj_106, n30_adj_107, n33_adj_108, 
            n32_adj_109, n35_adj_110, n34_adj_111, n37_adj_112, n36_adj_113, 
            \cic_cosine_out[1] , \cic_cosine_out[0] ) /* synthesis syn_module_defined=1 */ ;
    input [11:0]n67_adj_114;
    input \cic_gain[1] ;
    output \comb10[60] ;
    output n62;
    output \comb10[59] ;
    output [71:0]integrator_tmp;
    input clk_80mhz;
    output [71:0]integrator5;
    output [71:0]integrator_d_tmp;
    output [71:0]integrator2;
    input [71:0]integrator2_71__N_1032;
    output [71:0]integrator3;
    input [71:0]integrator3_71__N_1104;
    output [71:0]integrator4;
    input [71:0]integrator4_71__N_1176;
    input [71:0]integrator5_71__N_1248;
    output [71:0]comb6;
    input [71:0]comb6_71__N_1993;
    output [71:0]comb_d6;
    output [71:0]comb7;
    input [71:0]comb7_71__N_2065;
    output [71:0]comb_d7;
    output [71:0]comb8;
    input [71:0]comb8_71__N_2137;
    output [71:0]comb_d8;
    output [71:0]comb9;
    input [71:0]comb9_71__N_2209;
    output [71:0]comb_d9;
    output [71:0]integrator1;
    input [71:0]integrator1_71__N_960;
    output n19;
    output n18;
    output n21;
    output n20;
    output n23;
    output n22;
    output n25;
    output n24;
    output n27;
    output n3;
    output n2;
    output n26;
    output n5;
    output n29;
    output n28_adj_1;
    output n31_adj_2;
    output \comb10[71] ;
    output \comb10[70] ;
    output \comb10[69] ;
    output \comb10[68] ;
    output \comb10[67] ;
    output \comb10[66] ;
    output \comb10[65] ;
    output \comb10[64] ;
    output \comb10[63] ;
    output \comb10[62] ;
    output \comb10[61] ;
    output n30;
    output n33;
    output n32;
    output n35;
    output n4;
    output n34_adj_3;
    output n37_adj_4;
    output n36;
    output n7;
    output n3_adj_5;
    output n6;
    output n2_adj_6;
    output n5_adj_7;
    output n4_adj_8;
    output n7_adj_9;
    output n6_adj_10;
    output n9;
    output n8;
    output n5_adj_11;
    output n11;
    input \cic_gain[0] ;
    output n4_adj_12;
    output n10;
    output n13;
    output n12;
    output n15;
    output n14;
    output n17;
    output n16;
    output n19_adj_13;
    output n18_adj_14;
    output n21_adj_15;
    output n20_adj_16;
    output n23_adj_17;
    output n22_adj_18;
    output n25_adj_19;
    output n24_adj_20;
    output n27_adj_21;
    output n26_adj_22;
    output n29_adj_23;
    output n28_adj_24;
    output n7_adj_25;
    output n31_adj_26;
    output n6_adj_27;
    output n30_adj_28;
    output n33_adj_29;
    output n32_adj_30;
    output n35_adj_31;
    output n9_adj_32;
    output n8_adj_33;
    output n34_adj_34;
    output n37_adj_35;
    output n36_adj_36;
    output n3_adj_37;
    output n2_adj_38;
    output n11_adj_39;
    output n5_adj_40;
    output n4_adj_41;
    output n7_adj_42;
    output n6_adj_43;
    output n10_adj_44;
    output n9_adj_45;
    output n8_adj_46;
    output n11_adj_47;
    output n10_adj_48;
    output n13_adj_49;
    output n12_adj_50;
    output n15_adj_51;
    output n13_adj_52;
    output n14_adj_53;
    output n17_adj_54;
    output n16_adj_55;
    output n19_adj_56;
    output n12_adj_57;
    output n18_adj_58;
    output n15_adj_59;
    output n21_adj_60;
    output [11:0]count;
    output n20_adj_61;
    output n23_adj_62;
    output n22_adj_63;
    output n25_adj_64;
    output n24_adj_65;
    output n27_adj_66;
    output n26_adj_67;
    output n29_adj_68;
    output n28_adj_69;
    output n31_adj_70;
    output n30_adj_71;
    output n9_adj_72;
    output n8_adj_73;
    output n33_adj_74;
    output n11_adj_75;
    output n10_adj_76;
    output n32_adj_77;
    output n35_adj_78;
    output n70;
    output n68;
    output n67;
    output n66;
    output n65;
    output n64;
    output n63;
    output n34_adj_79;
    output n37_adj_80;
    output n36_adj_81;
    output n13_adj_82;
    output n12_adj_83;
    output n14_adj_84;
    output n15_adj_85;
    output n17_adj_86;
    output n16_adj_87;
    output n14_adj_88;
    output n19_adj_89;
    output n18_adj_90;
    output n21_adj_91;
    output n20_adj_92;
    output n61_adj_93;
    output n23_adj_94;
    output n22_adj_95;
    output n25_adj_96;
    output n17_adj_97;
    output n16_adj_98;
    output n24_adj_99;
    output n27_adj_100;
    output n26_adj_101;
    input n76;
    input n78;
    input cout;
    input n79;
    input n81;
    input n82;
    input n84;
    input n85;
    input n87;
    input n88;
    input n90;
    input n91;
    input n93;
    input n94;
    input n96;
    input n97;
    input n99;
    input n100;
    input n102;
    input n103;
    input n105;
    input n106;
    input n108;
    input n109;
    input n111;
    input n112;
    input n114;
    input n115;
    input n117;
    input n118;
    input n120;
    output n29_adj_102;
    output n28_adj_103;
    output n2_adj_104;
    output n3_adj_105;
    output n31_adj_106;
    output n30_adj_107;
    output n33_adj_108;
    output n32_adj_109;
    output n35_adj_110;
    output n34_adj_111;
    output n37_adj_112;
    output n36_adj_113;
    output \cic_cosine_out[1] ;
    output \cic_cosine_out[0] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/top.v(61[34:43])
    
    wire n23_c;
    wire [11:0]count_11__N_1980;
    wire [71:0]comb10;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(62[99:105])
    
    wire n19866, n19865, clk_80mhz_enable_850, clk_80mhz_enable_71, 
        valid_comb;
    wire [71:0]comb10_71__N_2281;
    
    wire clk_80mhz_enable_136, clk_80mhz_enable_195, clk_80mhz_enable_341, 
        clk_80mhz_enable_394, clk_80mhz_enable_449, clk_80mhz_enable_499, 
        clk_80mhz_enable_550, clk_80mhz_enable_600, clk_80mhz_enable_652, 
        clk_80mhz_enable_702, clk_80mhz_enable_752, clk_80mhz_enable_802, 
        count_11__N_1992, n18778, n18762, n18774, n18760, n20267, 
        n14290, n18816, n18800, n18808, n18812, n19854, n19853;
    
    LUT4 i4941_2_lut (.A(n67_adj_114[11]), .B(n23_c), .Z(count_11__N_1980[11])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(92[14] 95[8])
    defparam i4941_2_lut.init = 16'hbbbb;
    LUT4 i8630_then_3_lut (.A(\cic_gain[1] ), .B(\comb10[60] ), .C(comb10[58]), 
         .Z(n19866)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i8630_then_3_lut.init = 16'he4e4;
    LUT4 i8630_else_3_lut (.A(n62), .B(\cic_gain[1] ), .C(\comb10[59] ), 
         .Z(n19865)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i8630_else_3_lut.init = 16'he2e2;
    FD1P3AX integrator_tmp_i0_i0 (.D(integrator5[0]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i0 (.D(integrator_tmp[0]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i0.GSR = "ENABLED";
    FD1S3AX integrator2_i0 (.D(integrator2_71__N_1032[0]), .CK(clk_80mhz), 
            .Q(integrator2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i0.GSR = "ENABLED";
    FD1S3AX integrator3_i0 (.D(integrator3_71__N_1104[0]), .CK(clk_80mhz), 
            .Q(integrator3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i0.GSR = "ENABLED";
    FD1S3AX integrator4_i0 (.D(integrator4_71__N_1176[0]), .CK(clk_80mhz), 
            .Q(integrator4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i0.GSR = "ENABLED";
    FD1S3AX integrator5_i0 (.D(integrator5_71__N_1248[0]), .CK(clk_80mhz), 
            .Q(integrator5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i0.GSR = "ENABLED";
    FD1P3AX comb6_i0_i0 (.D(comb6_71__N_1993[0]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(comb6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i0 (.D(comb6[0]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i0.GSR = "ENABLED";
    FD1S3AX valid_comb_63 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), .Q(valid_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63.GSR = "ENABLED";
    FD1P3AX comb7_i0_i0 (.D(comb7_71__N_2065[0]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(comb7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i0 (.D(comb7[0]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX comb8_i0_i0 (.D(comb8_71__N_2137[0]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(comb8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i0 (.D(comb8[0]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX comb9_i0_i0 (.D(comb9_71__N_2209[0]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(comb9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i0 (.D(comb9[0]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i0.GSR = "ENABLED";
    FD1S3AX integrator1_i0 (.D(integrator1_71__N_960[0]), .CK(clk_80mhz), 
            .Q(integrator1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i0.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i55_1_lut (.A(integrator_d_tmp[54]), .Z(n19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i55_1_lut.init = 16'h5555;
    FD1S3AX integrator1_i71 (.D(integrator1_71__N_960[71]), .CK(clk_80mhz), 
            .Q(integrator1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i71.GSR = "ENABLED";
    FD1S3AX integrator1_i70 (.D(integrator1_71__N_960[70]), .CK(clk_80mhz), 
            .Q(integrator1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i70.GSR = "ENABLED";
    FD1S3AX integrator1_i69 (.D(integrator1_71__N_960[69]), .CK(clk_80mhz), 
            .Q(integrator1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i69.GSR = "ENABLED";
    FD1S3AX integrator1_i68 (.D(integrator1_71__N_960[68]), .CK(clk_80mhz), 
            .Q(integrator1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i68.GSR = "ENABLED";
    FD1S3AX integrator1_i67 (.D(integrator1_71__N_960[67]), .CK(clk_80mhz), 
            .Q(integrator1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i67.GSR = "ENABLED";
    FD1S3AX integrator1_i66 (.D(integrator1_71__N_960[66]), .CK(clk_80mhz), 
            .Q(integrator1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i66.GSR = "ENABLED";
    FD1S3AX integrator1_i65 (.D(integrator1_71__N_960[65]), .CK(clk_80mhz), 
            .Q(integrator1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i65.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i56_1_lut (.A(integrator_d_tmp[55]), .Z(n18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i56_1_lut.init = 16'h5555;
    FD1S3AX integrator1_i64 (.D(integrator1_71__N_960[64]), .CK(clk_80mhz), 
            .Q(integrator1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i64.GSR = "ENABLED";
    FD1S3AX integrator1_i63 (.D(integrator1_71__N_960[63]), .CK(clk_80mhz), 
            .Q(integrator1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i63.GSR = "ENABLED";
    FD1S3AX integrator1_i62 (.D(integrator1_71__N_960[62]), .CK(clk_80mhz), 
            .Q(integrator1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i62.GSR = "ENABLED";
    FD1S3AX integrator1_i61 (.D(integrator1_71__N_960[61]), .CK(clk_80mhz), 
            .Q(integrator1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i61.GSR = "ENABLED";
    FD1S3AX integrator1_i60 (.D(integrator1_71__N_960[60]), .CK(clk_80mhz), 
            .Q(integrator1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i60.GSR = "ENABLED";
    FD1S3AX integrator1_i59 (.D(integrator1_71__N_960[59]), .CK(clk_80mhz), 
            .Q(integrator1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i59.GSR = "ENABLED";
    FD1S3AX integrator1_i58 (.D(integrator1_71__N_960[58]), .CK(clk_80mhz), 
            .Q(integrator1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i58.GSR = "ENABLED";
    FD1S3AX integrator1_i57 (.D(integrator1_71__N_960[57]), .CK(clk_80mhz), 
            .Q(integrator1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i57.GSR = "ENABLED";
    FD1S3AX integrator1_i56 (.D(integrator1_71__N_960[56]), .CK(clk_80mhz), 
            .Q(integrator1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i56.GSR = "ENABLED";
    FD1S3AX integrator1_i55 (.D(integrator1_71__N_960[55]), .CK(clk_80mhz), 
            .Q(integrator1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i55.GSR = "ENABLED";
    FD1S3AX integrator1_i54 (.D(integrator1_71__N_960[54]), .CK(clk_80mhz), 
            .Q(integrator1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i54.GSR = "ENABLED";
    FD1S3AX integrator1_i53 (.D(integrator1_71__N_960[53]), .CK(clk_80mhz), 
            .Q(integrator1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i53.GSR = "ENABLED";
    FD1S3AX integrator1_i52 (.D(integrator1_71__N_960[52]), .CK(clk_80mhz), 
            .Q(integrator1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i52.GSR = "ENABLED";
    FD1S3AX integrator1_i51 (.D(integrator1_71__N_960[51]), .CK(clk_80mhz), 
            .Q(integrator1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i51.GSR = "ENABLED";
    FD1S3AX integrator1_i50 (.D(integrator1_71__N_960[50]), .CK(clk_80mhz), 
            .Q(integrator1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i50.GSR = "ENABLED";
    FD1S3AX integrator1_i49 (.D(integrator1_71__N_960[49]), .CK(clk_80mhz), 
            .Q(integrator1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i49.GSR = "ENABLED";
    FD1S3AX integrator1_i48 (.D(integrator1_71__N_960[48]), .CK(clk_80mhz), 
            .Q(integrator1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i48.GSR = "ENABLED";
    FD1S3AX integrator1_i47 (.D(integrator1_71__N_960[47]), .CK(clk_80mhz), 
            .Q(integrator1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i47.GSR = "ENABLED";
    FD1S3AX integrator1_i46 (.D(integrator1_71__N_960[46]), .CK(clk_80mhz), 
            .Q(integrator1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i46.GSR = "ENABLED";
    FD1S3AX integrator1_i45 (.D(integrator1_71__N_960[45]), .CK(clk_80mhz), 
            .Q(integrator1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i45.GSR = "ENABLED";
    FD1S3AX integrator1_i44 (.D(integrator1_71__N_960[44]), .CK(clk_80mhz), 
            .Q(integrator1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i44.GSR = "ENABLED";
    FD1S3AX integrator1_i43 (.D(integrator1_71__N_960[43]), .CK(clk_80mhz), 
            .Q(integrator1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i43.GSR = "ENABLED";
    FD1S3AX integrator1_i42 (.D(integrator1_71__N_960[42]), .CK(clk_80mhz), 
            .Q(integrator1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i42.GSR = "ENABLED";
    FD1S3AX integrator1_i41 (.D(integrator1_71__N_960[41]), .CK(clk_80mhz), 
            .Q(integrator1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i41.GSR = "ENABLED";
    FD1S3AX integrator1_i40 (.D(integrator1_71__N_960[40]), .CK(clk_80mhz), 
            .Q(integrator1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i40.GSR = "ENABLED";
    FD1S3AX integrator1_i39 (.D(integrator1_71__N_960[39]), .CK(clk_80mhz), 
            .Q(integrator1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i39.GSR = "ENABLED";
    FD1S3AX integrator1_i38 (.D(integrator1_71__N_960[38]), .CK(clk_80mhz), 
            .Q(integrator1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i38.GSR = "ENABLED";
    FD1S3AX integrator1_i37 (.D(integrator1_71__N_960[37]), .CK(clk_80mhz), 
            .Q(integrator1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i37.GSR = "ENABLED";
    FD1S3AX integrator1_i36 (.D(integrator1_71__N_960[36]), .CK(clk_80mhz), 
            .Q(integrator1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i36.GSR = "ENABLED";
    FD1S3AX integrator1_i35 (.D(integrator1_71__N_960[35]), .CK(clk_80mhz), 
            .Q(integrator1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i35.GSR = "ENABLED";
    FD1S3AX integrator1_i34 (.D(integrator1_71__N_960[34]), .CK(clk_80mhz), 
            .Q(integrator1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i34.GSR = "ENABLED";
    FD1S3AX integrator1_i33 (.D(integrator1_71__N_960[33]), .CK(clk_80mhz), 
            .Q(integrator1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i33.GSR = "ENABLED";
    FD1S3AX integrator1_i32 (.D(integrator1_71__N_960[32]), .CK(clk_80mhz), 
            .Q(integrator1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i32.GSR = "ENABLED";
    FD1S3AX integrator1_i31 (.D(integrator1_71__N_960[31]), .CK(clk_80mhz), 
            .Q(integrator1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i31.GSR = "ENABLED";
    FD1S3AX integrator1_i30 (.D(integrator1_71__N_960[30]), .CK(clk_80mhz), 
            .Q(integrator1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i30.GSR = "ENABLED";
    FD1S3AX integrator1_i29 (.D(integrator1_71__N_960[29]), .CK(clk_80mhz), 
            .Q(integrator1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i29.GSR = "ENABLED";
    FD1S3AX integrator1_i28 (.D(integrator1_71__N_960[28]), .CK(clk_80mhz), 
            .Q(integrator1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i28.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i53_1_lut (.A(integrator_d_tmp[52]), .Z(n21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i53_1_lut.init = 16'h5555;
    FD1S3AX integrator1_i27 (.D(integrator1_71__N_960[27]), .CK(clk_80mhz), 
            .Q(integrator1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i27.GSR = "ENABLED";
    FD1S3AX integrator1_i26 (.D(integrator1_71__N_960[26]), .CK(clk_80mhz), 
            .Q(integrator1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i26.GSR = "ENABLED";
    FD1S3AX integrator1_i25 (.D(integrator1_71__N_960[25]), .CK(clk_80mhz), 
            .Q(integrator1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i25.GSR = "ENABLED";
    FD1S3AX integrator1_i24 (.D(integrator1_71__N_960[24]), .CK(clk_80mhz), 
            .Q(integrator1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i24.GSR = "ENABLED";
    FD1S3AX integrator1_i23 (.D(integrator1_71__N_960[23]), .CK(clk_80mhz), 
            .Q(integrator1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i23.GSR = "ENABLED";
    FD1S3AX integrator1_i22 (.D(integrator1_71__N_960[22]), .CK(clk_80mhz), 
            .Q(integrator1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i22.GSR = "ENABLED";
    FD1S3AX integrator1_i21 (.D(integrator1_71__N_960[21]), .CK(clk_80mhz), 
            .Q(integrator1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i21.GSR = "ENABLED";
    FD1S3AX integrator1_i20 (.D(integrator1_71__N_960[20]), .CK(clk_80mhz), 
            .Q(integrator1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i20.GSR = "ENABLED";
    FD1S3AX integrator1_i19 (.D(integrator1_71__N_960[19]), .CK(clk_80mhz), 
            .Q(integrator1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i19.GSR = "ENABLED";
    FD1S3AX integrator1_i18 (.D(integrator1_71__N_960[18]), .CK(clk_80mhz), 
            .Q(integrator1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i18.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i54_1_lut (.A(integrator_d_tmp[53]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i54_1_lut.init = 16'h5555;
    FD1S3AX integrator1_i17 (.D(integrator1_71__N_960[17]), .CK(clk_80mhz), 
            .Q(integrator1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i17.GSR = "ENABLED";
    FD1S3AX integrator1_i16 (.D(integrator1_71__N_960[16]), .CK(clk_80mhz), 
            .Q(integrator1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i16.GSR = "ENABLED";
    FD1S3AX integrator1_i15 (.D(integrator1_71__N_960[15]), .CK(clk_80mhz), 
            .Q(integrator1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i15.GSR = "ENABLED";
    FD1S3AX integrator1_i14 (.D(integrator1_71__N_960[14]), .CK(clk_80mhz), 
            .Q(integrator1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i14.GSR = "ENABLED";
    FD1S3AX integrator1_i13 (.D(integrator1_71__N_960[13]), .CK(clk_80mhz), 
            .Q(integrator1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i13.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i51_1_lut (.A(integrator_d_tmp[50]), .Z(n23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i52_1_lut (.A(integrator_d_tmp[51]), .Z(n22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i49_1_lut (.A(integrator_d_tmp[48]), .Z(n25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i50_1_lut (.A(integrator_d_tmp[49]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i47_1_lut (.A(integrator_d_tmp[46]), .Z(n27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i71_1_lut (.A(comb_d8[70]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i72_1_lut (.A(comb_d8[71]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i48_1_lut (.A(integrator_d_tmp[47]), .Z(n26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i69_1_lut (.A(comb_d8[68]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i45_1_lut (.A(integrator_d_tmp[44]), .Z(n29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i46_1_lut (.A(integrator_d_tmp[45]), .Z(n28_adj_1)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i46_1_lut.init = 16'h5555;
    FD1S3AX integrator1_i12 (.D(integrator1_71__N_960[12]), .CK(clk_80mhz), 
            .Q(integrator1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i12.GSR = "ENABLED";
    FD1S3AX integrator1_i11 (.D(integrator1_71__N_960[11]), .CK(clk_80mhz), 
            .Q(integrator1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i11.GSR = "ENABLED";
    FD1S3AX integrator1_i10 (.D(integrator1_71__N_960[10]), .CK(clk_80mhz), 
            .Q(integrator1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i10.GSR = "ENABLED";
    FD1S3AX integrator1_i9 (.D(integrator1_71__N_960[9]), .CK(clk_80mhz), 
            .Q(integrator1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i9.GSR = "ENABLED";
    FD1S3AX integrator1_i8 (.D(integrator1_71__N_960[8]), .CK(clk_80mhz), 
            .Q(integrator1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i8.GSR = "ENABLED";
    FD1S3AX integrator1_i7 (.D(integrator1_71__N_960[7]), .CK(clk_80mhz), 
            .Q(integrator1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i7.GSR = "ENABLED";
    FD1S3AX integrator1_i6 (.D(integrator1_71__N_960[6]), .CK(clk_80mhz), 
            .Q(integrator1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i6.GSR = "ENABLED";
    FD1S3AX integrator1_i5 (.D(integrator1_71__N_960[5]), .CK(clk_80mhz), 
            .Q(integrator1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i5.GSR = "ENABLED";
    FD1S3AX integrator1_i4 (.D(integrator1_71__N_960[4]), .CK(clk_80mhz), 
            .Q(integrator1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i4.GSR = "ENABLED";
    FD1S3AX integrator1_i3 (.D(integrator1_71__N_960[3]), .CK(clk_80mhz), 
            .Q(integrator1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i3.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i43_1_lut (.A(integrator_d_tmp[42]), .Z(n31_adj_2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i43_1_lut.init = 16'h5555;
    FD1S3AX integrator1_i2 (.D(integrator1_71__N_960[2]), .CK(clk_80mhz), 
            .Q(integrator1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i2.GSR = "ENABLED";
    FD1S3AX integrator1_i1 (.D(integrator1_71__N_960[1]), .CK(clk_80mhz), 
            .Q(integrator1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator1_i1.GSR = "ENABLED";
    FD1P3AX comb10__i16 (.D(comb10_71__N_2281[71]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[71] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i16.GSR = "ENABLED";
    FD1P3AX comb10__i15 (.D(comb10_71__N_2281[70]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[70] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i15.GSR = "ENABLED";
    FD1P3AX comb10__i14 (.D(comb10_71__N_2281[69]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[69] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i14.GSR = "ENABLED";
    FD1P3AX comb10__i13 (.D(comb10_71__N_2281[68]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[68] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i13.GSR = "ENABLED";
    FD1P3AX comb10__i12 (.D(comb10_71__N_2281[67]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[67] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i12.GSR = "ENABLED";
    FD1P3AX comb10__i11 (.D(comb10_71__N_2281[66]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[66] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i11.GSR = "ENABLED";
    FD1P3AX comb10__i10 (.D(comb10_71__N_2281[65]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[65] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i10.GSR = "ENABLED";
    FD1P3AX comb10__i9 (.D(comb10_71__N_2281[64]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[64] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i9.GSR = "ENABLED";
    FD1P3AX comb10__i8 (.D(comb10_71__N_2281[63]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[63] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i8.GSR = "ENABLED";
    FD1P3AX comb10__i7 (.D(comb10_71__N_2281[62]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[62] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i7.GSR = "ENABLED";
    FD1P3AX comb10__i6 (.D(comb10_71__N_2281[61]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[61] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i6.GSR = "ENABLED";
    FD1P3AX comb10__i5 (.D(comb10_71__N_2281[60]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i5.GSR = "ENABLED";
    FD1P3AX comb10__i4 (.D(comb10_71__N_2281[59]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(\comb10[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i4.GSR = "ENABLED";
    FD1P3AX comb10__i3 (.D(comb10_71__N_2281[58]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(comb10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i3.GSR = "ENABLED";
    FD1P3AX comb10__i2 (.D(comb10_71__N_2281[57]), .SP(clk_80mhz_enable_71), 
            .CK(clk_80mhz), .Q(comb10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb10__i2.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i71 (.D(comb9[71]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i71.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i44_1_lut (.A(integrator_d_tmp[43]), .Z(n30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i44_1_lut.init = 16'h5555;
    FD1P3AX comb_d9_i0_i70 (.D(comb9[70]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i69 (.D(comb9[69]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i68 (.D(comb9[68]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i67 (.D(comb9[67]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i66 (.D(comb9[66]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i65 (.D(comb9[65]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i64 (.D(comb9[64]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i63 (.D(comb9[63]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i62 (.D(comb9[62]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i61 (.D(comb9[61]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i60 (.D(comb9[60]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i59 (.D(comb9[59]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i58 (.D(comb9[58]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i57 (.D(comb9[57]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i56 (.D(comb9[56]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i55 (.D(comb9[55]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i54 (.D(comb9[54]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i53 (.D(comb9[53]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i52 (.D(comb9[52]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i51 (.D(comb9[51]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i51.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i41_1_lut (.A(integrator_d_tmp[40]), .Z(n33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i41_1_lut.init = 16'h5555;
    FD1P3AX comb_d9_i0_i50 (.D(comb9[50]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i50.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i42_1_lut (.A(integrator_d_tmp[41]), .Z(n32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i42_1_lut.init = 16'h5555;
    FD1P3AX comb_d9_i0_i49 (.D(comb9[49]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i48 (.D(comb9[48]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i47 (.D(comb9[47]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i46 (.D(comb9[46]), .SP(clk_80mhz_enable_71), .CK(clk_80mhz), 
            .Q(comb_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i46.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i39_1_lut (.A(integrator_d_tmp[38]), .Z(n35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i39_1_lut.init = 16'h5555;
    FD1P3AX comb_d9_i0_i45 (.D(comb9[45]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i45.GSR = "ENABLED";
    LUT4 sub_29_inv_0_i70_1_lut (.A(comb_d8[69]), .Z(n4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i70_1_lut.init = 16'h5555;
    FD1P3AX comb_d9_i0_i44 (.D(comb9[44]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i43 (.D(comb9[43]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i42 (.D(comb9[42]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i41 (.D(comb9[41]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i40 (.D(comb9[40]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i40.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i40_1_lut (.A(integrator_d_tmp[39]), .Z(n34_adj_3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i37_1_lut (.A(integrator_d_tmp[36]), .Z(n37_adj_4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i37_1_lut.init = 16'h5555;
    FD1P3AX comb_d9_i0_i39 (.D(comb9[39]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i38 (.D(comb9[38]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i37 (.D(comb9[37]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i36 (.D(comb9[36]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i35 (.D(comb9[35]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i34 (.D(comb9[34]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i33 (.D(comb9[33]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i32 (.D(comb9[32]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i31 (.D(comb9[31]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i30 (.D(comb9[30]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i29 (.D(comb9[29]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i28 (.D(comb9[28]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i27 (.D(comb9[27]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i26 (.D(comb9[26]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i25 (.D(comb9[25]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i24 (.D(comb9[24]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i23 (.D(comb9[23]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i22 (.D(comb9[22]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i21 (.D(comb9[21]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i20 (.D(comb9[20]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i19 (.D(comb9[19]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i18 (.D(comb9[18]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i18.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i38_1_lut (.A(integrator_d_tmp[37]), .Z(n36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i38_1_lut.init = 16'h5555;
    FD1P3AX comb_d9_i0_i17 (.D(comb9[17]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i17.GSR = "ENABLED";
    LUT4 sub_29_inv_0_i67_1_lut (.A(comb_d8[66]), .Z(n7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i67_1_lut.init = 16'h5555;
    FD1P3AX comb_d9_i0_i16 (.D(comb9[16]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i16.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i71_1_lut (.A(comb_d6[70]), .Z(n3_adj_5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i71_1_lut.init = 16'h5555;
    FD1P3AX comb_d9_i0_i15 (.D(comb9[15]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i15.GSR = "ENABLED";
    LUT4 sub_29_inv_0_i68_1_lut (.A(comb_d8[67]), .Z(n6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i68_1_lut.init = 16'h5555;
    FD1P3AX comb_d9_i0_i14 (.D(comb9[14]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i13 (.D(comb9[13]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i12 (.D(comb9[12]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i12.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i72_1_lut (.A(comb_d6[71]), .Z(n2_adj_6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i72_1_lut.init = 16'h5555;
    FD1P3AX comb_d9_i0_i11 (.D(comb9[11]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i11.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i69_1_lut (.A(comb_d6[68]), .Z(n5_adj_7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i69_1_lut.init = 16'h5555;
    FD1P3AX comb_d9_i0_i10 (.D(comb9[10]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i9 (.D(comb9[9]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i8 (.D(comb9[8]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i7 (.D(comb9[7]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i6 (.D(comb9[6]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i5 (.D(comb9[5]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i4 (.D(comb9[4]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i3 (.D(comb9[3]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i2 (.D(comb9[2]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i1 (.D(comb9[1]), .SP(clk_80mhz_enable_136), .CK(clk_80mhz), 
            .Q(comb_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX comb9_i0_i71 (.D(comb9_71__N_2209[71]), .SP(clk_80mhz_enable_136), 
            .CK(clk_80mhz), .Q(comb9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i71.GSR = "ENABLED";
    FD1P3AX comb9_i0_i70 (.D(comb9_71__N_2209[70]), .SP(clk_80mhz_enable_136), 
            .CK(clk_80mhz), .Q(comb9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i70.GSR = "ENABLED";
    FD1P3AX comb9_i0_i69 (.D(comb9_71__N_2209[69]), .SP(clk_80mhz_enable_136), 
            .CK(clk_80mhz), .Q(comb9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i69.GSR = "ENABLED";
    FD1P3AX comb9_i0_i68 (.D(comb9_71__N_2209[68]), .SP(clk_80mhz_enable_136), 
            .CK(clk_80mhz), .Q(comb9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i68.GSR = "ENABLED";
    FD1P3AX comb9_i0_i67 (.D(comb9_71__N_2209[67]), .SP(clk_80mhz_enable_136), 
            .CK(clk_80mhz), .Q(comb9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i67.GSR = "ENABLED";
    FD1P3AX comb9_i0_i66 (.D(comb9_71__N_2209[66]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i66.GSR = "ENABLED";
    FD1P3AX comb9_i0_i65 (.D(comb9_71__N_2209[65]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i65.GSR = "ENABLED";
    FD1P3AX comb9_i0_i64 (.D(comb9_71__N_2209[64]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i64.GSR = "ENABLED";
    FD1P3AX comb9_i0_i63 (.D(comb9_71__N_2209[63]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i63.GSR = "ENABLED";
    FD1P3AX comb9_i0_i62 (.D(comb9_71__N_2209[62]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i62.GSR = "ENABLED";
    FD1P3AX comb9_i0_i61 (.D(comb9_71__N_2209[61]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i61.GSR = "ENABLED";
    FD1P3AX comb9_i0_i60 (.D(comb9_71__N_2209[60]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i60.GSR = "ENABLED";
    FD1P3AX comb9_i0_i59 (.D(comb9_71__N_2209[59]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i59.GSR = "ENABLED";
    FD1P3AX comb9_i0_i58 (.D(comb9_71__N_2209[58]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i58.GSR = "ENABLED";
    FD1P3AX comb9_i0_i57 (.D(comb9_71__N_2209[57]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i57.GSR = "ENABLED";
    FD1P3AX comb9_i0_i56 (.D(comb9_71__N_2209[56]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i56.GSR = "ENABLED";
    FD1P3AX comb9_i0_i55 (.D(comb9_71__N_2209[55]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i55.GSR = "ENABLED";
    FD1P3AX comb9_i0_i54 (.D(comb9_71__N_2209[54]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i54.GSR = "ENABLED";
    FD1P3AX comb9_i0_i53 (.D(comb9_71__N_2209[53]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i53.GSR = "ENABLED";
    FD1P3AX comb9_i0_i52 (.D(comb9_71__N_2209[52]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i52.GSR = "ENABLED";
    FD1P3AX comb9_i0_i51 (.D(comb9_71__N_2209[51]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i51.GSR = "ENABLED";
    FD1P3AX comb9_i0_i50 (.D(comb9_71__N_2209[50]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i50.GSR = "ENABLED";
    FD1P3AX comb9_i0_i49 (.D(comb9_71__N_2209[49]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i49.GSR = "ENABLED";
    FD1P3AX comb9_i0_i48 (.D(comb9_71__N_2209[48]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i48.GSR = "ENABLED";
    FD1P3AX comb9_i0_i47 (.D(comb9_71__N_2209[47]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i47.GSR = "ENABLED";
    FD1P3AX comb9_i0_i46 (.D(comb9_71__N_2209[46]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i46.GSR = "ENABLED";
    FD1P3AX comb9_i0_i45 (.D(comb9_71__N_2209[45]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i45.GSR = "ENABLED";
    FD1P3AX comb9_i0_i44 (.D(comb9_71__N_2209[44]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i44.GSR = "ENABLED";
    FD1P3AX comb9_i0_i43 (.D(comb9_71__N_2209[43]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i43.GSR = "ENABLED";
    FD1P3AX comb9_i0_i42 (.D(comb9_71__N_2209[42]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i42.GSR = "ENABLED";
    FD1P3AX comb9_i0_i41 (.D(comb9_71__N_2209[41]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i41.GSR = "ENABLED";
    FD1P3AX comb9_i0_i40 (.D(comb9_71__N_2209[40]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i40.GSR = "ENABLED";
    FD1P3AX comb9_i0_i39 (.D(comb9_71__N_2209[39]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i39.GSR = "ENABLED";
    FD1P3AX comb9_i0_i38 (.D(comb9_71__N_2209[38]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i38.GSR = "ENABLED";
    FD1P3AX comb9_i0_i37 (.D(comb9_71__N_2209[37]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i37.GSR = "ENABLED";
    FD1P3AX comb9_i0_i36 (.D(comb9_71__N_2209[36]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i36.GSR = "ENABLED";
    FD1P3AX comb9_i0_i35 (.D(comb9_71__N_2209[35]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i35.GSR = "ENABLED";
    FD1P3AX comb9_i0_i34 (.D(comb9_71__N_2209[34]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i34.GSR = "ENABLED";
    FD1P3AX comb9_i0_i33 (.D(comb9_71__N_2209[33]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i33.GSR = "ENABLED";
    FD1P3AX comb9_i0_i32 (.D(comb9_71__N_2209[32]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i32.GSR = "ENABLED";
    FD1P3AX comb9_i0_i31 (.D(comb9_71__N_2209[31]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i31.GSR = "ENABLED";
    FD1P3AX comb9_i0_i30 (.D(comb9_71__N_2209[30]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i30.GSR = "ENABLED";
    FD1P3AX comb9_i0_i29 (.D(comb9_71__N_2209[29]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i29.GSR = "ENABLED";
    FD1P3AX comb9_i0_i28 (.D(comb9_71__N_2209[28]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i28.GSR = "ENABLED";
    FD1P3AX comb9_i0_i27 (.D(comb9_71__N_2209[27]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i27.GSR = "ENABLED";
    FD1P3AX comb9_i0_i26 (.D(comb9_71__N_2209[26]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i26.GSR = "ENABLED";
    FD1P3AX comb9_i0_i25 (.D(comb9_71__N_2209[25]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i25.GSR = "ENABLED";
    FD1P3AX comb9_i0_i24 (.D(comb9_71__N_2209[24]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i24.GSR = "ENABLED";
    FD1P3AX comb9_i0_i23 (.D(comb9_71__N_2209[23]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i23.GSR = "ENABLED";
    FD1P3AX comb9_i0_i22 (.D(comb9_71__N_2209[22]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i22.GSR = "ENABLED";
    FD1P3AX comb9_i0_i21 (.D(comb9_71__N_2209[21]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i21.GSR = "ENABLED";
    FD1P3AX comb9_i0_i20 (.D(comb9_71__N_2209[20]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i20.GSR = "ENABLED";
    FD1P3AX comb9_i0_i19 (.D(comb9_71__N_2209[19]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i19.GSR = "ENABLED";
    FD1P3AX comb9_i0_i18 (.D(comb9_71__N_2209[18]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i18.GSR = "ENABLED";
    FD1P3AX comb9_i0_i17 (.D(comb9_71__N_2209[17]), .SP(clk_80mhz_enable_195), 
            .CK(clk_80mhz), .Q(comb9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i17.GSR = "ENABLED";
    FD1P3AX comb9_i0_i16 (.D(comb9_71__N_2209[16]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i16.GSR = "ENABLED";
    FD1P3AX comb9_i0_i15 (.D(comb9_71__N_2209[15]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i15.GSR = "ENABLED";
    FD1P3AX comb9_i0_i14 (.D(comb9_71__N_2209[14]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i14.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i70_1_lut (.A(comb_d6[69]), .Z(n4_adj_8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i67_1_lut (.A(comb_d6[66]), .Z(n7_adj_9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i68_1_lut (.A(comb_d6[67]), .Z(n6_adj_10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i65_1_lut (.A(comb_d6[64]), .Z(n9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i65_1_lut.init = 16'h5555;
    FD1P3AX comb9_i0_i13 (.D(comb9_71__N_2209[13]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i13.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i66_1_lut (.A(comb_d6[65]), .Z(n8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i69_1_lut (.A(integrator_d_tmp[68]), .Z(n5_adj_11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i69_1_lut.init = 16'h5555;
    FD1P3AX comb9_i0_i12 (.D(comb9_71__N_2209[12]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i12.GSR = "ENABLED";
    FD1P3AX comb9_i0_i11 (.D(comb9_71__N_2209[11]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i11.GSR = "ENABLED";
    FD1P3AX comb9_i0_i10 (.D(comb9_71__N_2209[10]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i10.GSR = "ENABLED";
    FD1P3AX comb9_i0_i9 (.D(comb9_71__N_2209[9]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i9.GSR = "ENABLED";
    FD1P3AX comb9_i0_i8 (.D(comb9_71__N_2209[8]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i8.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i63_1_lut (.A(comb_d6[62]), .Z(n11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i63_1_lut.init = 16'h5555;
    FD1P3AX comb9_i0_i7 (.D(comb9_71__N_2209[7]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i7.GSR = "ENABLED";
    FD1P3AX comb9_i0_i6 (.D(comb9_71__N_2209[6]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i6.GSR = "ENABLED";
    FD1P3AX comb9_i0_i5 (.D(comb9_71__N_2209[5]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i5.GSR = "ENABLED";
    FD1P3AX comb9_i0_i4 (.D(comb9_71__N_2209[4]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i4.GSR = "ENABLED";
    FD1P3AX comb9_i0_i3 (.D(comb9_71__N_2209[3]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i3.GSR = "ENABLED";
    FD1P3AX comb9_i0_i2 (.D(comb9_71__N_2209[2]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i2.GSR = "ENABLED";
    FD1P3AX comb9_i0_i1 (.D(comb9_71__N_2209[1]), .SP(clk_80mhz_enable_341), 
            .CK(clk_80mhz), .Q(comb9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb9_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i71 (.D(comb8[71]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i70 (.D(comb8[70]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i69 (.D(comb8[69]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i68 (.D(comb8[68]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i67 (.D(comb8[67]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i66 (.D(comb8[66]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i65 (.D(comb8[65]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i64 (.D(comb8[64]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i63 (.D(comb8[63]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i62 (.D(comb8[62]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i61 (.D(comb8[61]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i60 (.D(comb8[60]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i59 (.D(comb8[59]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i58 (.D(comb8[58]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i57 (.D(comb8[57]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i56 (.D(comb8[56]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i55 (.D(comb8[55]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i54 (.D(comb8[54]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i53 (.D(comb8[53]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i52 (.D(comb8[52]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i51 (.D(comb8[51]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i50 (.D(comb8[50]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i49 (.D(comb8[49]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i48 (.D(comb8[48]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i47 (.D(comb8[47]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i46 (.D(comb8[46]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i45 (.D(comb8[45]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i44 (.D(comb8[44]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i43 (.D(comb8[43]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i42 (.D(comb8[42]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i41 (.D(comb8[41]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i40 (.D(comb8[40]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i39 (.D(comb8[39]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i38 (.D(comb8[38]), .SP(clk_80mhz_enable_341), .CK(clk_80mhz), 
            .Q(comb_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i38.GSR = "ENABLED";
    LUT4 comb10_71__I_0_77_i62_3_lut (.A(\comb10[61] ), .B(\comb10[62] ), 
         .C(\cic_gain[0] ), .Z(n62)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i62_3_lut.init = 16'hcaca;
    FD1P3AX comb_d8_i0_i37 (.D(comb8[37]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i36 (.D(comb8[36]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i35 (.D(comb8[35]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i34 (.D(comb8[34]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i33 (.D(comb8[33]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i32 (.D(comb8[32]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i31 (.D(comb8[31]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i30 (.D(comb8[30]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i29 (.D(comb8[29]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i28 (.D(comb8[28]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i27 (.D(comb8[27]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i26 (.D(comb8[26]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i25 (.D(comb8[25]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i24 (.D(comb8[24]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i23 (.D(comb8[23]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i22 (.D(comb8[22]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i21 (.D(comb8[21]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i20 (.D(comb8[20]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i19 (.D(comb8[19]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i18 (.D(comb8[18]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i17 (.D(comb8[17]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i16 (.D(comb8[16]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i15 (.D(comb8[15]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i14 (.D(comb8[14]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i13 (.D(comb8[13]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i12 (.D(comb8[12]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i11 (.D(comb8[11]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i10 (.D(comb8[10]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i9 (.D(comb8[9]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i8 (.D(comb8[8]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i7 (.D(comb8[7]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i6 (.D(comb8[6]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i5 (.D(comb8[5]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i4 (.D(comb8[4]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i3 (.D(comb8[3]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i2 (.D(comb8[2]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i1 (.D(comb8[1]), .SP(clk_80mhz_enable_394), .CK(clk_80mhz), 
            .Q(comb_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX comb8_i0_i71 (.D(comb8_71__N_2137[71]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i71.GSR = "ENABLED";
    FD1P3AX comb8_i0_i70 (.D(comb8_71__N_2137[70]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i70.GSR = "ENABLED";
    FD1P3AX comb8_i0_i69 (.D(comb8_71__N_2137[69]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i69.GSR = "ENABLED";
    FD1P3AX comb8_i0_i68 (.D(comb8_71__N_2137[68]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i68.GSR = "ENABLED";
    FD1P3AX comb8_i0_i67 (.D(comb8_71__N_2137[67]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i67.GSR = "ENABLED";
    FD1P3AX comb8_i0_i66 (.D(comb8_71__N_2137[66]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i66.GSR = "ENABLED";
    FD1P3AX comb8_i0_i65 (.D(comb8_71__N_2137[65]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i65.GSR = "ENABLED";
    FD1P3AX comb8_i0_i64 (.D(comb8_71__N_2137[64]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i64.GSR = "ENABLED";
    FD1P3AX comb8_i0_i63 (.D(comb8_71__N_2137[63]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i63.GSR = "ENABLED";
    FD1P3AX comb8_i0_i62 (.D(comb8_71__N_2137[62]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i62.GSR = "ENABLED";
    FD1P3AX comb8_i0_i61 (.D(comb8_71__N_2137[61]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i61.GSR = "ENABLED";
    FD1P3AX comb8_i0_i60 (.D(comb8_71__N_2137[60]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i60.GSR = "ENABLED";
    FD1P3AX comb8_i0_i59 (.D(comb8_71__N_2137[59]), .SP(clk_80mhz_enable_394), 
            .CK(clk_80mhz), .Q(comb8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i59.GSR = "ENABLED";
    FD1P3AX comb8_i0_i58 (.D(comb8_71__N_2137[58]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i58.GSR = "ENABLED";
    FD1P3AX comb8_i0_i57 (.D(comb8_71__N_2137[57]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i57.GSR = "ENABLED";
    FD1P3AX comb8_i0_i56 (.D(comb8_71__N_2137[56]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i56.GSR = "ENABLED";
    FD1P3AX comb8_i0_i55 (.D(comb8_71__N_2137[55]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i55.GSR = "ENABLED";
    FD1P3AX comb8_i0_i54 (.D(comb8_71__N_2137[54]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i54.GSR = "ENABLED";
    FD1P3AX comb8_i0_i53 (.D(comb8_71__N_2137[53]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i53.GSR = "ENABLED";
    FD1P3AX comb8_i0_i52 (.D(comb8_71__N_2137[52]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i52.GSR = "ENABLED";
    FD1P3AX comb8_i0_i51 (.D(comb8_71__N_2137[51]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i51.GSR = "ENABLED";
    FD1P3AX comb8_i0_i50 (.D(comb8_71__N_2137[50]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i50.GSR = "ENABLED";
    FD1P3AX comb8_i0_i49 (.D(comb8_71__N_2137[49]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i49.GSR = "ENABLED";
    FD1P3AX comb8_i0_i48 (.D(comb8_71__N_2137[48]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i48.GSR = "ENABLED";
    FD1P3AX comb8_i0_i47 (.D(comb8_71__N_2137[47]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i47.GSR = "ENABLED";
    FD1P3AX comb8_i0_i46 (.D(comb8_71__N_2137[46]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i46.GSR = "ENABLED";
    FD1P3AX comb8_i0_i45 (.D(comb8_71__N_2137[45]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i45.GSR = "ENABLED";
    FD1P3AX comb8_i0_i44 (.D(comb8_71__N_2137[44]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i44.GSR = "ENABLED";
    FD1P3AX comb8_i0_i43 (.D(comb8_71__N_2137[43]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i43.GSR = "ENABLED";
    FD1P3AX comb8_i0_i42 (.D(comb8_71__N_2137[42]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i42.GSR = "ENABLED";
    FD1P3AX comb8_i0_i41 (.D(comb8_71__N_2137[41]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i41.GSR = "ENABLED";
    FD1P3AX comb8_i0_i40 (.D(comb8_71__N_2137[40]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i40.GSR = "ENABLED";
    FD1P3AX comb8_i0_i39 (.D(comb8_71__N_2137[39]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i39.GSR = "ENABLED";
    FD1P3AX comb8_i0_i38 (.D(comb8_71__N_2137[38]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i38.GSR = "ENABLED";
    FD1P3AX comb8_i0_i37 (.D(comb8_71__N_2137[37]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i37.GSR = "ENABLED";
    FD1P3AX comb8_i0_i36 (.D(comb8_71__N_2137[36]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i36.GSR = "ENABLED";
    FD1P3AX comb8_i0_i35 (.D(comb8_71__N_2137[35]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i35.GSR = "ENABLED";
    FD1P3AX comb8_i0_i34 (.D(comb8_71__N_2137[34]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i34.GSR = "ENABLED";
    FD1P3AX comb8_i0_i33 (.D(comb8_71__N_2137[33]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i33.GSR = "ENABLED";
    FD1P3AX comb8_i0_i32 (.D(comb8_71__N_2137[32]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i32.GSR = "ENABLED";
    FD1P3AX comb8_i0_i31 (.D(comb8_71__N_2137[31]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i31.GSR = "ENABLED";
    FD1P3AX comb8_i0_i30 (.D(comb8_71__N_2137[30]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i30.GSR = "ENABLED";
    FD1P3AX comb8_i0_i29 (.D(comb8_71__N_2137[29]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i29.GSR = "ENABLED";
    FD1P3AX comb8_i0_i28 (.D(comb8_71__N_2137[28]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i28.GSR = "ENABLED";
    FD1P3AX comb8_i0_i27 (.D(comb8_71__N_2137[27]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i27.GSR = "ENABLED";
    FD1P3AX comb8_i0_i26 (.D(comb8_71__N_2137[26]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i26.GSR = "ENABLED";
    FD1P3AX comb8_i0_i25 (.D(comb8_71__N_2137[25]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i25.GSR = "ENABLED";
    FD1P3AX comb8_i0_i24 (.D(comb8_71__N_2137[24]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i24.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i70_1_lut (.A(integrator_d_tmp[69]), .Z(n4_adj_12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i70_1_lut.init = 16'h5555;
    FD1P3AX comb8_i0_i23 (.D(comb8_71__N_2137[23]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i23.GSR = "ENABLED";
    FD1P3AX comb8_i0_i22 (.D(comb8_71__N_2137[22]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i22.GSR = "ENABLED";
    FD1P3AX comb8_i0_i21 (.D(comb8_71__N_2137[21]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i21.GSR = "ENABLED";
    FD1P3AX comb8_i0_i20 (.D(comb8_71__N_2137[20]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i20.GSR = "ENABLED";
    FD1P3AX comb8_i0_i19 (.D(comb8_71__N_2137[19]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i19.GSR = "ENABLED";
    FD1P3AX comb8_i0_i18 (.D(comb8_71__N_2137[18]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i18.GSR = "ENABLED";
    FD1P3AX comb8_i0_i17 (.D(comb8_71__N_2137[17]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i17.GSR = "ENABLED";
    FD1P3AX comb8_i0_i16 (.D(comb8_71__N_2137[16]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i16.GSR = "ENABLED";
    FD1P3AX comb8_i0_i15 (.D(comb8_71__N_2137[15]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i15.GSR = "ENABLED";
    FD1P3AX comb8_i0_i14 (.D(comb8_71__N_2137[14]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i14.GSR = "ENABLED";
    FD1P3AX comb8_i0_i13 (.D(comb8_71__N_2137[13]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i13.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i64_1_lut (.A(comb_d6[63]), .Z(n10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i61_1_lut (.A(comb_d6[60]), .Z(n13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i61_1_lut.init = 16'h5555;
    FD1P3AX comb8_i0_i12 (.D(comb8_71__N_2137[12]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i12.GSR = "ENABLED";
    FD1P3AX comb8_i0_i11 (.D(comb8_71__N_2137[11]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i11.GSR = "ENABLED";
    FD1P3AX comb8_i0_i10 (.D(comb8_71__N_2137[10]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i10.GSR = "ENABLED";
    FD1P3AX comb8_i0_i9 (.D(comb8_71__N_2137[9]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(comb8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i9.GSR = "ENABLED";
    FD1P3AX comb8_i0_i8 (.D(comb8_71__N_2137[8]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(comb8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i8.GSR = "ENABLED";
    FD1P3AX comb8_i0_i7 (.D(comb8_71__N_2137[7]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(comb8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i7.GSR = "ENABLED";
    FD1P3AX comb8_i0_i6 (.D(comb8_71__N_2137[6]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(comb8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i6.GSR = "ENABLED";
    FD1P3AX comb8_i0_i5 (.D(comb8_71__N_2137[5]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(comb8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i5.GSR = "ENABLED";
    FD1P3AX comb8_i0_i4 (.D(comb8_71__N_2137[4]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(comb8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i4.GSR = "ENABLED";
    FD1P3AX comb8_i0_i3 (.D(comb8_71__N_2137[3]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(comb8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i3.GSR = "ENABLED";
    FD1P3AX comb8_i0_i2 (.D(comb8_71__N_2137[2]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(comb8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i2.GSR = "ENABLED";
    FD1P3AX comb8_i0_i1 (.D(comb8_71__N_2137[1]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(comb8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb8_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i71 (.D(comb7[71]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i70 (.D(comb7[70]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i69 (.D(comb7[69]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i68 (.D(comb7[68]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i67 (.D(comb7[67]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i66 (.D(comb7[66]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i65 (.D(comb7[65]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i64 (.D(comb7[64]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i63 (.D(comb7[63]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i62 (.D(comb7[62]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i61 (.D(comb7[61]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i60 (.D(comb7[60]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i59 (.D(comb7[59]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i58 (.D(comb7[58]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i57 (.D(comb7[57]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i57.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i62_1_lut (.A(comb_d6[61]), .Z(n12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i59_1_lut (.A(comb_d6[58]), .Z(n15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i59_1_lut.init = 16'h5555;
    FD1P3AX comb_d7_i0_i56 (.D(comb7[56]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i56.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i60_1_lut (.A(comb_d6[59]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i57_1_lut (.A(comb_d6[56]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i57_1_lut.init = 16'h5555;
    FD1P3AX comb_d7_i0_i55 (.D(comb7[55]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i55.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i58_1_lut (.A(comb_d6[57]), .Z(n16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i58_1_lut.init = 16'h5555;
    FD1P3AX comb_d7_i0_i54 (.D(comb7[54]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i53 (.D(comb7[53]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i52 (.D(comb7[52]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i52.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i55_1_lut (.A(comb_d6[54]), .Z(n19_adj_13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i55_1_lut.init = 16'h5555;
    FD1P3AX comb_d7_i0_i51 (.D(comb7[51]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i50 (.D(comb7[50]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i49 (.D(comb7[49]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i49.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i56_1_lut (.A(comb_d6[55]), .Z(n18_adj_14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i56_1_lut.init = 16'h5555;
    FD1P3AX comb_d7_i0_i48 (.D(comb7[48]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i47 (.D(comb7[47]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i46 (.D(comb7[46]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i45 (.D(comb7[45]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i44 (.D(comb7[44]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i43 (.D(comb7[43]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i42 (.D(comb7[42]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i42.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i53_1_lut (.A(comb_d6[52]), .Z(n21_adj_15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i53_1_lut.init = 16'h5555;
    FD1P3AX comb_d7_i0_i41 (.D(comb7[41]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i40 (.D(comb7[40]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i39 (.D(comb7[39]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i38 (.D(comb7[38]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i37 (.D(comb7[37]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i37.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i54_1_lut (.A(comb_d6[53]), .Z(n20_adj_16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i51_1_lut (.A(comb_d6[50]), .Z(n23_adj_17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i51_1_lut.init = 16'h5555;
    FD1P3AX comb_d7_i0_i36 (.D(comb7[36]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i35 (.D(comb7[35]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i34 (.D(comb7[34]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i33 (.D(comb7[33]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i32 (.D(comb7[32]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i31 (.D(comb7[31]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i31.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i52_1_lut (.A(comb_d6[51]), .Z(n22_adj_18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i52_1_lut.init = 16'h5555;
    FD1P3AX comb_d7_i0_i30 (.D(comb7[30]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(comb_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i30.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i49_1_lut (.A(comb_d6[48]), .Z(n25_adj_19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i50_1_lut (.A(comb_d6[49]), .Z(n24_adj_20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i50_1_lut.init = 16'h5555;
    FD1P3AX comb_d7_i0_i29 (.D(comb7[29]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i28 (.D(comb7[28]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i27 (.D(comb7[27]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i26 (.D(comb7[26]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i25 (.D(comb7[25]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i24 (.D(comb7[24]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i23 (.D(comb7[23]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i22 (.D(comb7[22]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i21 (.D(comb7[21]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i20 (.D(comb7[20]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i19 (.D(comb7[19]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i18 (.D(comb7[18]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i17 (.D(comb7[17]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i16 (.D(comb7[16]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i15 (.D(comb7[15]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i14 (.D(comb7[14]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i13 (.D(comb7[13]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i12 (.D(comb7[12]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i11 (.D(comb7[11]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i10 (.D(comb7[10]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i9 (.D(comb7[9]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i8 (.D(comb7[8]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i7 (.D(comb7[7]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i6 (.D(comb7[6]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i5 (.D(comb7[5]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i5.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i47_1_lut (.A(comb_d6[46]), .Z(n27_adj_21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i48_1_lut (.A(comb_d6[47]), .Z(n26_adj_22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i48_1_lut.init = 16'h5555;
    FD1P3AX comb_d7_i0_i4 (.D(comb7[4]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i3 (.D(comb7[3]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i2 (.D(comb7[2]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i1 (.D(comb7[1]), .SP(clk_80mhz_enable_550), .CK(clk_80mhz), 
            .Q(comb_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX comb7_i0_i71 (.D(comb7_71__N_2065[71]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i71.GSR = "ENABLED";
    FD1P3AX comb7_i0_i70 (.D(comb7_71__N_2065[70]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i70.GSR = "ENABLED";
    FD1P3AX comb7_i0_i69 (.D(comb7_71__N_2065[69]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i69.GSR = "ENABLED";
    FD1P3AX comb7_i0_i68 (.D(comb7_71__N_2065[68]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i68.GSR = "ENABLED";
    FD1P3AX comb7_i0_i67 (.D(comb7_71__N_2065[67]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i67.GSR = "ENABLED";
    FD1P3AX comb7_i0_i66 (.D(comb7_71__N_2065[66]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i66.GSR = "ENABLED";
    FD1P3AX comb7_i0_i65 (.D(comb7_71__N_2065[65]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i65.GSR = "ENABLED";
    FD1P3AX comb7_i0_i64 (.D(comb7_71__N_2065[64]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i64.GSR = "ENABLED";
    FD1P3AX comb7_i0_i63 (.D(comb7_71__N_2065[63]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i63.GSR = "ENABLED";
    FD1P3AX comb7_i0_i62 (.D(comb7_71__N_2065[62]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i62.GSR = "ENABLED";
    FD1P3AX comb7_i0_i61 (.D(comb7_71__N_2065[61]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i61.GSR = "ENABLED";
    FD1P3AX comb7_i0_i60 (.D(comb7_71__N_2065[60]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i60.GSR = "ENABLED";
    FD1P3AX comb7_i0_i59 (.D(comb7_71__N_2065[59]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i59.GSR = "ENABLED";
    FD1P3AX comb7_i0_i58 (.D(comb7_71__N_2065[58]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i58.GSR = "ENABLED";
    FD1P3AX comb7_i0_i57 (.D(comb7_71__N_2065[57]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i57.GSR = "ENABLED";
    FD1P3AX comb7_i0_i56 (.D(comb7_71__N_2065[56]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i56.GSR = "ENABLED";
    FD1P3AX comb7_i0_i55 (.D(comb7_71__N_2065[55]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i55.GSR = "ENABLED";
    FD1P3AX comb7_i0_i54 (.D(comb7_71__N_2065[54]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i54.GSR = "ENABLED";
    FD1P3AX comb7_i0_i53 (.D(comb7_71__N_2065[53]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i53.GSR = "ENABLED";
    FD1P3AX comb7_i0_i52 (.D(comb7_71__N_2065[52]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i52.GSR = "ENABLED";
    FD1P3AX comb7_i0_i51 (.D(comb7_71__N_2065[51]), .SP(clk_80mhz_enable_550), 
            .CK(clk_80mhz), .Q(comb7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i51.GSR = "ENABLED";
    FD1P3AX comb7_i0_i50 (.D(comb7_71__N_2065[50]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i50.GSR = "ENABLED";
    FD1P3AX comb7_i0_i49 (.D(comb7_71__N_2065[49]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i49.GSR = "ENABLED";
    FD1P3AX comb7_i0_i48 (.D(comb7_71__N_2065[48]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i48.GSR = "ENABLED";
    FD1P3AX comb7_i0_i47 (.D(comb7_71__N_2065[47]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i47.GSR = "ENABLED";
    FD1P3AX comb7_i0_i46 (.D(comb7_71__N_2065[46]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i46.GSR = "ENABLED";
    FD1P3AX comb7_i0_i45 (.D(comb7_71__N_2065[45]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i45.GSR = "ENABLED";
    FD1P3AX comb7_i0_i44 (.D(comb7_71__N_2065[44]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i44.GSR = "ENABLED";
    FD1P3AX comb7_i0_i43 (.D(comb7_71__N_2065[43]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i43.GSR = "ENABLED";
    FD1P3AX comb7_i0_i42 (.D(comb7_71__N_2065[42]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i42.GSR = "ENABLED";
    FD1P3AX comb7_i0_i41 (.D(comb7_71__N_2065[41]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i41.GSR = "ENABLED";
    FD1P3AX comb7_i0_i40 (.D(comb7_71__N_2065[40]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i40.GSR = "ENABLED";
    FD1P3AX comb7_i0_i39 (.D(comb7_71__N_2065[39]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i39.GSR = "ENABLED";
    FD1P3AX comb7_i0_i38 (.D(comb7_71__N_2065[38]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i38.GSR = "ENABLED";
    FD1P3AX comb7_i0_i37 (.D(comb7_71__N_2065[37]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i37.GSR = "ENABLED";
    FD1P3AX comb7_i0_i36 (.D(comb7_71__N_2065[36]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i36.GSR = "ENABLED";
    FD1P3AX comb7_i0_i35 (.D(comb7_71__N_2065[35]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i35.GSR = "ENABLED";
    FD1P3AX comb7_i0_i34 (.D(comb7_71__N_2065[34]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i34.GSR = "ENABLED";
    FD1P3AX comb7_i0_i33 (.D(comb7_71__N_2065[33]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i33.GSR = "ENABLED";
    FD1P3AX comb7_i0_i32 (.D(comb7_71__N_2065[32]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i32.GSR = "ENABLED";
    FD1P3AX comb7_i0_i31 (.D(comb7_71__N_2065[31]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i31.GSR = "ENABLED";
    FD1P3AX comb7_i0_i30 (.D(comb7_71__N_2065[30]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i30.GSR = "ENABLED";
    FD1P3AX comb7_i0_i29 (.D(comb7_71__N_2065[29]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i29.GSR = "ENABLED";
    FD1P3AX comb7_i0_i28 (.D(comb7_71__N_2065[28]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i28.GSR = "ENABLED";
    FD1P3AX comb7_i0_i27 (.D(comb7_71__N_2065[27]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i27.GSR = "ENABLED";
    FD1P3AX comb7_i0_i26 (.D(comb7_71__N_2065[26]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i26.GSR = "ENABLED";
    FD1P3AX comb7_i0_i25 (.D(comb7_71__N_2065[25]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i25.GSR = "ENABLED";
    FD1P3AX comb7_i0_i24 (.D(comb7_71__N_2065[24]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i24.GSR = "ENABLED";
    FD1P3AX comb7_i0_i23 (.D(comb7_71__N_2065[23]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i23.GSR = "ENABLED";
    FD1P3AX comb7_i0_i22 (.D(comb7_71__N_2065[22]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i22.GSR = "ENABLED";
    FD1P3AX comb7_i0_i21 (.D(comb7_71__N_2065[21]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i21.GSR = "ENABLED";
    FD1P3AX comb7_i0_i20 (.D(comb7_71__N_2065[20]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i20.GSR = "ENABLED";
    FD1P3AX comb7_i0_i19 (.D(comb7_71__N_2065[19]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i19.GSR = "ENABLED";
    FD1P3AX comb7_i0_i18 (.D(comb7_71__N_2065[18]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i18.GSR = "ENABLED";
    FD1P3AX comb7_i0_i17 (.D(comb7_71__N_2065[17]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i17.GSR = "ENABLED";
    FD1P3AX comb7_i0_i16 (.D(comb7_71__N_2065[16]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i16.GSR = "ENABLED";
    FD1P3AX comb7_i0_i15 (.D(comb7_71__N_2065[15]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i15.GSR = "ENABLED";
    FD1P3AX comb7_i0_i14 (.D(comb7_71__N_2065[14]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i14.GSR = "ENABLED";
    FD1P3AX comb7_i0_i13 (.D(comb7_71__N_2065[13]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i13.GSR = "ENABLED";
    FD1P3AX comb7_i0_i12 (.D(comb7_71__N_2065[12]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i12.GSR = "ENABLED";
    FD1P3AX comb7_i0_i11 (.D(comb7_71__N_2065[11]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i11.GSR = "ENABLED";
    FD1P3AX comb7_i0_i10 (.D(comb7_71__N_2065[10]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i10.GSR = "ENABLED";
    FD1P3AX comb7_i0_i9 (.D(comb7_71__N_2065[9]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i9.GSR = "ENABLED";
    FD1P3AX comb7_i0_i8 (.D(comb7_71__N_2065[8]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i8.GSR = "ENABLED";
    FD1P3AX comb7_i0_i7 (.D(comb7_71__N_2065[7]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i7.GSR = "ENABLED";
    FD1P3AX comb7_i0_i6 (.D(comb7_71__N_2065[6]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i6.GSR = "ENABLED";
    FD1P3AX comb7_i0_i5 (.D(comb7_71__N_2065[5]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i5.GSR = "ENABLED";
    FD1P3AX comb7_i0_i4 (.D(comb7_71__N_2065[4]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i4.GSR = "ENABLED";
    FD1P3AX comb7_i0_i3 (.D(comb7_71__N_2065[3]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i3.GSR = "ENABLED";
    FD1P3AX comb7_i0_i2 (.D(comb7_71__N_2065[2]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i2.GSR = "ENABLED";
    FD1P3AX comb7_i0_i1 (.D(comb7_71__N_2065[1]), .SP(clk_80mhz_enable_600), 
            .CK(clk_80mhz), .Q(comb7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb7_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i71 (.D(comb6[71]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i70 (.D(comb6[70]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i69 (.D(comb6[69]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i68 (.D(comb6[68]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i67 (.D(comb6[67]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i66 (.D(comb6[66]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i65 (.D(comb6[65]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i64 (.D(comb6[64]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i63 (.D(comb6[63]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i62 (.D(comb6[62]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i61 (.D(comb6[61]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i60 (.D(comb6[60]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i59 (.D(comb6[59]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i58 (.D(comb6[58]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i57 (.D(comb6[57]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i56 (.D(comb6[56]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i55 (.D(comb6[55]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i54 (.D(comb6[54]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i53 (.D(comb6[53]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i52 (.D(comb6[52]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i51 (.D(comb6[51]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i50 (.D(comb6[50]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i49 (.D(comb6[49]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i48 (.D(comb6[48]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i47 (.D(comb6[47]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i46 (.D(comb6[46]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i45 (.D(comb6[45]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i45.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i45_1_lut (.A(comb_d6[44]), .Z(n29_adj_23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i45_1_lut.init = 16'h5555;
    FD1P3AX comb_d6_i0_i44 (.D(comb6[44]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i43 (.D(comb6[43]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i42 (.D(comb6[42]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i41 (.D(comb6[41]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i40 (.D(comb6[40]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i39 (.D(comb6[39]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i38 (.D(comb6[38]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i37 (.D(comb6[37]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i36 (.D(comb6[36]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i35 (.D(comb6[35]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i34 (.D(comb6[34]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i33 (.D(comb6[33]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i32 (.D(comb6[32]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i31 (.D(comb6[31]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i30 (.D(comb6[30]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i29 (.D(comb6[29]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i28 (.D(comb6[28]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i27 (.D(comb6[27]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i26 (.D(comb6[26]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i25 (.D(comb6[25]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i24 (.D(comb6[24]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i23 (.D(comb6[23]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i22 (.D(comb6[22]), .SP(clk_80mhz_enable_652), .CK(clk_80mhz), 
            .Q(comb_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i21 (.D(comb6[21]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i20 (.D(comb6[20]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i19 (.D(comb6[19]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i18 (.D(comb6[18]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i17 (.D(comb6[17]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i16 (.D(comb6[16]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i15 (.D(comb6[15]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i14 (.D(comb6[14]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i13 (.D(comb6[13]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i12 (.D(comb6[12]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i11 (.D(comb6[11]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i10 (.D(comb6[10]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i9 (.D(comb6[9]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i8 (.D(comb6[8]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i7 (.D(comb6[7]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i6 (.D(comb6[6]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i5 (.D(comb6[5]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i4 (.D(comb6[4]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i3 (.D(comb6[3]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i2 (.D(comb6[2]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i1 (.D(comb6[1]), .SP(clk_80mhz_enable_702), .CK(clk_80mhz), 
            .Q(comb_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX comb6_i0_i71 (.D(comb6_71__N_1993[71]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i71.GSR = "ENABLED";
    FD1P3AX comb6_i0_i70 (.D(comb6_71__N_1993[70]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i70.GSR = "ENABLED";
    FD1P3AX comb6_i0_i69 (.D(comb6_71__N_1993[69]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i69.GSR = "ENABLED";
    FD1P3AX comb6_i0_i68 (.D(comb6_71__N_1993[68]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i68.GSR = "ENABLED";
    FD1P3AX comb6_i0_i67 (.D(comb6_71__N_1993[67]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i67.GSR = "ENABLED";
    FD1P3AX comb6_i0_i66 (.D(comb6_71__N_1993[66]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i66.GSR = "ENABLED";
    FD1P3AX comb6_i0_i65 (.D(comb6_71__N_1993[65]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i65.GSR = "ENABLED";
    FD1P3AX comb6_i0_i64 (.D(comb6_71__N_1993[64]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i64.GSR = "ENABLED";
    FD1P3AX comb6_i0_i63 (.D(comb6_71__N_1993[63]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i63.GSR = "ENABLED";
    FD1P3AX comb6_i0_i62 (.D(comb6_71__N_1993[62]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i62.GSR = "ENABLED";
    FD1P3AX comb6_i0_i61 (.D(comb6_71__N_1993[61]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i61.GSR = "ENABLED";
    FD1P3AX comb6_i0_i60 (.D(comb6_71__N_1993[60]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i60.GSR = "ENABLED";
    FD1P3AX comb6_i0_i59 (.D(comb6_71__N_1993[59]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i59.GSR = "ENABLED";
    FD1P3AX comb6_i0_i58 (.D(comb6_71__N_1993[58]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i58.GSR = "ENABLED";
    FD1P3AX comb6_i0_i57 (.D(comb6_71__N_1993[57]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i57.GSR = "ENABLED";
    FD1P3AX comb6_i0_i56 (.D(comb6_71__N_1993[56]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i56.GSR = "ENABLED";
    FD1P3AX comb6_i0_i55 (.D(comb6_71__N_1993[55]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i55.GSR = "ENABLED";
    FD1P3AX comb6_i0_i54 (.D(comb6_71__N_1993[54]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i54.GSR = "ENABLED";
    FD1P3AX comb6_i0_i53 (.D(comb6_71__N_1993[53]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i53.GSR = "ENABLED";
    FD1P3AX comb6_i0_i52 (.D(comb6_71__N_1993[52]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i52.GSR = "ENABLED";
    FD1P3AX comb6_i0_i51 (.D(comb6_71__N_1993[51]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i51.GSR = "ENABLED";
    FD1P3AX comb6_i0_i50 (.D(comb6_71__N_1993[50]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i50.GSR = "ENABLED";
    FD1P3AX comb6_i0_i49 (.D(comb6_71__N_1993[49]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i49.GSR = "ENABLED";
    FD1P3AX comb6_i0_i48 (.D(comb6_71__N_1993[48]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i48.GSR = "ENABLED";
    FD1P3AX comb6_i0_i47 (.D(comb6_71__N_1993[47]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i47.GSR = "ENABLED";
    FD1P3AX comb6_i0_i46 (.D(comb6_71__N_1993[46]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i46.GSR = "ENABLED";
    FD1P3AX comb6_i0_i45 (.D(comb6_71__N_1993[45]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i45.GSR = "ENABLED";
    FD1P3AX comb6_i0_i44 (.D(comb6_71__N_1993[44]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i44.GSR = "ENABLED";
    FD1P3AX comb6_i0_i43 (.D(comb6_71__N_1993[43]), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(comb6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i43.GSR = "ENABLED";
    FD1P3AX comb6_i0_i42 (.D(comb6_71__N_1993[42]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i42.GSR = "ENABLED";
    FD1P3AX comb6_i0_i41 (.D(comb6_71__N_1993[41]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i41.GSR = "ENABLED";
    FD1P3AX comb6_i0_i40 (.D(comb6_71__N_1993[40]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i40.GSR = "ENABLED";
    FD1P3AX comb6_i0_i39 (.D(comb6_71__N_1993[39]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i39.GSR = "ENABLED";
    FD1P3AX comb6_i0_i38 (.D(comb6_71__N_1993[38]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i38.GSR = "ENABLED";
    FD1P3AX comb6_i0_i37 (.D(comb6_71__N_1993[37]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i37.GSR = "ENABLED";
    FD1P3AX comb6_i0_i36 (.D(comb6_71__N_1993[36]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i36.GSR = "ENABLED";
    FD1P3AX comb6_i0_i35 (.D(comb6_71__N_1993[35]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i35.GSR = "ENABLED";
    FD1P3AX comb6_i0_i34 (.D(comb6_71__N_1993[34]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i34.GSR = "ENABLED";
    FD1P3AX comb6_i0_i33 (.D(comb6_71__N_1993[33]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i33.GSR = "ENABLED";
    FD1P3AX comb6_i0_i32 (.D(comb6_71__N_1993[32]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i32.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i46_1_lut (.A(comb_d6[45]), .Z(n28_adj_24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i46_1_lut.init = 16'h5555;
    FD1P3AX comb6_i0_i31 (.D(comb6_71__N_1993[31]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i31.GSR = "ENABLED";
    FD1P3AX comb6_i0_i30 (.D(comb6_71__N_1993[30]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i30.GSR = "ENABLED";
    FD1P3AX comb6_i0_i29 (.D(comb6_71__N_1993[29]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i29.GSR = "ENABLED";
    FD1P3AX comb6_i0_i28 (.D(comb6_71__N_1993[28]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i28.GSR = "ENABLED";
    FD1P3AX comb6_i0_i27 (.D(comb6_71__N_1993[27]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i27.GSR = "ENABLED";
    FD1P3AX comb6_i0_i26 (.D(comb6_71__N_1993[26]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i26.GSR = "ENABLED";
    FD1P3AX comb6_i0_i25 (.D(comb6_71__N_1993[25]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i25.GSR = "ENABLED";
    FD1P3AX comb6_i0_i24 (.D(comb6_71__N_1993[24]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i24.GSR = "ENABLED";
    FD1P3AX comb6_i0_i23 (.D(comb6_71__N_1993[23]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i23.GSR = "ENABLED";
    FD1P3AX comb6_i0_i22 (.D(comb6_71__N_1993[22]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i22.GSR = "ENABLED";
    FD1P3AX comb6_i0_i21 (.D(comb6_71__N_1993[21]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i21.GSR = "ENABLED";
    FD1P3AX comb6_i0_i20 (.D(comb6_71__N_1993[20]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i20.GSR = "ENABLED";
    FD1P3AX comb6_i0_i19 (.D(comb6_71__N_1993[19]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i19.GSR = "ENABLED";
    FD1P3AX comb6_i0_i18 (.D(comb6_71__N_1993[18]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i18.GSR = "ENABLED";
    FD1P3AX comb6_i0_i17 (.D(comb6_71__N_1993[17]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i17.GSR = "ENABLED";
    FD1P3AX comb6_i0_i16 (.D(comb6_71__N_1993[16]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i16.GSR = "ENABLED";
    FD1P3AX comb6_i0_i15 (.D(comb6_71__N_1993[15]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i15.GSR = "ENABLED";
    FD1P3AX comb6_i0_i14 (.D(comb6_71__N_1993[14]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i14.GSR = "ENABLED";
    FD1P3AX comb6_i0_i13 (.D(comb6_71__N_1993[13]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i13.GSR = "ENABLED";
    FD1P3AX comb6_i0_i12 (.D(comb6_71__N_1993[12]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i12.GSR = "ENABLED";
    FD1P3AX comb6_i0_i11 (.D(comb6_71__N_1993[11]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i11.GSR = "ENABLED";
    FD1P3AX comb6_i0_i10 (.D(comb6_71__N_1993[10]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i10.GSR = "ENABLED";
    FD1P3AX comb6_i0_i9 (.D(comb6_71__N_1993[9]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i9.GSR = "ENABLED";
    FD1P3AX comb6_i0_i8 (.D(comb6_71__N_1993[8]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i8.GSR = "ENABLED";
    FD1P3AX comb6_i0_i7 (.D(comb6_71__N_1993[7]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i7.GSR = "ENABLED";
    FD1P3AX comb6_i0_i6 (.D(comb6_71__N_1993[6]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i6.GSR = "ENABLED";
    FD1P3AX comb6_i0_i5 (.D(comb6_71__N_1993[5]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i5.GSR = "ENABLED";
    FD1P3AX comb6_i0_i4 (.D(comb6_71__N_1993[4]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i4.GSR = "ENABLED";
    FD1P3AX comb6_i0_i3 (.D(comb6_71__N_1993[3]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i3.GSR = "ENABLED";
    FD1P3AX comb6_i0_i2 (.D(comb6_71__N_1993[2]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i2.GSR = "ENABLED";
    FD1P3AX comb6_i0_i1 (.D(comb6_71__N_1993[1]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(comb6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam comb6_i0_i1.GSR = "ENABLED";
    FD1S3AX integrator5_i71 (.D(integrator5_71__N_1248[71]), .CK(clk_80mhz), 
            .Q(integrator5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i71.GSR = "ENABLED";
    FD1S3AX integrator5_i70 (.D(integrator5_71__N_1248[70]), .CK(clk_80mhz), 
            .Q(integrator5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i70.GSR = "ENABLED";
    FD1S3AX integrator5_i69 (.D(integrator5_71__N_1248[69]), .CK(clk_80mhz), 
            .Q(integrator5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i69.GSR = "ENABLED";
    FD1S3AX integrator5_i68 (.D(integrator5_71__N_1248[68]), .CK(clk_80mhz), 
            .Q(integrator5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i68.GSR = "ENABLED";
    FD1S3AX integrator5_i67 (.D(integrator5_71__N_1248[67]), .CK(clk_80mhz), 
            .Q(integrator5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i67.GSR = "ENABLED";
    FD1S3AX integrator5_i66 (.D(integrator5_71__N_1248[66]), .CK(clk_80mhz), 
            .Q(integrator5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i66.GSR = "ENABLED";
    FD1S3AX integrator5_i65 (.D(integrator5_71__N_1248[65]), .CK(clk_80mhz), 
            .Q(integrator5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i65.GSR = "ENABLED";
    FD1S3AX integrator5_i64 (.D(integrator5_71__N_1248[64]), .CK(clk_80mhz), 
            .Q(integrator5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i64.GSR = "ENABLED";
    FD1S3AX integrator5_i63 (.D(integrator5_71__N_1248[63]), .CK(clk_80mhz), 
            .Q(integrator5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i63.GSR = "ENABLED";
    FD1S3AX integrator5_i62 (.D(integrator5_71__N_1248[62]), .CK(clk_80mhz), 
            .Q(integrator5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i62.GSR = "ENABLED";
    FD1S3AX integrator5_i61 (.D(integrator5_71__N_1248[61]), .CK(clk_80mhz), 
            .Q(integrator5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i61.GSR = "ENABLED";
    FD1S3AX integrator5_i60 (.D(integrator5_71__N_1248[60]), .CK(clk_80mhz), 
            .Q(integrator5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i60.GSR = "ENABLED";
    FD1S3AX integrator5_i59 (.D(integrator5_71__N_1248[59]), .CK(clk_80mhz), 
            .Q(integrator5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i59.GSR = "ENABLED";
    FD1S3AX integrator5_i58 (.D(integrator5_71__N_1248[58]), .CK(clk_80mhz), 
            .Q(integrator5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i58.GSR = "ENABLED";
    FD1S3AX integrator5_i57 (.D(integrator5_71__N_1248[57]), .CK(clk_80mhz), 
            .Q(integrator5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i57.GSR = "ENABLED";
    FD1S3AX integrator5_i56 (.D(integrator5_71__N_1248[56]), .CK(clk_80mhz), 
            .Q(integrator5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i56.GSR = "ENABLED";
    FD1S3AX integrator5_i55 (.D(integrator5_71__N_1248[55]), .CK(clk_80mhz), 
            .Q(integrator5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i55.GSR = "ENABLED";
    FD1S3AX integrator5_i54 (.D(integrator5_71__N_1248[54]), .CK(clk_80mhz), 
            .Q(integrator5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i54.GSR = "ENABLED";
    FD1S3AX integrator5_i53 (.D(integrator5_71__N_1248[53]), .CK(clk_80mhz), 
            .Q(integrator5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i53.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i67_1_lut (.A(integrator_d_tmp[66]), .Z(n7_adj_25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i67_1_lut.init = 16'h5555;
    FD1S3AX integrator5_i52 (.D(integrator5_71__N_1248[52]), .CK(clk_80mhz), 
            .Q(integrator5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i52.GSR = "ENABLED";
    FD1S3AX integrator5_i51 (.D(integrator5_71__N_1248[51]), .CK(clk_80mhz), 
            .Q(integrator5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i51.GSR = "ENABLED";
    FD1S3AX integrator5_i50 (.D(integrator5_71__N_1248[50]), .CK(clk_80mhz), 
            .Q(integrator5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i50.GSR = "ENABLED";
    FD1S3AX integrator5_i49 (.D(integrator5_71__N_1248[49]), .CK(clk_80mhz), 
            .Q(integrator5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i49.GSR = "ENABLED";
    FD1S3AX integrator5_i48 (.D(integrator5_71__N_1248[48]), .CK(clk_80mhz), 
            .Q(integrator5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i48.GSR = "ENABLED";
    FD1S3AX integrator5_i47 (.D(integrator5_71__N_1248[47]), .CK(clk_80mhz), 
            .Q(integrator5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i47.GSR = "ENABLED";
    FD1S3AX integrator5_i46 (.D(integrator5_71__N_1248[46]), .CK(clk_80mhz), 
            .Q(integrator5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i46.GSR = "ENABLED";
    FD1S3AX integrator5_i45 (.D(integrator5_71__N_1248[45]), .CK(clk_80mhz), 
            .Q(integrator5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i45.GSR = "ENABLED";
    FD1S3AX integrator5_i44 (.D(integrator5_71__N_1248[44]), .CK(clk_80mhz), 
            .Q(integrator5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i44.GSR = "ENABLED";
    FD1S3AX integrator5_i43 (.D(integrator5_71__N_1248[43]), .CK(clk_80mhz), 
            .Q(integrator5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i43.GSR = "ENABLED";
    FD1S3AX integrator5_i42 (.D(integrator5_71__N_1248[42]), .CK(clk_80mhz), 
            .Q(integrator5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i42.GSR = "ENABLED";
    FD1S3AX integrator5_i41 (.D(integrator5_71__N_1248[41]), .CK(clk_80mhz), 
            .Q(integrator5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i41.GSR = "ENABLED";
    FD1S3AX integrator5_i40 (.D(integrator5_71__N_1248[40]), .CK(clk_80mhz), 
            .Q(integrator5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i40.GSR = "ENABLED";
    FD1S3AX integrator5_i39 (.D(integrator5_71__N_1248[39]), .CK(clk_80mhz), 
            .Q(integrator5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i39.GSR = "ENABLED";
    FD1S3AX integrator5_i38 (.D(integrator5_71__N_1248[38]), .CK(clk_80mhz), 
            .Q(integrator5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i38.GSR = "ENABLED";
    FD1S3AX integrator5_i37 (.D(integrator5_71__N_1248[37]), .CK(clk_80mhz), 
            .Q(integrator5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i37.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i43_1_lut (.A(comb_d6[42]), .Z(n31_adj_26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i43_1_lut.init = 16'h5555;
    FD1S3AX integrator5_i36 (.D(integrator5_71__N_1248[36]), .CK(clk_80mhz), 
            .Q(integrator5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i36.GSR = "ENABLED";
    FD1S3AX integrator5_i35 (.D(integrator5_71__N_1248[35]), .CK(clk_80mhz), 
            .Q(integrator5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i35.GSR = "ENABLED";
    FD1S3AX integrator5_i34 (.D(integrator5_71__N_1248[34]), .CK(clk_80mhz), 
            .Q(integrator5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i34.GSR = "ENABLED";
    FD1S3AX integrator5_i33 (.D(integrator5_71__N_1248[33]), .CK(clk_80mhz), 
            .Q(integrator5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i33.GSR = "ENABLED";
    FD1S3AX integrator5_i32 (.D(integrator5_71__N_1248[32]), .CK(clk_80mhz), 
            .Q(integrator5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i32.GSR = "ENABLED";
    FD1S3AX integrator5_i31 (.D(integrator5_71__N_1248[31]), .CK(clk_80mhz), 
            .Q(integrator5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i31.GSR = "ENABLED";
    FD1S3AX integrator5_i30 (.D(integrator5_71__N_1248[30]), .CK(clk_80mhz), 
            .Q(integrator5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i30.GSR = "ENABLED";
    FD1S3AX integrator5_i29 (.D(integrator5_71__N_1248[29]), .CK(clk_80mhz), 
            .Q(integrator5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i29.GSR = "ENABLED";
    FD1S3AX integrator5_i28 (.D(integrator5_71__N_1248[28]), .CK(clk_80mhz), 
            .Q(integrator5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i28.GSR = "ENABLED";
    FD1S3AX integrator5_i27 (.D(integrator5_71__N_1248[27]), .CK(clk_80mhz), 
            .Q(integrator5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i27.GSR = "ENABLED";
    FD1S3AX integrator5_i26 (.D(integrator5_71__N_1248[26]), .CK(clk_80mhz), 
            .Q(integrator5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i26.GSR = "ENABLED";
    FD1S3AX integrator5_i25 (.D(integrator5_71__N_1248[25]), .CK(clk_80mhz), 
            .Q(integrator5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i25.GSR = "ENABLED";
    FD1S3AX integrator5_i24 (.D(integrator5_71__N_1248[24]), .CK(clk_80mhz), 
            .Q(integrator5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i24.GSR = "ENABLED";
    FD1S3AX integrator5_i23 (.D(integrator5_71__N_1248[23]), .CK(clk_80mhz), 
            .Q(integrator5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i23.GSR = "ENABLED";
    FD1S3AX integrator5_i22 (.D(integrator5_71__N_1248[22]), .CK(clk_80mhz), 
            .Q(integrator5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i22.GSR = "ENABLED";
    FD1S3AX integrator5_i21 (.D(integrator5_71__N_1248[21]), .CK(clk_80mhz), 
            .Q(integrator5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i21.GSR = "ENABLED";
    FD1S3AX integrator5_i20 (.D(integrator5_71__N_1248[20]), .CK(clk_80mhz), 
            .Q(integrator5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i20.GSR = "ENABLED";
    FD1S3AX integrator5_i19 (.D(integrator5_71__N_1248[19]), .CK(clk_80mhz), 
            .Q(integrator5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i19.GSR = "ENABLED";
    FD1S3AX integrator5_i18 (.D(integrator5_71__N_1248[18]), .CK(clk_80mhz), 
            .Q(integrator5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i18.GSR = "ENABLED";
    FD1S3AX integrator5_i17 (.D(integrator5_71__N_1248[17]), .CK(clk_80mhz), 
            .Q(integrator5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i17.GSR = "ENABLED";
    FD1S3AX integrator5_i16 (.D(integrator5_71__N_1248[16]), .CK(clk_80mhz), 
            .Q(integrator5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i16.GSR = "ENABLED";
    FD1S3AX integrator5_i15 (.D(integrator5_71__N_1248[15]), .CK(clk_80mhz), 
            .Q(integrator5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i15.GSR = "ENABLED";
    FD1S3AX integrator5_i14 (.D(integrator5_71__N_1248[14]), .CK(clk_80mhz), 
            .Q(integrator5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i14.GSR = "ENABLED";
    FD1S3AX integrator5_i13 (.D(integrator5_71__N_1248[13]), .CK(clk_80mhz), 
            .Q(integrator5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i13.GSR = "ENABLED";
    FD1S3AX integrator5_i12 (.D(integrator5_71__N_1248[12]), .CK(clk_80mhz), 
            .Q(integrator5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i12.GSR = "ENABLED";
    FD1S3AX integrator5_i11 (.D(integrator5_71__N_1248[11]), .CK(clk_80mhz), 
            .Q(integrator5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i11.GSR = "ENABLED";
    FD1S3AX integrator5_i10 (.D(integrator5_71__N_1248[10]), .CK(clk_80mhz), 
            .Q(integrator5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i10.GSR = "ENABLED";
    FD1S3AX integrator5_i9 (.D(integrator5_71__N_1248[9]), .CK(clk_80mhz), 
            .Q(integrator5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i9.GSR = "ENABLED";
    FD1S3AX integrator5_i8 (.D(integrator5_71__N_1248[8]), .CK(clk_80mhz), 
            .Q(integrator5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i8.GSR = "ENABLED";
    FD1S3AX integrator5_i7 (.D(integrator5_71__N_1248[7]), .CK(clk_80mhz), 
            .Q(integrator5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i7.GSR = "ENABLED";
    FD1S3AX integrator5_i6 (.D(integrator5_71__N_1248[6]), .CK(clk_80mhz), 
            .Q(integrator5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i6.GSR = "ENABLED";
    FD1S3AX integrator5_i5 (.D(integrator5_71__N_1248[5]), .CK(clk_80mhz), 
            .Q(integrator5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i5.GSR = "ENABLED";
    FD1S3AX integrator5_i4 (.D(integrator5_71__N_1248[4]), .CK(clk_80mhz), 
            .Q(integrator5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i4.GSR = "ENABLED";
    FD1S3AX integrator5_i3 (.D(integrator5_71__N_1248[3]), .CK(clk_80mhz), 
            .Q(integrator5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i3.GSR = "ENABLED";
    FD1S3AX integrator5_i2 (.D(integrator5_71__N_1248[2]), .CK(clk_80mhz), 
            .Q(integrator5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i2.GSR = "ENABLED";
    FD1S3AX integrator5_i1 (.D(integrator5_71__N_1248[1]), .CK(clk_80mhz), 
            .Q(integrator5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator5_i1.GSR = "ENABLED";
    FD1S3AX integrator4_i71 (.D(integrator4_71__N_1176[71]), .CK(clk_80mhz), 
            .Q(integrator4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i71.GSR = "ENABLED";
    FD1S3AX integrator4_i70 (.D(integrator4_71__N_1176[70]), .CK(clk_80mhz), 
            .Q(integrator4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i70.GSR = "ENABLED";
    FD1S3AX integrator4_i69 (.D(integrator4_71__N_1176[69]), .CK(clk_80mhz), 
            .Q(integrator4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i69.GSR = "ENABLED";
    FD1S3AX integrator4_i68 (.D(integrator4_71__N_1176[68]), .CK(clk_80mhz), 
            .Q(integrator4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i68.GSR = "ENABLED";
    FD1S3AX integrator4_i67 (.D(integrator4_71__N_1176[67]), .CK(clk_80mhz), 
            .Q(integrator4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i67.GSR = "ENABLED";
    FD1S3AX integrator4_i66 (.D(integrator4_71__N_1176[66]), .CK(clk_80mhz), 
            .Q(integrator4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i66.GSR = "ENABLED";
    FD1S3AX integrator4_i65 (.D(integrator4_71__N_1176[65]), .CK(clk_80mhz), 
            .Q(integrator4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i65.GSR = "ENABLED";
    FD1S3AX integrator4_i64 (.D(integrator4_71__N_1176[64]), .CK(clk_80mhz), 
            .Q(integrator4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i64.GSR = "ENABLED";
    FD1S3AX integrator4_i63 (.D(integrator4_71__N_1176[63]), .CK(clk_80mhz), 
            .Q(integrator4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i63.GSR = "ENABLED";
    FD1S3AX integrator4_i62 (.D(integrator4_71__N_1176[62]), .CK(clk_80mhz), 
            .Q(integrator4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i62.GSR = "ENABLED";
    FD1S3AX integrator4_i61 (.D(integrator4_71__N_1176[61]), .CK(clk_80mhz), 
            .Q(integrator4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i61.GSR = "ENABLED";
    FD1S3AX integrator4_i60 (.D(integrator4_71__N_1176[60]), .CK(clk_80mhz), 
            .Q(integrator4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i60.GSR = "ENABLED";
    FD1S3AX integrator4_i59 (.D(integrator4_71__N_1176[59]), .CK(clk_80mhz), 
            .Q(integrator4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i59.GSR = "ENABLED";
    FD1S3AX integrator4_i58 (.D(integrator4_71__N_1176[58]), .CK(clk_80mhz), 
            .Q(integrator4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i58.GSR = "ENABLED";
    FD1S3AX integrator4_i57 (.D(integrator4_71__N_1176[57]), .CK(clk_80mhz), 
            .Q(integrator4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i57.GSR = "ENABLED";
    FD1S3AX integrator4_i56 (.D(integrator4_71__N_1176[56]), .CK(clk_80mhz), 
            .Q(integrator4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i56.GSR = "ENABLED";
    FD1S3AX integrator4_i55 (.D(integrator4_71__N_1176[55]), .CK(clk_80mhz), 
            .Q(integrator4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i55.GSR = "ENABLED";
    FD1S3AX integrator4_i54 (.D(integrator4_71__N_1176[54]), .CK(clk_80mhz), 
            .Q(integrator4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i54.GSR = "ENABLED";
    FD1S3AX integrator4_i53 (.D(integrator4_71__N_1176[53]), .CK(clk_80mhz), 
            .Q(integrator4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i53.GSR = "ENABLED";
    FD1S3AX integrator4_i52 (.D(integrator4_71__N_1176[52]), .CK(clk_80mhz), 
            .Q(integrator4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i52.GSR = "ENABLED";
    FD1S3AX integrator4_i51 (.D(integrator4_71__N_1176[51]), .CK(clk_80mhz), 
            .Q(integrator4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i51.GSR = "ENABLED";
    FD1S3AX integrator4_i50 (.D(integrator4_71__N_1176[50]), .CK(clk_80mhz), 
            .Q(integrator4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i50.GSR = "ENABLED";
    FD1S3AX integrator4_i49 (.D(integrator4_71__N_1176[49]), .CK(clk_80mhz), 
            .Q(integrator4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i49.GSR = "ENABLED";
    FD1S3AX integrator4_i48 (.D(integrator4_71__N_1176[48]), .CK(clk_80mhz), 
            .Q(integrator4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i48.GSR = "ENABLED";
    FD1S3AX integrator4_i47 (.D(integrator4_71__N_1176[47]), .CK(clk_80mhz), 
            .Q(integrator4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i47.GSR = "ENABLED";
    FD1S3AX integrator4_i46 (.D(integrator4_71__N_1176[46]), .CK(clk_80mhz), 
            .Q(integrator4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i46.GSR = "ENABLED";
    FD1S3AX integrator4_i45 (.D(integrator4_71__N_1176[45]), .CK(clk_80mhz), 
            .Q(integrator4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i45.GSR = "ENABLED";
    FD1S3AX integrator4_i44 (.D(integrator4_71__N_1176[44]), .CK(clk_80mhz), 
            .Q(integrator4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i44.GSR = "ENABLED";
    FD1S3AX integrator4_i43 (.D(integrator4_71__N_1176[43]), .CK(clk_80mhz), 
            .Q(integrator4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i43.GSR = "ENABLED";
    FD1S3AX integrator4_i42 (.D(integrator4_71__N_1176[42]), .CK(clk_80mhz), 
            .Q(integrator4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i42.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i68_1_lut (.A(integrator_d_tmp[67]), .Z(n6_adj_27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i68_1_lut.init = 16'h5555;
    FD1S3AX integrator4_i41 (.D(integrator4_71__N_1176[41]), .CK(clk_80mhz), 
            .Q(integrator4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i41.GSR = "ENABLED";
    FD1S3AX integrator4_i40 (.D(integrator4_71__N_1176[40]), .CK(clk_80mhz), 
            .Q(integrator4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i40.GSR = "ENABLED";
    FD1S3AX integrator4_i39 (.D(integrator4_71__N_1176[39]), .CK(clk_80mhz), 
            .Q(integrator4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i39.GSR = "ENABLED";
    FD1S3AX integrator4_i38 (.D(integrator4_71__N_1176[38]), .CK(clk_80mhz), 
            .Q(integrator4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i38.GSR = "ENABLED";
    FD1S3AX integrator4_i37 (.D(integrator4_71__N_1176[37]), .CK(clk_80mhz), 
            .Q(integrator4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i37.GSR = "ENABLED";
    FD1S3AX integrator4_i36 (.D(integrator4_71__N_1176[36]), .CK(clk_80mhz), 
            .Q(integrator4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i36.GSR = "ENABLED";
    FD1S3AX integrator4_i35 (.D(integrator4_71__N_1176[35]), .CK(clk_80mhz), 
            .Q(integrator4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i35.GSR = "ENABLED";
    FD1S3AX integrator4_i34 (.D(integrator4_71__N_1176[34]), .CK(clk_80mhz), 
            .Q(integrator4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i34.GSR = "ENABLED";
    FD1S3AX integrator4_i33 (.D(integrator4_71__N_1176[33]), .CK(clk_80mhz), 
            .Q(integrator4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i33.GSR = "ENABLED";
    FD1S3AX integrator4_i32 (.D(integrator4_71__N_1176[32]), .CK(clk_80mhz), 
            .Q(integrator4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i32.GSR = "ENABLED";
    FD1S3AX integrator4_i31 (.D(integrator4_71__N_1176[31]), .CK(clk_80mhz), 
            .Q(integrator4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i31.GSR = "ENABLED";
    FD1S3AX integrator4_i30 (.D(integrator4_71__N_1176[30]), .CK(clk_80mhz), 
            .Q(integrator4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i30.GSR = "ENABLED";
    FD1S3AX integrator4_i29 (.D(integrator4_71__N_1176[29]), .CK(clk_80mhz), 
            .Q(integrator4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i29.GSR = "ENABLED";
    FD1S3AX integrator4_i28 (.D(integrator4_71__N_1176[28]), .CK(clk_80mhz), 
            .Q(integrator4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i28.GSR = "ENABLED";
    FD1S3AX integrator4_i27 (.D(integrator4_71__N_1176[27]), .CK(clk_80mhz), 
            .Q(integrator4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i27.GSR = "ENABLED";
    FD1S3AX integrator4_i26 (.D(integrator4_71__N_1176[26]), .CK(clk_80mhz), 
            .Q(integrator4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i26.GSR = "ENABLED";
    FD1S3AX integrator4_i25 (.D(integrator4_71__N_1176[25]), .CK(clk_80mhz), 
            .Q(integrator4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i25.GSR = "ENABLED";
    FD1S3AX integrator4_i24 (.D(integrator4_71__N_1176[24]), .CK(clk_80mhz), 
            .Q(integrator4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i24.GSR = "ENABLED";
    FD1S3AX integrator4_i23 (.D(integrator4_71__N_1176[23]), .CK(clk_80mhz), 
            .Q(integrator4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i23.GSR = "ENABLED";
    FD1S3AX integrator4_i22 (.D(integrator4_71__N_1176[22]), .CK(clk_80mhz), 
            .Q(integrator4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i22.GSR = "ENABLED";
    FD1S3AX integrator4_i21 (.D(integrator4_71__N_1176[21]), .CK(clk_80mhz), 
            .Q(integrator4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i21.GSR = "ENABLED";
    FD1S3AX integrator4_i20 (.D(integrator4_71__N_1176[20]), .CK(clk_80mhz), 
            .Q(integrator4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i20.GSR = "ENABLED";
    FD1S3AX integrator4_i19 (.D(integrator4_71__N_1176[19]), .CK(clk_80mhz), 
            .Q(integrator4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i19.GSR = "ENABLED";
    FD1S3AX integrator4_i18 (.D(integrator4_71__N_1176[18]), .CK(clk_80mhz), 
            .Q(integrator4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i18.GSR = "ENABLED";
    FD1S3AX integrator4_i17 (.D(integrator4_71__N_1176[17]), .CK(clk_80mhz), 
            .Q(integrator4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i17.GSR = "ENABLED";
    FD1S3AX integrator4_i16 (.D(integrator4_71__N_1176[16]), .CK(clk_80mhz), 
            .Q(integrator4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i16.GSR = "ENABLED";
    FD1S3AX integrator4_i15 (.D(integrator4_71__N_1176[15]), .CK(clk_80mhz), 
            .Q(integrator4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i15.GSR = "ENABLED";
    FD1S3AX integrator4_i14 (.D(integrator4_71__N_1176[14]), .CK(clk_80mhz), 
            .Q(integrator4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i14.GSR = "ENABLED";
    FD1S3AX integrator4_i13 (.D(integrator4_71__N_1176[13]), .CK(clk_80mhz), 
            .Q(integrator4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i13.GSR = "ENABLED";
    FD1S3AX integrator4_i12 (.D(integrator4_71__N_1176[12]), .CK(clk_80mhz), 
            .Q(integrator4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i12.GSR = "ENABLED";
    FD1S3AX integrator4_i11 (.D(integrator4_71__N_1176[11]), .CK(clk_80mhz), 
            .Q(integrator4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i11.GSR = "ENABLED";
    FD1S3AX integrator4_i10 (.D(integrator4_71__N_1176[10]), .CK(clk_80mhz), 
            .Q(integrator4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i10.GSR = "ENABLED";
    FD1S3AX integrator4_i9 (.D(integrator4_71__N_1176[9]), .CK(clk_80mhz), 
            .Q(integrator4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i9.GSR = "ENABLED";
    FD1S3AX integrator4_i8 (.D(integrator4_71__N_1176[8]), .CK(clk_80mhz), 
            .Q(integrator4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i8.GSR = "ENABLED";
    FD1S3AX integrator4_i7 (.D(integrator4_71__N_1176[7]), .CK(clk_80mhz), 
            .Q(integrator4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i7.GSR = "ENABLED";
    FD1S3AX integrator4_i6 (.D(integrator4_71__N_1176[6]), .CK(clk_80mhz), 
            .Q(integrator4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i6.GSR = "ENABLED";
    FD1S3AX integrator4_i5 (.D(integrator4_71__N_1176[5]), .CK(clk_80mhz), 
            .Q(integrator4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i5.GSR = "ENABLED";
    FD1S3AX integrator4_i4 (.D(integrator4_71__N_1176[4]), .CK(clk_80mhz), 
            .Q(integrator4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i4.GSR = "ENABLED";
    FD1S3AX integrator4_i3 (.D(integrator4_71__N_1176[3]), .CK(clk_80mhz), 
            .Q(integrator4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i3.GSR = "ENABLED";
    FD1S3AX integrator4_i2 (.D(integrator4_71__N_1176[2]), .CK(clk_80mhz), 
            .Q(integrator4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i2.GSR = "ENABLED";
    FD1S3AX integrator4_i1 (.D(integrator4_71__N_1176[1]), .CK(clk_80mhz), 
            .Q(integrator4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator4_i1.GSR = "ENABLED";
    FD1S3AX integrator3_i71 (.D(integrator3_71__N_1104[71]), .CK(clk_80mhz), 
            .Q(integrator3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i71.GSR = "ENABLED";
    FD1S3AX integrator3_i70 (.D(integrator3_71__N_1104[70]), .CK(clk_80mhz), 
            .Q(integrator3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i70.GSR = "ENABLED";
    FD1S3AX integrator3_i69 (.D(integrator3_71__N_1104[69]), .CK(clk_80mhz), 
            .Q(integrator3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i69.GSR = "ENABLED";
    FD1S3AX integrator3_i68 (.D(integrator3_71__N_1104[68]), .CK(clk_80mhz), 
            .Q(integrator3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i68.GSR = "ENABLED";
    FD1S3AX integrator3_i67 (.D(integrator3_71__N_1104[67]), .CK(clk_80mhz), 
            .Q(integrator3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i67.GSR = "ENABLED";
    FD1S3AX integrator3_i66 (.D(integrator3_71__N_1104[66]), .CK(clk_80mhz), 
            .Q(integrator3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i66.GSR = "ENABLED";
    FD1S3AX integrator3_i65 (.D(integrator3_71__N_1104[65]), .CK(clk_80mhz), 
            .Q(integrator3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i65.GSR = "ENABLED";
    FD1S3AX integrator3_i64 (.D(integrator3_71__N_1104[64]), .CK(clk_80mhz), 
            .Q(integrator3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i64.GSR = "ENABLED";
    FD1S3AX integrator3_i63 (.D(integrator3_71__N_1104[63]), .CK(clk_80mhz), 
            .Q(integrator3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i63.GSR = "ENABLED";
    FD1S3AX integrator3_i62 (.D(integrator3_71__N_1104[62]), .CK(clk_80mhz), 
            .Q(integrator3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i62.GSR = "ENABLED";
    FD1S3AX integrator3_i61 (.D(integrator3_71__N_1104[61]), .CK(clk_80mhz), 
            .Q(integrator3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i61.GSR = "ENABLED";
    FD1S3AX integrator3_i60 (.D(integrator3_71__N_1104[60]), .CK(clk_80mhz), 
            .Q(integrator3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i60.GSR = "ENABLED";
    FD1S3AX integrator3_i59 (.D(integrator3_71__N_1104[59]), .CK(clk_80mhz), 
            .Q(integrator3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i59.GSR = "ENABLED";
    FD1S3AX integrator3_i58 (.D(integrator3_71__N_1104[58]), .CK(clk_80mhz), 
            .Q(integrator3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i58.GSR = "ENABLED";
    FD1S3AX integrator3_i57 (.D(integrator3_71__N_1104[57]), .CK(clk_80mhz), 
            .Q(integrator3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i57.GSR = "ENABLED";
    FD1S3AX integrator3_i56 (.D(integrator3_71__N_1104[56]), .CK(clk_80mhz), 
            .Q(integrator3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i56.GSR = "ENABLED";
    FD1S3AX integrator3_i55 (.D(integrator3_71__N_1104[55]), .CK(clk_80mhz), 
            .Q(integrator3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i55.GSR = "ENABLED";
    FD1S3AX integrator3_i54 (.D(integrator3_71__N_1104[54]), .CK(clk_80mhz), 
            .Q(integrator3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i54.GSR = "ENABLED";
    FD1S3AX integrator3_i53 (.D(integrator3_71__N_1104[53]), .CK(clk_80mhz), 
            .Q(integrator3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i53.GSR = "ENABLED";
    FD1S3AX integrator3_i52 (.D(integrator3_71__N_1104[52]), .CK(clk_80mhz), 
            .Q(integrator3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i52.GSR = "ENABLED";
    FD1S3AX integrator3_i51 (.D(integrator3_71__N_1104[51]), .CK(clk_80mhz), 
            .Q(integrator3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i51.GSR = "ENABLED";
    FD1S3AX integrator3_i50 (.D(integrator3_71__N_1104[50]), .CK(clk_80mhz), 
            .Q(integrator3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i50.GSR = "ENABLED";
    FD1S3AX integrator3_i49 (.D(integrator3_71__N_1104[49]), .CK(clk_80mhz), 
            .Q(integrator3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i49.GSR = "ENABLED";
    FD1S3AX integrator3_i48 (.D(integrator3_71__N_1104[48]), .CK(clk_80mhz), 
            .Q(integrator3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i48.GSR = "ENABLED";
    FD1S3AX integrator3_i47 (.D(integrator3_71__N_1104[47]), .CK(clk_80mhz), 
            .Q(integrator3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i47.GSR = "ENABLED";
    FD1S3AX integrator3_i46 (.D(integrator3_71__N_1104[46]), .CK(clk_80mhz), 
            .Q(integrator3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i46.GSR = "ENABLED";
    FD1S3AX integrator3_i45 (.D(integrator3_71__N_1104[45]), .CK(clk_80mhz), 
            .Q(integrator3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i45.GSR = "ENABLED";
    FD1S3AX integrator3_i44 (.D(integrator3_71__N_1104[44]), .CK(clk_80mhz), 
            .Q(integrator3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i44.GSR = "ENABLED";
    FD1S3AX integrator3_i43 (.D(integrator3_71__N_1104[43]), .CK(clk_80mhz), 
            .Q(integrator3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i43.GSR = "ENABLED";
    FD1S3AX integrator3_i42 (.D(integrator3_71__N_1104[42]), .CK(clk_80mhz), 
            .Q(integrator3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i42.GSR = "ENABLED";
    FD1S3AX integrator3_i41 (.D(integrator3_71__N_1104[41]), .CK(clk_80mhz), 
            .Q(integrator3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i41.GSR = "ENABLED";
    FD1S3AX integrator3_i40 (.D(integrator3_71__N_1104[40]), .CK(clk_80mhz), 
            .Q(integrator3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i40.GSR = "ENABLED";
    FD1S3AX integrator3_i39 (.D(integrator3_71__N_1104[39]), .CK(clk_80mhz), 
            .Q(integrator3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i39.GSR = "ENABLED";
    FD1S3AX integrator3_i38 (.D(integrator3_71__N_1104[38]), .CK(clk_80mhz), 
            .Q(integrator3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i38.GSR = "ENABLED";
    FD1S3AX integrator3_i37 (.D(integrator3_71__N_1104[37]), .CK(clk_80mhz), 
            .Q(integrator3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i37.GSR = "ENABLED";
    FD1S3AX integrator3_i36 (.D(integrator3_71__N_1104[36]), .CK(clk_80mhz), 
            .Q(integrator3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i36.GSR = "ENABLED";
    FD1S3AX integrator3_i35 (.D(integrator3_71__N_1104[35]), .CK(clk_80mhz), 
            .Q(integrator3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i35.GSR = "ENABLED";
    FD1S3AX integrator3_i34 (.D(integrator3_71__N_1104[34]), .CK(clk_80mhz), 
            .Q(integrator3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i34.GSR = "ENABLED";
    FD1S3AX integrator3_i33 (.D(integrator3_71__N_1104[33]), .CK(clk_80mhz), 
            .Q(integrator3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i33.GSR = "ENABLED";
    FD1S3AX integrator3_i32 (.D(integrator3_71__N_1104[32]), .CK(clk_80mhz), 
            .Q(integrator3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i32.GSR = "ENABLED";
    FD1S3AX integrator3_i31 (.D(integrator3_71__N_1104[31]), .CK(clk_80mhz), 
            .Q(integrator3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i31.GSR = "ENABLED";
    FD1S3AX integrator3_i30 (.D(integrator3_71__N_1104[30]), .CK(clk_80mhz), 
            .Q(integrator3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i30.GSR = "ENABLED";
    FD1S3AX integrator3_i29 (.D(integrator3_71__N_1104[29]), .CK(clk_80mhz), 
            .Q(integrator3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i29.GSR = "ENABLED";
    FD1S3AX integrator3_i28 (.D(integrator3_71__N_1104[28]), .CK(clk_80mhz), 
            .Q(integrator3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i28.GSR = "ENABLED";
    FD1S3AX integrator3_i27 (.D(integrator3_71__N_1104[27]), .CK(clk_80mhz), 
            .Q(integrator3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i27.GSR = "ENABLED";
    FD1S3AX integrator3_i26 (.D(integrator3_71__N_1104[26]), .CK(clk_80mhz), 
            .Q(integrator3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i26.GSR = "ENABLED";
    FD1S3AX integrator3_i25 (.D(integrator3_71__N_1104[25]), .CK(clk_80mhz), 
            .Q(integrator3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i25.GSR = "ENABLED";
    FD1S3AX integrator3_i24 (.D(integrator3_71__N_1104[24]), .CK(clk_80mhz), 
            .Q(integrator3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i24.GSR = "ENABLED";
    FD1S3AX integrator3_i23 (.D(integrator3_71__N_1104[23]), .CK(clk_80mhz), 
            .Q(integrator3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i23.GSR = "ENABLED";
    FD1S3AX integrator3_i22 (.D(integrator3_71__N_1104[22]), .CK(clk_80mhz), 
            .Q(integrator3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i22.GSR = "ENABLED";
    FD1S3AX integrator3_i21 (.D(integrator3_71__N_1104[21]), .CK(clk_80mhz), 
            .Q(integrator3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i21.GSR = "ENABLED";
    FD1S3AX integrator3_i20 (.D(integrator3_71__N_1104[20]), .CK(clk_80mhz), 
            .Q(integrator3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i20.GSR = "ENABLED";
    FD1S3AX integrator3_i19 (.D(integrator3_71__N_1104[19]), .CK(clk_80mhz), 
            .Q(integrator3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i19.GSR = "ENABLED";
    FD1S3AX integrator3_i18 (.D(integrator3_71__N_1104[18]), .CK(clk_80mhz), 
            .Q(integrator3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i18.GSR = "ENABLED";
    FD1S3AX integrator3_i17 (.D(integrator3_71__N_1104[17]), .CK(clk_80mhz), 
            .Q(integrator3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i17.GSR = "ENABLED";
    FD1S3AX integrator3_i16 (.D(integrator3_71__N_1104[16]), .CK(clk_80mhz), 
            .Q(integrator3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i16.GSR = "ENABLED";
    FD1S3AX integrator3_i15 (.D(integrator3_71__N_1104[15]), .CK(clk_80mhz), 
            .Q(integrator3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i15.GSR = "ENABLED";
    FD1S3AX integrator3_i14 (.D(integrator3_71__N_1104[14]), .CK(clk_80mhz), 
            .Q(integrator3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i14.GSR = "ENABLED";
    FD1S3AX integrator3_i13 (.D(integrator3_71__N_1104[13]), .CK(clk_80mhz), 
            .Q(integrator3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i13.GSR = "ENABLED";
    FD1S3AX integrator3_i12 (.D(integrator3_71__N_1104[12]), .CK(clk_80mhz), 
            .Q(integrator3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i12.GSR = "ENABLED";
    FD1S3AX integrator3_i11 (.D(integrator3_71__N_1104[11]), .CK(clk_80mhz), 
            .Q(integrator3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i11.GSR = "ENABLED";
    FD1S3AX integrator3_i10 (.D(integrator3_71__N_1104[10]), .CK(clk_80mhz), 
            .Q(integrator3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i10.GSR = "ENABLED";
    FD1S3AX integrator3_i9 (.D(integrator3_71__N_1104[9]), .CK(clk_80mhz), 
            .Q(integrator3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i9.GSR = "ENABLED";
    FD1S3AX integrator3_i8 (.D(integrator3_71__N_1104[8]), .CK(clk_80mhz), 
            .Q(integrator3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i8.GSR = "ENABLED";
    FD1S3AX integrator3_i7 (.D(integrator3_71__N_1104[7]), .CK(clk_80mhz), 
            .Q(integrator3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i7.GSR = "ENABLED";
    FD1S3AX integrator3_i6 (.D(integrator3_71__N_1104[6]), .CK(clk_80mhz), 
            .Q(integrator3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i6.GSR = "ENABLED";
    FD1S3AX integrator3_i5 (.D(integrator3_71__N_1104[5]), .CK(clk_80mhz), 
            .Q(integrator3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i5.GSR = "ENABLED";
    FD1S3AX integrator3_i4 (.D(integrator3_71__N_1104[4]), .CK(clk_80mhz), 
            .Q(integrator3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i4.GSR = "ENABLED";
    FD1S3AX integrator3_i3 (.D(integrator3_71__N_1104[3]), .CK(clk_80mhz), 
            .Q(integrator3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i3.GSR = "ENABLED";
    FD1S3AX integrator3_i2 (.D(integrator3_71__N_1104[2]), .CK(clk_80mhz), 
            .Q(integrator3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i2.GSR = "ENABLED";
    FD1S3AX integrator3_i1 (.D(integrator3_71__N_1104[1]), .CK(clk_80mhz), 
            .Q(integrator3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator3_i1.GSR = "ENABLED";
    FD1S3AX integrator2_i71 (.D(integrator2_71__N_1032[71]), .CK(clk_80mhz), 
            .Q(integrator2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i71.GSR = "ENABLED";
    FD1S3AX integrator2_i70 (.D(integrator2_71__N_1032[70]), .CK(clk_80mhz), 
            .Q(integrator2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i70.GSR = "ENABLED";
    FD1S3AX integrator2_i69 (.D(integrator2_71__N_1032[69]), .CK(clk_80mhz), 
            .Q(integrator2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i69.GSR = "ENABLED";
    FD1S3AX integrator2_i68 (.D(integrator2_71__N_1032[68]), .CK(clk_80mhz), 
            .Q(integrator2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i68.GSR = "ENABLED";
    FD1S3AX integrator2_i67 (.D(integrator2_71__N_1032[67]), .CK(clk_80mhz), 
            .Q(integrator2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i67.GSR = "ENABLED";
    FD1S3AX integrator2_i66 (.D(integrator2_71__N_1032[66]), .CK(clk_80mhz), 
            .Q(integrator2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i66.GSR = "ENABLED";
    FD1S3AX integrator2_i65 (.D(integrator2_71__N_1032[65]), .CK(clk_80mhz), 
            .Q(integrator2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i65.GSR = "ENABLED";
    FD1S3AX integrator2_i64 (.D(integrator2_71__N_1032[64]), .CK(clk_80mhz), 
            .Q(integrator2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i64.GSR = "ENABLED";
    FD1S3AX integrator2_i63 (.D(integrator2_71__N_1032[63]), .CK(clk_80mhz), 
            .Q(integrator2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i63.GSR = "ENABLED";
    FD1S3AX integrator2_i62 (.D(integrator2_71__N_1032[62]), .CK(clk_80mhz), 
            .Q(integrator2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i62.GSR = "ENABLED";
    FD1S3AX integrator2_i61 (.D(integrator2_71__N_1032[61]), .CK(clk_80mhz), 
            .Q(integrator2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i61.GSR = "ENABLED";
    FD1S3AX integrator2_i60 (.D(integrator2_71__N_1032[60]), .CK(clk_80mhz), 
            .Q(integrator2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i60.GSR = "ENABLED";
    FD1S3AX integrator2_i59 (.D(integrator2_71__N_1032[59]), .CK(clk_80mhz), 
            .Q(integrator2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i59.GSR = "ENABLED";
    FD1S3AX integrator2_i58 (.D(integrator2_71__N_1032[58]), .CK(clk_80mhz), 
            .Q(integrator2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i58.GSR = "ENABLED";
    FD1S3AX integrator2_i57 (.D(integrator2_71__N_1032[57]), .CK(clk_80mhz), 
            .Q(integrator2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i57.GSR = "ENABLED";
    FD1S3AX integrator2_i56 (.D(integrator2_71__N_1032[56]), .CK(clk_80mhz), 
            .Q(integrator2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i56.GSR = "ENABLED";
    FD1S3AX integrator2_i55 (.D(integrator2_71__N_1032[55]), .CK(clk_80mhz), 
            .Q(integrator2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i55.GSR = "ENABLED";
    FD1S3AX integrator2_i54 (.D(integrator2_71__N_1032[54]), .CK(clk_80mhz), 
            .Q(integrator2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i54.GSR = "ENABLED";
    FD1S3AX integrator2_i53 (.D(integrator2_71__N_1032[53]), .CK(clk_80mhz), 
            .Q(integrator2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i53.GSR = "ENABLED";
    FD1S3AX integrator2_i52 (.D(integrator2_71__N_1032[52]), .CK(clk_80mhz), 
            .Q(integrator2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i52.GSR = "ENABLED";
    FD1S3AX integrator2_i51 (.D(integrator2_71__N_1032[51]), .CK(clk_80mhz), 
            .Q(integrator2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i51.GSR = "ENABLED";
    FD1S3AX integrator2_i50 (.D(integrator2_71__N_1032[50]), .CK(clk_80mhz), 
            .Q(integrator2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i50.GSR = "ENABLED";
    FD1S3AX integrator2_i49 (.D(integrator2_71__N_1032[49]), .CK(clk_80mhz), 
            .Q(integrator2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i49.GSR = "ENABLED";
    FD1S3AX integrator2_i48 (.D(integrator2_71__N_1032[48]), .CK(clk_80mhz), 
            .Q(integrator2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i48.GSR = "ENABLED";
    FD1S3AX integrator2_i47 (.D(integrator2_71__N_1032[47]), .CK(clk_80mhz), 
            .Q(integrator2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i47.GSR = "ENABLED";
    FD1S3AX integrator2_i46 (.D(integrator2_71__N_1032[46]), .CK(clk_80mhz), 
            .Q(integrator2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i46.GSR = "ENABLED";
    FD1S3AX integrator2_i45 (.D(integrator2_71__N_1032[45]), .CK(clk_80mhz), 
            .Q(integrator2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i45.GSR = "ENABLED";
    FD1S3AX integrator2_i44 (.D(integrator2_71__N_1032[44]), .CK(clk_80mhz), 
            .Q(integrator2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i44.GSR = "ENABLED";
    FD1S3AX integrator2_i43 (.D(integrator2_71__N_1032[43]), .CK(clk_80mhz), 
            .Q(integrator2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i43.GSR = "ENABLED";
    FD1S3AX integrator2_i42 (.D(integrator2_71__N_1032[42]), .CK(clk_80mhz), 
            .Q(integrator2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i42.GSR = "ENABLED";
    FD1S3AX integrator2_i41 (.D(integrator2_71__N_1032[41]), .CK(clk_80mhz), 
            .Q(integrator2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i41.GSR = "ENABLED";
    FD1S3AX integrator2_i40 (.D(integrator2_71__N_1032[40]), .CK(clk_80mhz), 
            .Q(integrator2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i40.GSR = "ENABLED";
    FD1S3AX integrator2_i39 (.D(integrator2_71__N_1032[39]), .CK(clk_80mhz), 
            .Q(integrator2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i39.GSR = "ENABLED";
    FD1S3AX integrator2_i38 (.D(integrator2_71__N_1032[38]), .CK(clk_80mhz), 
            .Q(integrator2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i38.GSR = "ENABLED";
    FD1S3AX integrator2_i37 (.D(integrator2_71__N_1032[37]), .CK(clk_80mhz), 
            .Q(integrator2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i37.GSR = "ENABLED";
    FD1S3AX integrator2_i36 (.D(integrator2_71__N_1032[36]), .CK(clk_80mhz), 
            .Q(integrator2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i36.GSR = "ENABLED";
    FD1S3AX integrator2_i35 (.D(integrator2_71__N_1032[35]), .CK(clk_80mhz), 
            .Q(integrator2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i35.GSR = "ENABLED";
    FD1S3AX integrator2_i34 (.D(integrator2_71__N_1032[34]), .CK(clk_80mhz), 
            .Q(integrator2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i34.GSR = "ENABLED";
    FD1S3AX integrator2_i33 (.D(integrator2_71__N_1032[33]), .CK(clk_80mhz), 
            .Q(integrator2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i33.GSR = "ENABLED";
    FD1S3AX integrator2_i32 (.D(integrator2_71__N_1032[32]), .CK(clk_80mhz), 
            .Q(integrator2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i32.GSR = "ENABLED";
    FD1S3AX integrator2_i31 (.D(integrator2_71__N_1032[31]), .CK(clk_80mhz), 
            .Q(integrator2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i31.GSR = "ENABLED";
    FD1S3AX integrator2_i30 (.D(integrator2_71__N_1032[30]), .CK(clk_80mhz), 
            .Q(integrator2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i30.GSR = "ENABLED";
    FD1S3AX integrator2_i29 (.D(integrator2_71__N_1032[29]), .CK(clk_80mhz), 
            .Q(integrator2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i29.GSR = "ENABLED";
    FD1S3AX integrator2_i28 (.D(integrator2_71__N_1032[28]), .CK(clk_80mhz), 
            .Q(integrator2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i28.GSR = "ENABLED";
    FD1S3AX integrator2_i27 (.D(integrator2_71__N_1032[27]), .CK(clk_80mhz), 
            .Q(integrator2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i27.GSR = "ENABLED";
    FD1S3AX integrator2_i26 (.D(integrator2_71__N_1032[26]), .CK(clk_80mhz), 
            .Q(integrator2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i26.GSR = "ENABLED";
    FD1S3AX integrator2_i25 (.D(integrator2_71__N_1032[25]), .CK(clk_80mhz), 
            .Q(integrator2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i25.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i44_1_lut (.A(comb_d6[43]), .Z(n30_adj_28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i44_1_lut.init = 16'h5555;
    FD1S3AX integrator2_i24 (.D(integrator2_71__N_1032[24]), .CK(clk_80mhz), 
            .Q(integrator2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i24.GSR = "ENABLED";
    FD1S3AX integrator2_i23 (.D(integrator2_71__N_1032[23]), .CK(clk_80mhz), 
            .Q(integrator2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i23.GSR = "ENABLED";
    FD1S3AX integrator2_i22 (.D(integrator2_71__N_1032[22]), .CK(clk_80mhz), 
            .Q(integrator2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i22.GSR = "ENABLED";
    FD1S3AX integrator2_i21 (.D(integrator2_71__N_1032[21]), .CK(clk_80mhz), 
            .Q(integrator2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i21.GSR = "ENABLED";
    FD1S3AX integrator2_i20 (.D(integrator2_71__N_1032[20]), .CK(clk_80mhz), 
            .Q(integrator2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i20.GSR = "ENABLED";
    FD1S3AX integrator2_i19 (.D(integrator2_71__N_1032[19]), .CK(clk_80mhz), 
            .Q(integrator2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i19.GSR = "ENABLED";
    FD1S3AX integrator2_i18 (.D(integrator2_71__N_1032[18]), .CK(clk_80mhz), 
            .Q(integrator2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i18.GSR = "ENABLED";
    FD1S3AX integrator2_i17 (.D(integrator2_71__N_1032[17]), .CK(clk_80mhz), 
            .Q(integrator2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i17.GSR = "ENABLED";
    FD1S3AX integrator2_i16 (.D(integrator2_71__N_1032[16]), .CK(clk_80mhz), 
            .Q(integrator2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i16.GSR = "ENABLED";
    FD1S3AX integrator2_i15 (.D(integrator2_71__N_1032[15]), .CK(clk_80mhz), 
            .Q(integrator2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i15.GSR = "ENABLED";
    FD1S3AX integrator2_i14 (.D(integrator2_71__N_1032[14]), .CK(clk_80mhz), 
            .Q(integrator2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i14.GSR = "ENABLED";
    FD1S3AX integrator2_i13 (.D(integrator2_71__N_1032[13]), .CK(clk_80mhz), 
            .Q(integrator2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i13.GSR = "ENABLED";
    FD1S3AX integrator2_i12 (.D(integrator2_71__N_1032[12]), .CK(clk_80mhz), 
            .Q(integrator2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i12.GSR = "ENABLED";
    FD1S3AX integrator2_i11 (.D(integrator2_71__N_1032[11]), .CK(clk_80mhz), 
            .Q(integrator2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i11.GSR = "ENABLED";
    FD1S3AX integrator2_i10 (.D(integrator2_71__N_1032[10]), .CK(clk_80mhz), 
            .Q(integrator2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i10.GSR = "ENABLED";
    FD1S3AX integrator2_i9 (.D(integrator2_71__N_1032[9]), .CK(clk_80mhz), 
            .Q(integrator2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i9.GSR = "ENABLED";
    FD1S3AX integrator2_i8 (.D(integrator2_71__N_1032[8]), .CK(clk_80mhz), 
            .Q(integrator2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i8.GSR = "ENABLED";
    FD1S3AX integrator2_i7 (.D(integrator2_71__N_1032[7]), .CK(clk_80mhz), 
            .Q(integrator2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i7.GSR = "ENABLED";
    FD1S3AX integrator2_i6 (.D(integrator2_71__N_1032[6]), .CK(clk_80mhz), 
            .Q(integrator2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i6.GSR = "ENABLED";
    FD1S3AX integrator2_i5 (.D(integrator2_71__N_1032[5]), .CK(clk_80mhz), 
            .Q(integrator2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i5.GSR = "ENABLED";
    FD1S3AX integrator2_i4 (.D(integrator2_71__N_1032[4]), .CK(clk_80mhz), 
            .Q(integrator2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i4.GSR = "ENABLED";
    FD1S3AX integrator2_i3 (.D(integrator2_71__N_1032[3]), .CK(clk_80mhz), 
            .Q(integrator2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i3.GSR = "ENABLED";
    FD1S3AX integrator2_i2 (.D(integrator2_71__N_1032[2]), .CK(clk_80mhz), 
            .Q(integrator2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i2.GSR = "ENABLED";
    FD1S3AX integrator2_i1 (.D(integrator2_71__N_1032[1]), .CK(clk_80mhz), 
            .Q(integrator2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator2_i1.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i71 (.D(integrator_tmp[71]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i70 (.D(integrator_tmp[70]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i69 (.D(integrator_tmp[69]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i68 (.D(integrator_tmp[68]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i67 (.D(integrator_tmp[67]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i66 (.D(integrator_tmp[66]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i65 (.D(integrator_tmp[65]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i64 (.D(integrator_tmp[64]), .SP(clk_80mhz_enable_752), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i63 (.D(integrator_tmp[63]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i63.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i41_1_lut (.A(comb_d6[40]), .Z(n33_adj_29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i41_1_lut.init = 16'h5555;
    FD1P3AX integrator_d_tmp_i0_i62 (.D(integrator_tmp[62]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i61 (.D(integrator_tmp[61]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i60 (.D(integrator_tmp[60]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i59 (.D(integrator_tmp[59]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i58 (.D(integrator_tmp[58]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i57 (.D(integrator_tmp[57]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i56 (.D(integrator_tmp[56]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i55 (.D(integrator_tmp[55]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i54 (.D(integrator_tmp[54]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i53 (.D(integrator_tmp[53]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i52 (.D(integrator_tmp[52]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i51 (.D(integrator_tmp[51]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i50 (.D(integrator_tmp[50]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i49 (.D(integrator_tmp[49]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i48 (.D(integrator_tmp[48]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i47 (.D(integrator_tmp[47]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i46 (.D(integrator_tmp[46]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i45 (.D(integrator_tmp[45]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i45.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i42_1_lut (.A(comb_d6[41]), .Z(n32_adj_30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i39_1_lut (.A(comb_d6[38]), .Z(n35_adj_31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i39_1_lut.init = 16'h5555;
    FD1P3AX integrator_d_tmp_i0_i44 (.D(integrator_tmp[44]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i43 (.D(integrator_tmp[43]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i42 (.D(integrator_tmp[42]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i41 (.D(integrator_tmp[41]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i40 (.D(integrator_tmp[40]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i39 (.D(integrator_tmp[39]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i38 (.D(integrator_tmp[38]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i37 (.D(integrator_tmp[37]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i36 (.D(integrator_tmp[36]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i35 (.D(integrator_tmp[35]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i34 (.D(integrator_tmp[34]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i33 (.D(integrator_tmp[33]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i32 (.D(integrator_tmp[32]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i31 (.D(integrator_tmp[31]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i30 (.D(integrator_tmp[30]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i29 (.D(integrator_tmp[29]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i29.GSR = "ENABLED";
    LUT4 sub_29_inv_0_i65_1_lut (.A(comb_d8[64]), .Z(n9_adj_32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i65_1_lut.init = 16'h5555;
    FD1P3AX integrator_d_tmp_i0_i28 (.D(integrator_tmp[28]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i28.GSR = "ENABLED";
    LUT4 sub_29_inv_0_i66_1_lut (.A(comb_d8[65]), .Z(n8_adj_33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i66_1_lut.init = 16'h5555;
    FD1P3AX integrator_d_tmp_i0_i27 (.D(integrator_tmp[27]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i26 (.D(integrator_tmp[26]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i25 (.D(integrator_tmp[25]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i24 (.D(integrator_tmp[24]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i23 (.D(integrator_tmp[23]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i22 (.D(integrator_tmp[22]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i21 (.D(integrator_tmp[21]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i20 (.D(integrator_tmp[20]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i19 (.D(integrator_tmp[19]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i18 (.D(integrator_tmp[18]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i17 (.D(integrator_tmp[17]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i16 (.D(integrator_tmp[16]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i15 (.D(integrator_tmp[15]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i14 (.D(integrator_tmp[14]), .SP(clk_80mhz_enable_802), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i13 (.D(integrator_tmp[13]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i12 (.D(integrator_tmp[12]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i11 (.D(integrator_tmp[11]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i10 (.D(integrator_tmp[10]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i9 (.D(integrator_tmp[9]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i8 (.D(integrator_tmp[8]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i7 (.D(integrator_tmp[7]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i6 (.D(integrator_tmp[6]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i5 (.D(integrator_tmp[5]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i4 (.D(integrator_tmp[4]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i3 (.D(integrator_tmp[3]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i2 (.D(integrator_tmp[2]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i1 (.D(integrator_tmp[1]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(101[10] 116[6])
    defparam integrator_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i71 (.D(integrator5[71]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i70 (.D(integrator5[70]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i69 (.D(integrator5[69]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i68 (.D(integrator5[68]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i67 (.D(integrator5[67]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i66 (.D(integrator5[66]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i65 (.D(integrator5[65]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i64 (.D(integrator5[64]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i63 (.D(integrator5[63]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i62 (.D(integrator5[62]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i61 (.D(integrator5[61]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i60 (.D(integrator5[60]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i59 (.D(integrator5[59]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i58 (.D(integrator5[58]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i57 (.D(integrator5[57]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i56 (.D(integrator5[56]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i55 (.D(integrator5[55]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i54 (.D(integrator5[54]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i53 (.D(integrator5[53]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i52 (.D(integrator5[52]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i51 (.D(integrator5[51]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i50 (.D(integrator5[50]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i49 (.D(integrator5[49]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i48 (.D(integrator5[48]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i47 (.D(integrator5[47]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i46 (.D(integrator5[46]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i45 (.D(integrator5[45]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i44 (.D(integrator5[44]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i43 (.D(integrator5[43]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i42 (.D(integrator5[42]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i41 (.D(integrator5[41]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i40 (.D(integrator5[40]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i39 (.D(integrator5[39]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i38 (.D(integrator5[38]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i37 (.D(integrator5[37]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i36 (.D(integrator5[36]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i35 (.D(integrator5[35]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i34 (.D(integrator5[34]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i33 (.D(integrator5[33]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i32 (.D(integrator5[32]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i31 (.D(integrator5[31]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i30 (.D(integrator5[30]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i29 (.D(integrator5[29]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i28 (.D(integrator5[28]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i27 (.D(integrator5[27]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i26 (.D(integrator5[26]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i25 (.D(integrator5[25]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i24 (.D(integrator5[24]), .SP(clk_80mhz_enable_850), 
            .CK(clk_80mhz), .Q(integrator_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i23 (.D(integrator5[23]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i23.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i40_1_lut (.A(comb_d6[39]), .Z(n34_adj_34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i40_1_lut.init = 16'h5555;
    FD1P3AX integrator_tmp_i0_i22 (.D(integrator5[22]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i21 (.D(integrator5[21]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i20 (.D(integrator5[20]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i19 (.D(integrator5[19]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i18 (.D(integrator5[18]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i17 (.D(integrator5[17]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i16 (.D(integrator5[16]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i15 (.D(integrator5[15]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i14 (.D(integrator5[14]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i13 (.D(integrator5[13]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i12 (.D(integrator5[12]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i11 (.D(integrator5[11]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i10 (.D(integrator5[10]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i9 (.D(integrator5[9]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i8 (.D(integrator5[8]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i7 (.D(integrator5[7]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i6 (.D(integrator5[6]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i5 (.D(integrator5[5]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i4 (.D(integrator5[4]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i3 (.D(integrator5[3]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i2 (.D(integrator5[2]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i1 (.D(integrator5[1]), .SP(count_11__N_1992), 
            .CK(clk_80mhz), .Q(integrator_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam integrator_tmp_i0_i1.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i37_1_lut (.A(comb_d6[36]), .Z(n37_adj_35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i38_1_lut (.A(comb_d6[37]), .Z(n36_adj_36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(108[28:43])
    defparam sub_27_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i71_1_lut (.A(comb_d7[70]), .Z(n3_adj_37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i72_1_lut (.A(comb_d7[71]), .Z(n2_adj_38)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i63_1_lut (.A(comb_d8[62]), .Z(n11_adj_39)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i69_1_lut (.A(comb_d7[68]), .Z(n5_adj_40)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i70_1_lut (.A(comb_d7[69]), .Z(n4_adj_41)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i67_1_lut (.A(comb_d7[66]), .Z(n7_adj_42)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i68_1_lut (.A(comb_d7[67]), .Z(n6_adj_43)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i64_1_lut (.A(comb_d8[63]), .Z(n10_adj_44)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i65_1_lut (.A(comb_d7[64]), .Z(n9_adj_45)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i66_1_lut (.A(comb_d7[65]), .Z(n8_adj_46)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i63_1_lut (.A(comb_d7[62]), .Z(n11_adj_47)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i64_1_lut (.A(comb_d7[63]), .Z(n10_adj_48)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i61_1_lut (.A(comb_d7[60]), .Z(n13_adj_49)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i62_1_lut (.A(comb_d7[61]), .Z(n12_adj_50)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i59_1_lut (.A(comb_d7[58]), .Z(n15_adj_51)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i61_1_lut (.A(comb_d8[60]), .Z(n13_adj_52)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i60_1_lut (.A(comb_d7[59]), .Z(n14_adj_53)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i57_1_lut (.A(comb_d7[56]), .Z(n17_adj_54)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i58_1_lut (.A(comb_d7[57]), .Z(n16_adj_55)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i55_1_lut (.A(comb_d7[54]), .Z(n19_adj_56)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i62_1_lut (.A(comb_d8[61]), .Z(n12_adj_57)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i56_1_lut (.A(comb_d7[55]), .Z(n18_adj_58)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i59_1_lut (.A(comb_d8[58]), .Z(n15_adj_59)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i53_1_lut (.A(comb_d7[52]), .Z(n21_adj_60)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i53_1_lut.init = 16'h5555;
    FD1S3IX count__i0 (.D(count_11__N_1980[0]), .CK(clk_80mhz), .CD(count_11__N_1992), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i0.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i54_1_lut (.A(comb_d7[53]), .Z(n20_adj_61)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i51_1_lut (.A(comb_d7[50]), .Z(n23_adj_62)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i52_1_lut (.A(comb_d7[51]), .Z(n22_adj_63)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i49_1_lut (.A(comb_d7[48]), .Z(n25_adj_64)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i50_1_lut (.A(comb_d7[49]), .Z(n24_adj_65)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i47_1_lut (.A(comb_d7[46]), .Z(n27_adj_66)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i48_1_lut (.A(comb_d7[47]), .Z(n26_adj_67)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i45_1_lut (.A(comb_d7[44]), .Z(n29_adj_68)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i46_1_lut (.A(comb_d7[45]), .Z(n28_adj_69)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i43_1_lut (.A(comb_d7[42]), .Z(n31_adj_70)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i44_1_lut (.A(comb_d7[43]), .Z(n30_adj_71)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 i1_4_lut (.A(n18778), .B(count[6]), .C(n18762), .D(count[8]), 
         .Z(count_11__N_1992)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_186 (.A(count[2]), .B(n18774), .C(n18760), .D(count[4]), 
         .Z(n18778)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_186.init = 16'h8000;
    LUT4 i1_2_lut (.A(count[11]), .B(count[9]), .Z(n18762)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_187 (.A(count[1]), .B(count[3]), .C(count[0]), .D(count[10]), 
         .Z(n18774)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_187.init = 16'h8000;
    LUT4 sub_26_inv_0_i65_1_lut (.A(integrator_d_tmp[64]), .Z(n9_adj_72)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_adj_188 (.A(count[7]), .B(count[5]), .Z(n18760)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_188.init = 16'h8888;
    LUT4 sub_26_inv_0_i66_1_lut (.A(integrator_d_tmp[65]), .Z(n8_adj_73)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i41_1_lut (.A(comb_d7[40]), .Z(n33_adj_74)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i63_1_lut (.A(integrator_d_tmp[62]), .Z(n11_adj_75)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i64_1_lut (.A(integrator_d_tmp[63]), .Z(n10_adj_76)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i42_1_lut (.A(comb_d7[41]), .Z(n32_adj_77)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i39_1_lut (.A(comb_d7[38]), .Z(n35_adj_78)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 comb10_71__I_0_77_i70_3_lut (.A(\comb10[69] ), .B(\comb10[70] ), 
         .C(\cic_gain[0] ), .Z(n70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i70_3_lut.init = 16'hcaca;
    LUT4 comb10_71__I_0_77_i68_3_lut (.A(\comb10[67] ), .B(\comb10[68] ), 
         .C(\cic_gain[0] ), .Z(n68)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i68_3_lut.init = 16'hcaca;
    LUT4 comb10_71__I_0_77_i67_3_lut (.A(\comb10[66] ), .B(\comb10[67] ), 
         .C(\cic_gain[0] ), .Z(n67)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i67_3_lut.init = 16'hcaca;
    LUT4 comb10_71__I_0_77_i66_3_lut (.A(\comb10[65] ), .B(\comb10[66] ), 
         .C(\cic_gain[0] ), .Z(n66)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i66_3_lut.init = 16'hcaca;
    LUT4 comb10_71__I_0_77_i65_3_lut (.A(\comb10[64] ), .B(\comb10[65] ), 
         .C(\cic_gain[0] ), .Z(n65)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i65_3_lut.init = 16'hcaca;
    LUT4 comb10_71__I_0_77_i64_3_lut (.A(\comb10[63] ), .B(\comb10[64] ), 
         .C(\cic_gain[0] ), .Z(n64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i64_3_lut.init = 16'hcaca;
    LUT4 comb10_71__I_0_77_i63_3_lut (.A(\comb10[62] ), .B(\comb10[63] ), 
         .C(\cic_gain[0] ), .Z(n63)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i63_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i40_1_lut (.A(comb_d7[39]), .Z(n34_adj_79)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i37_1_lut (.A(comb_d7[36]), .Z(n37_adj_80)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i38_1_lut (.A(comb_d7[37]), .Z(n36_adj_81)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(110[28:43])
    defparam sub_28_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i61_1_lut (.A(integrator_d_tmp[60]), .Z(n13_adj_82)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i62_1_lut (.A(integrator_d_tmp[61]), .Z(n12_adj_83)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i60_1_lut (.A(comb_d8[59]), .Z(n14_adj_84)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i59_1_lut (.A(integrator_d_tmp[58]), .Z(n15_adj_85)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i57_1_lut (.A(comb_d8[56]), .Z(n17_adj_86)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 i8378_2_lut (.A(n23_c), .B(n20267), .Z(n14290)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam i8378_2_lut.init = 16'hdddd;
    LUT4 sub_29_inv_0_i58_1_lut (.A(comb_d8[57]), .Z(n16_adj_87)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i60_1_lut (.A(integrator_d_tmp[59]), .Z(n14_adj_88)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i55_1_lut (.A(comb_d8[54]), .Z(n19_adj_89)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i56_1_lut (.A(comb_d8[55]), .Z(n18_adj_90)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i53_1_lut (.A(comb_d8[52]), .Z(n21_adj_91)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i54_1_lut (.A(comb_d8[53]), .Z(n20_adj_92)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 comb10_71__I_0_77_i61_3_lut (.A(\comb10[60] ), .B(\comb10[61] ), 
         .C(\cic_gain[0] ), .Z(n61_adj_93)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(118[21:70])
    defparam comb10_71__I_0_77_i61_3_lut.init = 16'hcaca;
    LUT4 sub_29_inv_0_i51_1_lut (.A(comb_d8[50]), .Z(n23_adj_94)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i52_1_lut (.A(comb_d8[51]), .Z(n22_adj_95)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i49_1_lut (.A(comb_d8[48]), .Z(n25_adj_96)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i57_1_lut (.A(integrator_d_tmp[56]), .Z(n17_adj_97)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i58_1_lut (.A(integrator_d_tmp[57]), .Z(n16_adj_98)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i50_1_lut (.A(comb_d8[49]), .Z(n24_adj_99)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i47_1_lut (.A(comb_d8[46]), .Z(n27_adj_100)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i48_1_lut (.A(comb_d8[47]), .Z(n26_adj_101)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 mux_3409_i16_3_lut (.A(n76), .B(n78), .C(cout), .Z(comb10_71__N_2281[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i16_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i15_3_lut (.A(n79), .B(n81), .C(cout), .Z(comb10_71__N_2281[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i15_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i14_3_lut (.A(n82), .B(n84), .C(cout), .Z(comb10_71__N_2281[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i14_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i13_3_lut (.A(n85), .B(n87), .C(cout), .Z(comb10_71__N_2281[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i13_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i12_3_lut (.A(n88), .B(n90), .C(cout), .Z(comb10_71__N_2281[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i12_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i11_3_lut (.A(n91), .B(n93), .C(cout), .Z(comb10_71__N_2281[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i11_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i10_3_lut (.A(n94), .B(n96), .C(cout), .Z(comb10_71__N_2281[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i10_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i9_3_lut (.A(n97), .B(n99), .C(cout), .Z(comb10_71__N_2281[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i9_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i8_3_lut (.A(n100), .B(n102), .C(cout), .Z(comb10_71__N_2281[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i8_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i7_3_lut (.A(n103), .B(n105), .C(cout), .Z(comb10_71__N_2281[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i7_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i6_3_lut (.A(n106), .B(n108), .C(cout), .Z(comb10_71__N_2281[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i6_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i5_3_lut (.A(n109), .B(n111), .C(cout), .Z(comb10_71__N_2281[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i5_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i4_3_lut (.A(n112), .B(n114), .C(cout), .Z(comb10_71__N_2281[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i3_3_lut (.A(n115), .B(n117), .C(cout), .Z(comb10_71__N_2281[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i3_3_lut.init = 16'hcaca;
    LUT4 mux_3409_i2_3_lut (.A(n118), .B(n120), .C(cout), .Z(comb10_71__N_2281[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(114[28:43])
    defparam mux_3409_i2_3_lut.init = 16'hcaca;
    LUT4 sub_29_inv_0_i45_1_lut (.A(comb_d8[44]), .Z(n29_adj_102)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i46_1_lut (.A(comb_d8[45]), .Z(n28_adj_103)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i72_1_lut (.A(integrator_d_tmp[71]), .Z(n2_adj_104)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i71_1_lut (.A(integrator_d_tmp[70]), .Z(n3_adj_105)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(106[28:61])
    defparam sub_26_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i43_1_lut (.A(comb_d8[42]), .Z(n31_adj_106)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i44_1_lut (.A(comb_d8[43]), .Z(n30_adj_107)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i41_1_lut (.A(comb_d8[40]), .Z(n33_adj_108)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i42_1_lut (.A(comb_d8[41]), .Z(n32_adj_109)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i39_1_lut (.A(comb_d8[38]), .Z(n35_adj_110)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i40_1_lut (.A(comb_d8[39]), .Z(n34_adj_111)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 i4858_2_lut (.A(n67_adj_114[0]), .B(n23_c), .Z(count_11__N_1980[0])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(92[14] 95[8])
    defparam i4858_2_lut.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_189 (.A(count[11]), .B(n18816), .C(n18800), .D(n18808), 
         .Z(n23_c)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(88[18:48])
    defparam i1_4_lut_adj_189.init = 16'hfffd;
    LUT4 i1_4_lut_adj_190 (.A(count[6]), .B(n18812), .C(count[7]), .D(count[4]), 
         .Z(n18816)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(88[18:48])
    defparam i1_4_lut_adj_190.init = 16'hfffe;
    LUT4 i1_2_lut_adj_191 (.A(count[2]), .B(count[5]), .Z(n18800)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(88[18:48])
    defparam i1_2_lut_adj_191.init = 16'heeee;
    LUT4 i1_2_lut_adj_192 (.A(count[9]), .B(count[10]), .Z(n18808)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(88[18:48])
    defparam i1_2_lut_adj_192.init = 16'heeee;
    LUT4 i1_4_lut_adj_193 (.A(count[1]), .B(count[3]), .C(count[0]), .D(count[8]), 
         .Z(n18812)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(88[18:48])
    defparam i1_4_lut_adj_193.init = 16'hfffe;
    LUT4 sub_29_inv_0_i37_1_lut (.A(comb_d8[36]), .Z(n37_adj_112)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_29_inv_0_i38_1_lut (.A(comb_d8[37]), .Z(n36_adj_113)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(112[28:43])
    defparam sub_29_inv_0_i38_1_lut.init = 16'h5555;
    FD1S3IX count__i2 (.D(n67_adj_114[2]), .CK(clk_80mhz), .CD(n14290), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n67_adj_114[3]), .CK(clk_80mhz), .CD(n14290), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n67_adj_114[4]), .CK(clk_80mhz), .CD(n14290), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n67_adj_114[5]), .CK(clk_80mhz), .CD(n14290), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n67_adj_114[6]), .CK(clk_80mhz), .CD(n14290), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n67_adj_114[7]), .CK(clk_80mhz), .CD(n14290), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n67_adj_114[8]), .CK(clk_80mhz), .CD(n14290), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n67_adj_114[9]), .CK(clk_80mhz), .CD(n14290), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n67_adj_114[10]), .CK(clk_80mhz), .CD(n14290), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_11__N_1980[11]), .CK(clk_80mhz), .CD(count_11__N_1992), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i11.GSR = "ENABLED";
    LUT4 i8510_then_3_lut (.A(\cic_gain[1] ), .B(\comb10[59] ), .C(comb10[57]), 
         .Z(n19854)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i8510_then_3_lut.init = 16'he4e4;
    LUT4 i8510_else_3_lut (.A(n61_adj_93), .B(\cic_gain[1] ), .C(comb10[58]), 
         .Z(n19853)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i8510_else_3_lut.init = 16'he2e2;
    LUT4 i1_4_lut_rep_309 (.A(n18778), .B(count[6]), .C(n18762), .D(count[8]), 
         .Z(n20267)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_rep_309.init = 16'h8000;
    LUT4 i1_4_lut_rep_310 (.A(n18778), .B(count[6]), .C(n18762), .D(count[8]), 
         .Z(clk_80mhz_enable_850)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_rep_310.init = 16'h8000;
    FD1S3AX valid_comb_63_rep_324 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_802)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_324.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_323 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_752)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_323.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_322 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_702)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_322.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_321 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_652)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_321.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_320 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_600)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_320.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_319 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_550)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_319.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_318 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_499)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_318.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_317 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_449)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_317.GSR = "ENABLED";
    PFUMX i8769 (.BLUT(n19865), .ALUT(n19866), .C0(\cic_gain[0] ), .Z(\cic_cosine_out[1] ));
    FD1S3AX valid_comb_63_rep_316 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_394)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_316.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_315 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_341)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_315.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_314 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_195)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_314.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_313 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_136)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_313.GSR = "ENABLED";
    FD1S3AX valid_comb_63_rep_312 (.D(clk_80mhz_enable_850), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_71)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam valid_comb_63_rep_312.GSR = "ENABLED";
    PFUMX i8761 (.BLUT(n19853), .ALUT(n19854), .C0(\cic_gain[0] ), .Z(\cic_cosine_out[0] ));
    FD1S3IX count__i1 (.D(n67_adj_114[1]), .CK(clk_80mhz), .CD(n14290), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=206, LSE_RLINE=212 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version0-modified/impl1/source/CIC.v(71[10] 96[6])
    defparam count__i1.GSR = "ENABLED";
    
endmodule
