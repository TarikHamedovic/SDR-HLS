module cic#(
 parameter int IW = 5,
 parameter int OW = 10,
 parameter int R = 100,
 parameter int M = 10
)(
 input logic i_clk,
 input logic i_rest,
 input logic i_ce,
 input logic signed [IW-1:0 ]
)


endmodule