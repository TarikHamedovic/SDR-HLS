// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.13.0.56.2
// Netlist written on Sun Aug 25 17:35:18 2024
//
// Verilog Description of module top
//

module top (clk_25mhz, i_Rx_Serial, RFIn, o_Tx_Serial, led, XOut, 
            DiffOut, PWMOut, PWMOutP1, PWMOutP2, PWMOutP3, PWMOutP4, 
            PWMOutN1, PWMOutN2, PWMOutN3, PWMOutN4, sinGen, sin_out, 
            CIC_out_clkSin) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(39[8:11])
    input clk_25mhz;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(40[22:31])
    input i_Rx_Serial;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(41[22:33])
    input RFIn;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(42[22:26])
    output o_Tx_Serial;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(43[22:33])
    output [7:0]led;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(44[22:25])
    output XOut;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(45[22:26])
    output DiffOut;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(46[22:29])
    output PWMOut;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(47[22:28])
    output PWMOutP1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(48[22:30])
    output PWMOutP2;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(49[22:30])
    output PWMOutP3;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(50[22:30])
    output PWMOutP4;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(51[22:30])
    output PWMOutN1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(52[22:30])
    output PWMOutN2;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(53[22:30])
    output PWMOutN3;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(54[22:30])
    output PWMOutN4;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(55[22:30])
    output sinGen;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(56[22:28])
    output sin_out;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(57[22:29])
    output CIC_out_clkSin;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(58[22:36])
    
    wire clk_25mhz_c /* synthesis is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(40[22:31])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(61[23:32])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(74[23:38])
    
    wire GND_net, VCC_net, i_Rx_Serial_c, RFIn_c, led_c_7, led_c_6, 
        led_c_5, led_c_4, led_c_3, led_c_2, led_c_1, led_c_0, DiffOut_c, 
        PWMOutP4_c, PWMOutN4_c, sinGen_c, o_Rx_DV, o_Rx_DV1;
    wire [7:0]o_Rx_Byte1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(67[23:33])
    wire [11:0]MixerOutSin;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(70[23:34])
    wire [11:0]MixerOutCos;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(71[23:34])
    wire [11:0]CIC1_outCos;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(76[23:34])
    wire [63:0]phase_accum;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(78[23:34])
    wire [12:0]LOSine;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(79[23:29])
    wire [12:0]LOCosine;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(80[23:31])
    wire [63:0]phase_inc_carrGen;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(82[23:40])
    wire [63:0]phase_inc_carrGen1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(83[23:41])
    wire [11:0]DemodOut;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(85[23:31])
    wire [7:0]CICGain;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(86[23:30])
    
    wire n12609, n12611, n16114, n37, n36, n35, n34, n33, n32, 
        n31, n30, n29, n28, n27, n26, n25, n24, n23, n22, 
        n21, n20, n19, n18, n17, n16, n15, n14, n13, n12, 
        n11, n10, n9, n8, n7, n6, n5, n4, n3, n2, n16251, 
        n16250, n16249, n16438, n16437, n15_adj_2794, n60, n57, 
        n54, n51, n48, n45, n42, n39, n36_adj_2795, n33_adj_2796, 
        cout, n16436, n16435, n3901, n16434;
    wire [63:0]phase_accum_adj_5702;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(26[28:39])
    
    wire n12252, n26_adj_2797, n16433;
    wire [11:0]MixerOutSin_11__N_236;
    wire [11:0]MixerOutCos_11__N_250;
    
    wire n25_adj_2798;
    wire [71:0]d_tmp;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(52[28:33])
    wire [71:0]d_d_tmp;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(52[35:42])
    wire [71:0]d1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(53[28:30])
    wire [71:0]d2;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(53[32:34])
    wire [71:0]d3;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(53[36:38])
    wire [71:0]d4;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(53[40:42])
    wire [71:0]d5;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(53[44:46])
    wire [71:0]d6;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[28:30])
    wire [71:0]d_d6;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[32:36])
    wire [71:0]d7;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[38:40])
    wire [71:0]d_d7;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[42:46])
    wire [71:0]d8;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[48:50])
    wire [71:0]d_d8;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[52:56])
    wire [71:0]d9;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[58:60])
    wire [71:0]d_d9;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[62:66])
    
    wire n16113, n16112;
    wire [15:0]count;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(56[28:33])
    wire [71:0]d1_71__N_418;
    wire [71:0]d2_71__N_490;
    wire [71:0]d3_71__N_562;
    wire [71:0]d4_71__N_634;
    wire [71:0]d5_71__N_706;
    
    wire n16432, n16431, n16430, n16429, n16428, n16427, n16426, 
        n16425, n16424, n16423, n16422, n16421, n16420, n16419, 
        n81, n78, n75, n72, n69, n66, n63, n60_adj_2799, n57_adj_2800, 
        n54_adj_2801, n51_adj_2802, n48_adj_2803, n45_adj_2804, n42_adj_2805;
    wire [71:0]d6_71__N_1459;
    wire [71:0]d7_71__N_1531;
    wire [71:0]d8_71__N_1603;
    wire [71:0]d9_71__N_1675;
    
    wire n39_adj_2806, n36_adj_2807, cout_adj_2808, n16083, n16082, 
        n16081, n16080, n16079, n16078, n16077, n16076, n16075, 
        n16074, n16073, n16072, n16071, n16070, n16069, n16068, 
        n16067, n16066, n16061, n16060, n16059, n16058, n16057, 
        n16056, n16055, n16054, n16053, n16052, n16051, n16050, 
        n16049, cout_adj_2809, cout_adj_2810;
    wire [71:0]d_tmp_adj_5708;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(52[28:33])
    wire [71:0]d_d_tmp_adj_5709;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(52[35:42])
    wire [71:0]d1_adj_5710;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(53[28:30])
    wire [71:0]d2_adj_5711;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(53[32:34])
    wire [71:0]d3_adj_5712;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(53[36:38])
    wire [71:0]d4_adj_5713;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(53[40:42])
    wire [71:0]d5_adj_5714;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(53[44:46])
    wire [71:0]d6_adj_5715;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[28:30])
    wire [71:0]d_d6_adj_5716;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[32:36])
    wire [71:0]d7_adj_5717;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[38:40])
    wire [71:0]d_d7_adj_5718;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[42:46])
    wire [71:0]d8_adj_5719;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[48:50])
    wire [71:0]d_d8_adj_5720;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[52:56])
    wire [71:0]d9_adj_5721;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[58:60])
    wire [71:0]d_d9_adj_5722;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[62:66])
    wire [71:0]d10_adj_5723;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[68:71])
    
    wire n17523;
    wire [15:0]count_adj_5725;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(56[28:33])
    wire [71:0]d1_71__N_418_adj_5726;
    wire [71:0]d2_71__N_490_adj_5727;
    wire [71:0]d3_71__N_562_adj_5728;
    wire [71:0]d4_71__N_634_adj_5729;
    wire [71:0]d5_71__N_706_adj_5730;
    
    wire n16418, n16417, n16416, n16415, n16414, n16413, n16412, 
        n16411, n16410, n16409, n16408, n16407, cout_adj_4267;
    wire [71:0]d6_71__N_1459_adj_5742;
    wire [71:0]d7_71__N_1531_adj_5743;
    wire [71:0]d8_71__N_1603_adj_5744;
    wire [71:0]d9_71__N_1675_adj_5745;
    
    wire n16048, n16047, n16046, n16045, n16044, n16040, n16039, 
        n16038, n16037, n16036, n16035, n16034, n16033, n16032, 
        n16031, n16030, n16029, n16028, n16027, n16026, n16025, 
        n16024, n16023, n16022, n16021, n16020, n16019, n16018, 
        n24_adj_4556, n23_adj_4557, cout_adj_4558;
    wire [71:0]d_out_11__N_1819_adj_5748;
    
    wire n120, n117, n114, n111, n108, n105, n102, n99, n96, 
        n93, n90, n87, n84, n81_adj_4559, n78_adj_4560, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, 
        n153, n150, n147, n144, n141, n138, n135, n132, n129, 
        n126, n123, n120_adj_4561, n117_adj_4562, n114_adj_4563, n111_adj_4564, 
        n108_adj_4565, n105_adj_4566, n102_adj_4567, n99_adj_4568, n96_adj_4569, 
        n93_adj_4570, n90_adj_4571, n87_adj_4572, n84_adj_4573, n81_adj_4574, 
        n78_adj_4575, n22_adj_4576;
    wire [9:0]counter;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(36[12:19])
    wire [11:0]DataInReg;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(39[12:21])
    wire [11:0]DataInReg_11__N_1856;
    
    wire n16017, n16016;
    wire [31:0]ISquare;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(33[28:35])
    wire [11:0]MultDataB;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(38[28:37])
    wire [23:0]MultResult1;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(39[28:39])
    wire [23:0]MultResult2;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(43[28:39])
    
    wire n21_adj_4577, n20_adj_4578, n19_adj_4579, n18_adj_4580, n37_adj_4581, 
        n36_adj_4582, n35_adj_4583, n34_adj_4584, n33_adj_4585, n32_adj_4586, 
        n31_adj_4587, n30_adj_4588, n29_adj_4589, n28_adj_4590, n27_adj_4591, 
        n26_adj_4592, n25_adj_4593, n16248, n213, n24_adj_4594, n17_adj_4595, 
        n23_adj_4596, n22_adj_4597, n21_adj_4598, n20_adj_4599, n19_adj_4600, 
        n18_adj_4601, n17_adj_4602, n16_adj_4603, n15_adj_4604, n14_adj_4605, 
        n13_adj_4606, n12_adj_4607, n11_adj_4608, n10_adj_4609, n9_adj_4610, 
        n8_adj_4611, n7_adj_4612, n6_adj_4613, n5_adj_4614, n4_adj_4615, 
        n3_adj_4616, n2_adj_4617, n37_adj_4618, n36_adj_4619, n35_adj_4620, 
        n34_adj_4621, n33_adj_4622, n32_adj_4623, n31_adj_4624, n30_adj_4625, 
        n29_adj_4626, n28_adj_4627, n27_adj_4628, n26_adj_4629, n25_adj_4630, 
        n24_adj_4631, n23_adj_4632, n22_adj_4633, n21_adj_4634, n20_adj_4635, 
        n19_adj_4636, n18_adj_4637, n17_adj_4638, n16_adj_4639, n15_adj_4640, 
        n14_adj_4641, n13_adj_4642, n12_adj_4643, n11_adj_4644, n10_adj_4645, 
        n9_adj_4646, n8_adj_4647, n7_adj_4648, n6_adj_4649, n5_adj_4650, 
        n4_adj_4651, n3_adj_4652, n2_adj_4653, n16247;
    wire [17:0]d_out_d_11__N_1874;
    
    wire d_out_d_11__N_1873, n37_adj_4654, n36_adj_4655, n35_adj_4656;
    wire [17:0]d_out_d_11__N_1876;
    
    wire d_out_d_11__N_1875, n34_adj_4657, n33_adj_4658, n32_adj_4659, 
        n31_adj_4660, n30_adj_4661, n29_adj_4662, n28_adj_4663, n27_adj_4664, 
        n26_adj_4665, n25_adj_4666, n24_adj_4667, n23_adj_4668, n22_adj_4669, 
        n21_adj_4670, n20_adj_4671, n19_adj_4672, n18_adj_4673, n17_adj_4674, 
        n16_adj_4675, n15_adj_4676, n14_adj_4677, n13_adj_4678, n12_adj_4679, 
        n11_adj_4680, n10_adj_4681, n9_adj_4682, n8_adj_4683, n7_adj_4684, 
        n6_adj_4685, n5_adj_4686, n4_adj_4687, n3_adj_4688, n2_adj_4689;
    wire [17:0]d_out_d_11__N_1878;
    
    wire d_out_d_11__N_1877;
    wire [17:0]d_out_d_11__N_1880;
    
    wire d_out_d_11__N_1879, n37_adj_4690, n36_adj_4691, n35_adj_4692, 
        n34_adj_4693, n33_adj_4694, n32_adj_4695, n31_adj_4696, n30_adj_4697, 
        n29_adj_4698, n28_adj_4699, n27_adj_4700, n26_adj_4701, n25_adj_4702, 
        n24_adj_4703, n23_adj_4704, n22_adj_4705, n21_adj_4706, n20_adj_4707, 
        n19_adj_4708, n18_adj_4709, n17_adj_4710, n16_adj_4711, n15_adj_4712, 
        n14_adj_4713, n13_adj_4714, n12_adj_4715, n11_adj_4716, n10_adj_4717, 
        n9_adj_4718, n8_adj_4719, n7_adj_4720, n6_adj_4721;
    wire [17:0]d_out_d_11__N_1882;
    
    wire n5_adj_4722, n4_adj_4723, n3_adj_4724, n2_adj_4725, n16246, 
        n16245;
    wire [17:0]d_out_d_11__N_1884;
    
    wire n16099;
    wire [17:0]d_out_d_11__N_1886;
    
    wire n8_adj_4726, n8_adj_4727, n8_adj_4728, n8_adj_4729, n3728, 
        n8_adj_4730, n16090, n16091, n16093, n16094, n16095, n16096;
    wire [17:0]d_out_d_11__N_1888;
    
    wire n16097, n16244, n16243, n16111;
    wire [17:0]d_out_d_11__N_1890;
    
    wire clk_80mhz_enable_1388, n3674;
    wire [17:0]d_out_d_11__N_1892;
    
    wire n916, n917, n918, n919, n920, n921, n922, n923, n924, 
        n925, n926, n927, n928, n929, n930, n931;
    wire [17:0]d_out_d_11__N_2401;
    
    wire clk_80mhz_enable_1387, n16_adj_4731, n14_adj_4732;
    wire [17:0]d_out_d_11__N_2383;
    
    wire n33_adj_4733, n34_adj_4734, n35_adj_4735, n36_adj_4736, n37_adj_4737, 
        n16242, n16241, n16402, n16240, n16239, n16238, n39_adj_4738, 
        n16237, n16236, n16235, n16234, n16015, n16233, n16014, 
        n16401, n16400, n16399, n16398, n16397, n16396, n16395, 
        n8_adj_4739, n16389, n16388, n16387, n16386, n16385, n16384, 
        n16383, n16382, n16381, n17837, n17836, n16232, n16231, 
        n16230, n16229, n16228, n16227, n16226, n16375, n16374, 
        n16373, n16372, n16371, n16013, n16012, n16011, n16225, 
        n16224, n16110, n16223, n16222, n16370, n16010, n16009, 
        n16008, n16007, n16006, n16005, n16004, n16003, n16002, 
        n16001, n16000, n15999, n15998, n15997, n15996, n15995, 
        n15994, n15993, n15992, n16221, n16220, n17812, n16219, 
        n16218, n16217, n17835, n17834, n12613, n1962, n12583, 
        n1960, n12585, n12587, n12589, n12591, n12593, n12595, 
        n1953, n1952, n1951, n1950, n12597, n12599, n1947, n16364, 
        n3897, n16363, n3895, n3893, n16829, clk_80mhz_enable_23, 
        n15991, n16216, n16215, n16362, n50, n16361, n12254, n16360, 
        n12256, n2684, n2682, n2680, n2678, n12258, n16354, n16353, 
        n16352, n2668, n16351, n12260, n2663, n16350, n2659, n2657, 
        n16349, n2655, n16348, n16347, n16345, n16344, n15990, 
        n11962, n2641, n11964, n11966, n11968, n11970, n16343, 
        n11972, n11974, n11976, n12615, n1937, n1935, n1934, n1933, 
        n1932, n1931, n17389, n47, n15989, n16214, n15988, n16213, 
        n17810, n17809, n63_adj_4740, n65, n66_adj_4741, n44, n17832, 
        n41, n12601, n12603, n12605, n12607, n1942, n38, n16212, 
        n15987, n1994, n1993, n12543, n12545, n1989, n12547, n1987, 
        n12549, n12551, n12553, n1983, n12555, n12557, n12559, 
        n1979, n12561, n12563, n12565, n1975, n12567, n1973, n12569, 
        n12571, n1970, n12573, n1968, n12575, n12577, n12579, 
        n1964, n12581, n16342, n3949, n16341, n16340, n3945, n16339, 
        n16338, n16337, n3941, n3938, n3934, n3933, n16331, n16330, 
        n16329, n16328, n3922, n16327, n3920, n3918, n16326, n3916, 
        n16325, n16324, n16323, n3906, n2629, n16318, n11978, 
        n16317, n11980, n2622, n2621, n11982, n11984, n11986, 
        n2617, n11988, n2613, n11990, n2609, n11992, n2607, n2606, 
        n11994, n16316, n11996, n2602, n11998, n12000, n2598, 
        n12002, n12004, n2594, n16315, n12006, n16314, n2586, 
        n2585, n16313, n16312, n16311, n35_adj_4742, n32_adj_4743, 
        n16211, n13_adj_4744, n32_adj_4745, n31_adj_4746, n30_adj_4747, 
        n29_adj_4748, n28_adj_4749, n27_adj_4750, n16210, n16209, 
        n16208, n16207, n16206, n16205, n16204, n16203, n16202, 
        n16310, n16309, n2711, n12246, n16308, n2707, n16307, 
        n12248, n2703, n16306, n2700, n12250, n16305, n2696, n2695, 
        n16304, n16115, n16201, n16200, n12_adj_4751, n16199, n29_adj_4752, 
        n11_adj_4753, n16108, n10_adj_4754, n15985, n9_adj_4755, n15984, 
        n15983, n15982, n15981, n8_adj_4756, n15980, n15979, n15978, 
        n16198, n7_adj_4757, n15977, n16197, n15976, n6_adj_4758, 
        n5_adj_4759, n16196, n4_adj_4760, n15975, n3_adj_4761, n16195, 
        n2_adj_4762, n16107, n16303, n16194, n2_adj_4763, n3_adj_4764, 
        n4_adj_4765, n5_adj_4766, n6_adj_4767, n7_adj_4768, n8_adj_4769, 
        n9_adj_4770, n10_adj_4771, n11_adj_4772, n12_adj_4773, n13_adj_4774, 
        n14_adj_4775, n15_adj_4776, n16_adj_4777, n17_adj_4778, n18_adj_4779, 
        n19_adj_4780, n20_adj_4781, n21_adj_4782, n22_adj_4783, n23_adj_4784, 
        n24_adj_4785, n25_adj_4786, n26_adj_4787, n27_adj_4788, n28_adj_4789, 
        n29_adj_4790, n30_adj_4791, n31_adj_4792, n32_adj_4793, n33_adj_4794, 
        n34_adj_4795, n35_adj_4796, n36_adj_4797, n37_adj_4798, n2_adj_4799, 
        n3_adj_4800, n4_adj_4801, n5_adj_4802, n6_adj_4803, n7_adj_4804, 
        n8_adj_4805, n9_adj_4806, n10_adj_4807, n11_adj_4808, n12_adj_4809, 
        n13_adj_4810, n14_adj_4811, n15_adj_4812, n16_adj_4813, n17_adj_4814, 
        n18_adj_4815, n19_adj_4816, n20_adj_4817, n21_adj_4818, n22_adj_4819, 
        n23_adj_4820, n24_adj_4821, n25_adj_4822, n26_adj_4823, n27_adj_4824, 
        n28_adj_4825, n29_adj_4826, n30_adj_4827, n31_adj_4828, n32_adj_4829, 
        n33_adj_4830, n34_adj_4831, n35_adj_4832, n36_adj_4833, n37_adj_4834, 
        n16193, n15974, cout_adj_4835, cout_adj_4836, n41_adj_4837, 
        n44_adj_4838, n47_adj_4839, n50_adj_4840, n53, n56, n59, 
        n62, n65_adj_4841, n68, n71, n74, n77, n80, n78_adj_4842, 
        n81_adj_4843, n84_adj_4844, n87_adj_4845, n90_adj_4846, n93_adj_4847, 
        n96_adj_4848, n99_adj_4849, n102_adj_4850, n105_adj_4851, n108_adj_4852, 
        n111_adj_4853, n114_adj_4854, n117_adj_4855, n120_adj_4856, 
        n123_adj_4857, n126_adj_4858, n129_adj_4859, n132_adj_4860, 
        n135_adj_4861, n138_adj_4862, n141_adj_4863, n144_adj_4864, 
        n147_adj_4865, n150_adj_4866, n153_adj_4867, n156_adj_4868, 
        n159_adj_4869, n162_adj_4870, n165_adj_4871, n168_adj_4872, 
        n171_adj_4873, n174_adj_4874, n177_adj_4875, n180_adj_4876, 
        n183_adj_4877, n78_adj_4878, n81_adj_4879, n84_adj_4880, n87_adj_4881, 
        n90_adj_4882, n93_adj_4883, n96_adj_4884, n99_adj_4885, n102_adj_4886, 
        n105_adj_4887, n108_adj_4888, n111_adj_4889, n114_adj_4890, 
        n117_adj_4891, n120_adj_4892, n123_adj_4893, n126_adj_4894, 
        n129_adj_4895, n132_adj_4896, n135_adj_4897, n138_adj_4898, 
        n141_adj_4899, n144_adj_4900, n147_adj_4901, n150_adj_4902, 
        n153_adj_4903, n156_adj_4904, n159_adj_4905, n162_adj_4906, 
        n165_adj_4907, n168_adj_4908, n171_adj_4909, n174_adj_4910, 
        n177_adj_4911, n180_adj_4912, n183_adj_4913, n78_adj_4914, n81_adj_4915, 
        n84_adj_4916, n87_adj_4917, n90_adj_4918, n93_adj_4919, n96_adj_4920, 
        n99_adj_4921, n102_adj_4922, n105_adj_4923, n108_adj_4924, n111_adj_4925, 
        n114_adj_4926, n117_adj_4927, n120_adj_4928, n123_adj_4929, 
        n126_adj_4930, n129_adj_4931, n132_adj_4932, n135_adj_4933, 
        n138_adj_4934, n141_adj_4935, n144_adj_4936, n147_adj_4937, 
        n150_adj_4938, n153_adj_4939, n156_adj_4940, n159_adj_4941, 
        n162_adj_4942, n165_adj_4943, n168_adj_4944, n171_adj_4945, 
        n174_adj_4946, n177_adj_4947, n180_adj_4948, n183_adj_4949, 
        n78_adj_4950, n81_adj_4951, n84_adj_4952, n87_adj_4953, n90_adj_4954, 
        n93_adj_4955, n96_adj_4956, n99_adj_4957, n102_adj_4958, n105_adj_4959, 
        n108_adj_4960, n111_adj_4961, n114_adj_4962, n117_adj_4963, 
        n120_adj_4964, n123_adj_4965, n126_adj_4966, n129_adj_4967, 
        n132_adj_4968, n135_adj_4969, n138_adj_4970, n141_adj_4971, 
        n144_adj_4972, n147_adj_4973, n150_adj_4974, n153_adj_4975, 
        n156_adj_4976, n159_adj_4977, n162_adj_4978, n165_adj_4979, 
        n168_adj_4980, n171_adj_4981, n174_adj_4982, n177_adj_4983, 
        n180_adj_4984, n183_adj_4985, n78_adj_4986, n81_adj_4987, n84_adj_4988, 
        n87_adj_4989, n90_adj_4990, n93_adj_4991, n96_adj_4992, n99_adj_4993, 
        n102_adj_4994, n105_adj_4995, n108_adj_4996, n111_adj_4997, 
        n114_adj_4998, n117_adj_4999, n120_adj_5000, n18053, n134, 
        n137, n140, n143, n146, n149, n152, n155, n158, n161, 
        n164, n167, n170, n173, n176, n179, n182, n185, n188, 
        n191, n194, n197, n200, n203, n206, n209, n212, n215, 
        n218, n221, n224, n227, n230, n233, n236, n239, n242, 
        n245, n248, n251, n254, n257, n260, n263, n266, n269, 
        n272, n275, n278, n281, n284, n287, n290, n293, n296, 
        n299, n302, n305, n308, n311, n314, n317, n320, n323, 
        cout_adj_5001, n132_adj_5002, n135_adj_5003, n138_adj_5004, 
        n141_adj_5005, n144_adj_5006, n147_adj_5007, n150_adj_5008, 
        n153_adj_5009, n156_adj_5010, n159_adj_5011, n162_adj_5012, 
        n165_adj_5013, n168_adj_5014, n171_adj_5015, n174_adj_5016, 
        n177_adj_5017, n180_adj_5018, n183_adj_5019, n186, n189, n192, 
        n195, n198, n201, n204, n207, n210, n213_adj_5020, n216, 
        n219, n222, n225, n228, n231, n234, n237, n240, n243, 
        n246, n249, n252, n255, n258, n261, n264, n267, n270, 
        n273, n276, n279, n282, n285, n288, n291, n294, n297, 
        n300, n303, n306, n309, n312, n315, n318, n321, cout_adj_5021, 
        n130, n133, n136, n139, n142, n145, n148, n151, n154, 
        n157, n160, n163, n166, n169, n172, n175, n178, n181, 
        n184, n187, n190, n193, n196, n199, n202, n205, n208, 
        n211, n214, n217, n220, n223, n226, n229, n232, n235, 
        n238, n241, n244, n247, n250, n253, n256, n259, n262, 
        n265, n268, n271, n274, n277, n280, n283, n286, n289, 
        n292, n295, n298, n301, n304, n307, n310, n313, n316, 
        n23_adj_5022, n32_adj_5023, n124, n127, n130_adj_5024, n133_adj_5025, 
        n136_adj_5026, n139_adj_5027, n142_adj_5028, n145_adj_5029, 
        n148_adj_5030, n151_adj_5031, n154_adj_5032, n157_adj_5033, 
        n160_adj_5034, n163_adj_5035, n166_adj_5036, n169_adj_5037, 
        n172_adj_5038, n175_adj_5039, n178_adj_5040, n181_adj_5041, 
        n184_adj_5042, n187_adj_5043, n190_adj_5044, n193_adj_5045, 
        n196_adj_5046, n199_adj_5047, n202_adj_5048, n205_adj_5049, 
        n208_adj_5050, n211_adj_5051, n214_adj_5052, n217_adj_5053, 
        n220_adj_5054, n223_adj_5055, n226_adj_5056, n229_adj_5057, 
        n232_adj_5058, n235_adj_5059, n238_adj_5060, n241_adj_5061, 
        n244_adj_5062, n247_adj_5063, n250_adj_5064, n253_adj_5065, 
        n256_adj_5066, n259_adj_5067, n262_adj_5068, n265_adj_5069, 
        n268_adj_5070, n271_adj_5071, n274_adj_5072, n277_adj_5073, 
        n280_adj_5074, n283_adj_5075, n286_adj_5076, n289_adj_5077, 
        n292_adj_5078, n295_adj_5079, n298_adj_5080, n301_adj_5081, 
        n78_adj_5082, n81_adj_5083, n84_adj_5084, n87_adj_5085, n90_adj_5086, 
        n93_adj_5087, n96_adj_5088, n99_adj_5089, n102_adj_5090, n105_adj_5091, 
        n108_adj_5092, n111_adj_5093, n114_adj_5094, n117_adj_5095, 
        n120_adj_5096, n123_adj_5097, n126_adj_5098, n129_adj_5099, 
        n132_adj_5100, n135_adj_5101, n138_adj_5102, n141_adj_5103, 
        n144_adj_5104, n147_adj_5105, n150_adj_5106, n153_adj_5107, 
        n156_adj_5108, n159_adj_5109, n162_adj_5110, n165_adj_5111, 
        n168_adj_5112, n171_adj_5113, n174_adj_5114, n177_adj_5115, 
        n180_adj_5116, n183_adj_5117, n78_adj_5118, n81_adj_5119, n84_adj_5120, 
        n87_adj_5121, n90_adj_5122, n93_adj_5123, n96_adj_5124, n99_adj_5125, 
        n102_adj_5126, n105_adj_5127, n108_adj_5128, n111_adj_5129, 
        n114_adj_5130, n117_adj_5131, n120_adj_5132, n123_adj_5133, 
        n126_adj_5134, n129_adj_5135, n132_adj_5136, n135_adj_5137, 
        n138_adj_5138, n141_adj_5139, n144_adj_5140, n147_adj_5141, 
        n150_adj_5142, n153_adj_5143, n156_adj_5144, n159_adj_5145, 
        n162_adj_5146, n165_adj_5147, n168_adj_5148, n171_adj_5149, 
        n174_adj_5150, n177_adj_5151, n180_adj_5152, n183_adj_5153, 
        n76, n79, n82, n85, n88, n91, n94, n97, n100, n103, 
        n106, n109, n112, n115, n118, n78_adj_5154, n81_adj_5155, 
        n84_adj_5156, n87_adj_5157, n90_adj_5158, n93_adj_5159, n96_adj_5160, 
        n99_adj_5161, n102_adj_5162, n105_adj_5163, n108_adj_5164, n111_adj_5165, 
        n114_adj_5166, n117_adj_5167, n120_adj_5168, n123_adj_5169, 
        n126_adj_5170, n129_adj_5171, n132_adj_5172, n135_adj_5173, 
        n138_adj_5174, n141_adj_5175, n144_adj_5176, n147_adj_5177, 
        n150_adj_5178, n153_adj_5179, n156_adj_5180, n159_adj_5181, 
        n162_adj_5182, n165_adj_5183, n168_adj_5184, n171_adj_5185, 
        n174_adj_5186, n177_adj_5187, n180_adj_5188, n183_adj_5189, 
        n45_adj_5190, n48_adj_5191, n51_adj_5192, n54_adj_5193, n57_adj_5194, 
        n60_adj_5195, n63_adj_5196, n66_adj_5197, n69_adj_5198, n72_adj_5199, 
        n75_adj_5200, n78_adj_5201, n81_adj_5202, n84_adj_5203, n87_adj_5204, 
        n90_adj_5205, cout_adj_5206, cout_adj_5207, n36_adj_5208, n39_adj_5209, 
        n42_adj_5210, n45_adj_5211, n48_adj_5212, n51_adj_5213, n54_adj_5214, 
        n57_adj_5215, n60_adj_5216, n63_adj_5217, n66_adj_5218, n69_adj_5219, 
        n72_adj_5220, n75_adj_5221, n78_adj_5222, n81_adj_5223, n54_adj_5224, 
        n57_adj_5225, n60_adj_5226, n63_adj_5227, n66_adj_5228, n69_adj_5229, 
        n72_adj_5230, n75_adj_5231, n78_adj_5232, n81_adj_5233, n84_adj_5234, 
        n87_adj_5235, n90_adj_5236, n93_adj_5237, n96_adj_5238, n99_adj_5239, 
        n102_adj_5240, n105_adj_5241, n108_adj_5242, n111_adj_5243, 
        n114_adj_5244, n117_adj_5245, n120_adj_5246, n123_adj_5247, 
        n126_adj_5248, n78_adj_5249, n81_adj_5250, n84_adj_5251, n87_adj_5252, 
        n90_adj_5253, n93_adj_5254, n96_adj_5255, n99_adj_5256, n102_adj_5257, 
        n105_adj_5258, n108_adj_5259, n111_adj_5260, n114_adj_5261, 
        n117_adj_5262, n120_adj_5263, n123_adj_5264, n126_adj_5265, 
        n129_adj_5266, n132_adj_5267, n135_adj_5268, n138_adj_5269, 
        n141_adj_5270, n144_adj_5271, n147_adj_5272, n150_adj_5273, 
        n153_adj_5274, n156_adj_5275, n159_adj_5276, n162_adj_5277, 
        n165_adj_5278, n168_adj_5279, n171_adj_5280, n174_adj_5281, 
        n177_adj_5282, n180_adj_5283, n183_adj_5284, n78_adj_5285, n81_adj_5286, 
        n84_adj_5287, n87_adj_5288, n90_adj_5289, n93_adj_5290, n96_adj_5291, 
        n99_adj_5292, n102_adj_5293, n105_adj_5294, n108_adj_5295, n111_adj_5296, 
        n114_adj_5297, n117_adj_5298, n120_adj_5299, n123_adj_5300, 
        n126_adj_5301, n129_adj_5302, n132_adj_5303, n135_adj_5304, 
        n138_adj_5305, n141_adj_5306, n144_adj_5307, n147_adj_5308, 
        n150_adj_5309, n153_adj_5310, n156_adj_5311, n159_adj_5312, 
        n162_adj_5313, n165_adj_5314, n168_adj_5315, n171_adj_5316, 
        n174_adj_5317, n177_adj_5318, n180_adj_5319, n183_adj_5320, 
        n78_adj_5321, n81_adj_5322, n84_adj_5323, n87_adj_5324, n90_adj_5325, 
        n93_adj_5326, n96_adj_5327, n99_adj_5328, n102_adj_5329, n105_adj_5330, 
        n108_adj_5331, n111_adj_5332, n114_adj_5333, n117_adj_5334, 
        n120_adj_5335, n123_adj_5336, n126_adj_5337, n129_adj_5338, 
        n132_adj_5339, n135_adj_5340, n138_adj_5341, n141_adj_5342, 
        n144_adj_5343, n147_adj_5344, n150_adj_5345, n153_adj_5346, 
        n156_adj_5347, n159_adj_5348, n162_adj_5349, n165_adj_5350, 
        n168_adj_5351, n171_adj_5352, n174_adj_5353, n177_adj_5354, 
        n180_adj_5355, n183_adj_5356, n78_adj_5357, n81_adj_5358, n84_adj_5359, 
        n87_adj_5360, n90_adj_5361, n93_adj_5362, n96_adj_5363, n99_adj_5364, 
        n102_adj_5365, n105_adj_5366, n108_adj_5367, n111_adj_5368, 
        n114_adj_5369, n117_adj_5370, n120_adj_5371, n123_adj_5372, 
        n126_adj_5373, n129_adj_5374, n132_adj_5375, n135_adj_5376, 
        n138_adj_5377, n141_adj_5378, n144_adj_5379, n147_adj_5380, 
        n150_adj_5381, n153_adj_5382, n156_adj_5383, n159_adj_5384, 
        n162_adj_5385, n165_adj_5386, n168_adj_5387, n171_adj_5388, 
        n174_adj_5389, n177_adj_5390, n180_adj_5391, n183_adj_5392, 
        n45_adj_5393, n48_adj_5394, n51_adj_5395, n54_adj_5396, n57_adj_5397, 
        n60_adj_5398, n63_adj_5399, n66_adj_5400, n69_adj_5401, n72_adj_5402, 
        n75_adj_5403, n78_adj_5404, n81_adj_5405, n84_adj_5406, n87_adj_5407, 
        n90_adj_5408, n78_adj_5409, n81_adj_5410, n84_adj_5411, n87_adj_5412, 
        n90_adj_5413, n93_adj_5414, n96_adj_5415, n99_adj_5416, n102_adj_5417, 
        n105_adj_5418, n108_adj_5419, n111_adj_5420, n114_adj_5421, 
        n117_adj_5422, n120_adj_5423, n123_adj_5424, n126_adj_5425, 
        n129_adj_5426, n132_adj_5427, n135_adj_5428, n138_adj_5429, 
        n141_adj_5430, n144_adj_5431, n147_adj_5432, n150_adj_5433, 
        n153_adj_5434, n156_adj_5435, n159_adj_5436, n162_adj_5437, 
        n165_adj_5438, n168_adj_5439, n171_adj_5440, n174_adj_5441, 
        n177_adj_5442, n180_adj_5443, n183_adj_5444, n45_adj_5445, n48_adj_5446, 
        n51_adj_5447, n54_adj_5448, n57_adj_5449, n60_adj_5450, n63_adj_5451, 
        n66_adj_5452, n69_adj_5453, n72_adj_5454, n75_adj_5455, n78_adj_5456, 
        n81_adj_5457, n84_adj_5458, n87_adj_5459, n90_adj_5460, cout_adj_5461, 
        n15973, n15972, n15971, n15970, n15969, n15968, n15963, 
        n15962, n15961, n15960, n15959, n15958, n15957, n15956, 
        n15955, n15954, n15953, n15952, n15951, n15950, n15949, 
        n15948, n15947, n15946, n15941, n15940, n15939, n15938, 
        n15937, n15936, cout_adj_5462, cout_adj_5463, cout_adj_5464, 
        n12261, n12259, n12257, n12255, n12253, n12251, n12249, 
        n12247, n12245, n16109, n16106, n15022, n12542, n16259, 
        n16254, n16252, n16258, n16253, n16191, n16190, n78_adj_5465, 
        n81_adj_5466, n16092, n84_adj_5467, n87_adj_5468, n16189, 
        n90_adj_5469, n93_adj_5470, n16188, n96_adj_5471, n99_adj_5472, 
        n102_adj_5473, n105_adj_5474, n108_adj_5475, n16105, n111_adj_5476, 
        n114_adj_5477, n16187, n117_adj_5478, n120_adj_5479, n16186, 
        n123_adj_5480, n126_adj_5481, n15021, n129_adj_5482, n132_adj_5483, 
        n16257, n135_adj_5484, n138_adj_5485, n141_adj_5486, n16185, 
        n144_adj_5487, n147_adj_5488, n16184, n150_adj_5489, n153_adj_5490, 
        n156_adj_5491, n159_adj_5492, n16183, n162_adj_5493, n165_adj_5494, 
        n16182, n168_adj_5495, n171_adj_5496, n174_adj_5497, n177_adj_5498, 
        n16181, n180_adj_5499, n183_adj_5500, n16180, n16256, n12538, 
        n16179, n16178, n16104, n15020, n15935, n15934, n15933, 
        n15932, n15931, n15930, n15929, n15928, n15927, n15926, 
        n15925, n15924, n15920, n15919, n15019, n15018, cout_adj_5501, 
        n15017, n16177, n16176, n16175, n12701, n16174, n16170, 
        n16169, n16168, n16167, n16166, n16302, n78_adj_5502, n81_adj_5503, 
        n84_adj_5504, n87_adj_5505, n90_adj_5506, n93_adj_5507, n16165, 
        n96_adj_5508, n16164, n99_adj_5509, n16163, n102_adj_5510, 
        n16162, n105_adj_5511, n16161, n108_adj_5512, n16160, n111_adj_5513, 
        n16159, n114_adj_5514, n16158, n117_adj_5515, n16157, n120_adj_5516, 
        n16156, n123_adj_5517, n16155, n126_adj_5518, n16154, n129_adj_5519, 
        n16153, n132_adj_5520, n135_adj_5521, n138_adj_5522, n141_adj_5523, 
        n16151, n144_adj_5524, n147_adj_5525, n150_adj_5526, n153_adj_5527, 
        n156_adj_5528, n159_adj_5529, n162_adj_5530, n165_adj_5531, 
        n168_adj_5532, n171_adj_5533, n174_adj_5534, n177_adj_5535, 
        n180_adj_5536, n183_adj_5537, n16150, n16149, n16148, n16147, 
        n16146, n16145, n16144, n16143, n16142, n16141, n16140, 
        n16139, n16138, n16137, n16301, n16136, n16135, n16134, 
        n16098, n16130, n16129, n16128, n16127, n16126, n16125, 
        n16124, n16123, n16122, n16121, n16120, n16119, n16300, 
        n16299, n16118, n16117, n16298, n16297, n16116, n16103, 
        n16867, n16102, n16296, n16295, n15918, n16294, n16293, 
        n16101, n16100, n16292, n16291, n16290, n16289, n16288, 
        n16287, n16286, n17288, n16285, n16284, n16283, n16282, 
        n16281, n16280, n15016, n16279, n16278, n16277, n16276, 
        n78_adj_5538, n81_adj_5539, n16275, n84_adj_5540, n16274, 
        n87_adj_5541, n16273, n90_adj_5542, n93_adj_5543, n96_adj_5544, 
        n99_adj_5545, n102_adj_5546, n105_adj_5547, n16272, n108_adj_5548, 
        n111_adj_5549, n114_adj_5550, n117_adj_5551, n120_adj_5552, 
        n123_adj_5553, n126_adj_5554, n15917, n129_adj_5555, n132_adj_5556, 
        n135_adj_5557, n16492, n138_adj_5558, n141_adj_5559, n16491, 
        n144_adj_5560, n16490, n147_adj_5561, n150_adj_5562, n16489, 
        n153_adj_5563, n16271, n156_adj_5564, n16488, n159_adj_5565, 
        n16487, n162_adj_5566, n16270, n165_adj_5567, n16269, n168_adj_5568, 
        n16255, n171_adj_5569, n16486, n174_adj_5570, n177_adj_5571, 
        n180_adj_5572, n183_adj_5573, n16485, n16484, n12540, n16478, 
        n8_adj_5574, n16477, n16476, n12710, n11959, n16268, n11963, 
        n11965, n16267, n11969, n11971, n16266, n11975, n11977, 
        n16265, n16264, n11983, n16263, n11987, n11989, n11991, 
        n16262, n11995, n11997, n11999, n16475, n16261, n12003, 
        n16260, n12007, n16474, n16473, n16472, n15015, n16466, 
        n16465, n16464, n16463, n16462, clk_80mhz_enable_1408, n16461, 
        n16460, n16459, n16458, n15014, n12424, n16452, n16451, 
        n16450, n16449, n16448, n16447, n16446, n16445, n16444, 
        n15916, n15915, n15914, n15913, n15912, n15911, n15910, 
        n15909, n15908, n15907, n15906, n15905, n15904, n15903, 
        n15902, n15901, n15900, n15899, n15898, n15897, n15896, 
        n15895, n15894, n15893, n15892, n15891, n15890, n15889, 
        n15888, n15887, n15886, n15885, n15884, n15883, n15882, 
        n15881, n15880, n15879, n15878, n15877, n15876, n15875, 
        n15874, n15873, n15872, n15871, n15870, n15869, n15868, 
        n15867, n15866, n15865, n15864, n15863, n15862, n15861, 
        n15860, n15859, n15858, n15857, n15856, n15855, n15854, 
        n15853, n15852, n15851, n15850, n15849, n15848, n15847, 
        n15846, n15845, n15844, n15843, n15842, n15841, n15840, 
        n15839, n15838, n15837, n15836, n15835, n15834, n15833, 
        n15832, n15831, n15830, n15829, n15828, n15827, n15826, 
        n15825, n15824, n15823, n15822, n15812, n15811, n15810, 
        n15809, n15808, n15807, n15806, n15805, n15804, n15803, 
        n15802, cout_adj_5575, n15801, n15800, n15799, n15798, n15797, 
        n15796, n15795, n15791, n15790, n15789, n15788, n15787, 
        n15786, n15785, n15784, n15783, n15782, n15781, n15780, 
        n15779, n15778, n15777, n15776, n15775, n15774, n15772, 
        n15771, n15770, n15769, n15768, n15767, n15766, n15765, 
        n15764, n15763, n15762, n15761, n15760, n15759, n15758, 
        n15757, n15756, n15755, n15754, n15753, n15752, n15751, 
        n15750, n15749, n15748, n15747, n15744, n15743, n15742, 
        n15741, n15740, n15739, n15738, n15737, n15736, n15735, 
        n15734, n15733, n15732, n15731, cout_adj_5576, n15730, n15729, 
        n15728, n15727, n15723, n15722, n15721, n15720, n15719, 
        n15718, n15717, n15716, n15714, n15713, n15712, n15711, 
        n15710, n15709, n15708, n15707, n15706, n15705, n15704, 
        n15703, n15702, n15701, n15700, n15699, n15698, n15697, 
        n15693, n15692, n15691, n15690, n15689, n15688, n15687, 
        n15686, n15685, n15684, n15683, n15682, n76_adj_5577, n79_adj_5578, 
        n15679, n82_adj_5579, n15678, n85_adj_5580, n15677, n88_adj_5581, 
        n15676, n91_adj_5582, n15675, n94_adj_5583, n15674, n97_adj_5584, 
        n15673, n100_adj_5585, n15672, n103_adj_5586, n15671, n106_adj_5587, 
        n15670, n109_adj_5588, n15669, n112_adj_5589, n15668, n115_adj_5590, 
        n15667, n118_adj_5591, n15666, n15665, n15664, n15663, n15662, 
        n15658, n15657, n15656, n15655, n15654, n15653, n15652, 
        n15651, n15650, n15649, n15648, n15647, n15646, n15645, 
        n15644, n15643, n15642, n15641, n15640, n15639, n15638, 
        n15637, n15636, n15635, n15634, n15633, n15632, n15631, 
        n15630, n15629, n15628, n15627, n15626, n15625, n15624, 
        n15623, n15622, n15621, n15620, n15619, n15618, n15617, 
        n15616, n15615, n15614, n15613, n15612, n15611, n15610, 
        n15609, n15608, n15607, n15606, n15605, n15604, n15603, 
        n15602, n15601, n15600, n15599, n15598, n15597, n15596, 
        n15595, n15594, n15593, n15592, n15591, n15590, n15589, 
        n15588, n15587, n15585, n15584, n15583, n15582, n15581, 
        n15580, n15579, n15578, n15577, n15576, n15575, n15574, 
        n15573, n15572, n15571, n15570, n15569, n15568, n15566, 
        n15565, n15564, n15563, n15562, n15561, n15560, n15559, 
        n15558, n15557, n15556, n15555, n15554, n45_adj_5592, n15553, 
        n48_adj_5593, n15552, n51_adj_5594, n15551, n54_adj_5595, 
        n15550, n57_adj_5596, n15549, n60_adj_5597, n15547, n63_adj_5598, 
        n15546, n66_adj_5599, n15545, n69_adj_5600, n15544, n72_adj_5601, 
        n15543, n75_adj_5602, n15542, n78_adj_5603, n15541, n81_adj_5604, 
        n15540, n84_adj_5605, n15539, n87_adj_5606, n15538, n90_adj_5607, 
        n15537, n15536, n15535, n15534, n15533, n15532, n15531, 
        n15530, n15528, n15527, n15526, n15525, n15524, n15523, 
        n15521, n15520, n15519, n15518, n15517, n15516, n15515, 
        n15514, n15513, n15512, n15511, n15510, n15509, n15508, 
        n15507, n15506, n15505, n15504, n15499, n15498, n15497, 
        n15496, n15495, n15494, n15493, n15492, n15491, n15490, 
        n15489, n15488, n15487, n15486, n15485, n15484, n15483, 
        n15482, n15478, n15477, n15476, n15475, n15474, n15473, 
        n15472, n15471, n15470, n15469, n15468, n15467, n15466, 
        n15465, n15464, n15463, n15462, n15461, n15460, n15459, 
        n15458, n15457, n15456, n15455, n15454, n15453, n15452, 
        n15451, n15450, n15449, n15448, n15447, n15446, n15445, 
        n15444, n15443, n15442, n15441, n15440, n15439, n15438, 
        n15437, n15436, n15435, n15434, n15433, n15432, n15431, 
        n15430, n15429, n15428, n15427, n15426, n15425, n15424, 
        n15423, n15422, n15421, n15420, n15419, n15417, n15416, 
        n15415, n15414, n15413, n15412, n15411, n15410, n15409, 
        n15408, n15407, n15406, n15405, n15404, n15403, n15402, 
        n15401, n15400, n15393, n15392, n15391, n15390, n15389, 
        n15388, n15387, n15386, n15385, n15384, n15383, n15382, 
        n15381, n15380, n15379, n15378, n15377, n15376, n15372, 
        n15371, n15370, n15369, n15368, n15367, n15366, n15365, 
        n15364, n15363, n15362, n15361, n15360, n15359, n15358, 
        n15357, n15356, n15355, n15353, n15352, n15351, n15350, 
        n15349, n15348, n15347, n15346, n15345, n15344, n15343, 
        n15342, n15341, n15340, n15339, n15338, n15337, n15336, 
        n15331, n15330, n15329, n15328, n15327, n15326, n15325, 
        n15324, n15323, n15322, n15321, n15320, n15319, n15318, 
        n15317, n15316, n15315, n15314, n15310, n15309, n15308, 
        n15307, n15306, n15305, n15304, n15303, n15302, n15301, 
        n15300, n15299, n15298, n15297, n15296, n15295, n15294, 
        n15293, n15291, n15290, n15289, n15288, n15287, n15286, 
        n15285, n15284, n15283, n15282, n15281, n15280, n15279, 
        n15278, n15277, n15276, n15275, n15274, n15269, n15268, 
        n15267, n15266, n15265, n15264, n15263, n15262, n15261, 
        n15260, n15259, n15258, n15257, n15256, n15255, n15254, 
        n15253, n15252, n15251, n15250, n15249, n78_adj_5608, n15248, 
        n81_adj_5609, n15247, n84_adj_5610, n15246, n87_adj_5611, 
        n15245, n90_adj_5612, n15244, n93_adj_5613, n15243, n96_adj_5614, 
        n15242, n99_adj_5615, n15241, n102_adj_5616, n15240, n105_adj_5617, 
        n15239, n108_adj_5618, n15237, n111_adj_5619, n15236, n114_adj_5620, 
        n15235, n117_adj_5621, n15234, n120_adj_5622, n15233, n123_adj_5623, 
        n15232, n126_adj_5624, n15231, n129_adj_5625, n15230, n132_adj_5626, 
        n15229, n135_adj_5627, n15228, n138_adj_5628, n15227, n141_adj_5629, 
        n15226, n144_adj_5630, n15225, n147_adj_5631, n15224, n150_adj_5632, 
        n15223, n153_adj_5633, n15222, n156_adj_5634, n15221, n159_adj_5635, 
        n15220, n162_adj_5636, n165_adj_5637, n15217, n168_adj_5638, 
        n15216, n171_adj_5639, n15215, n174_adj_5640, n15214, n177_adj_5641, 
        n15213, n180_adj_5642, n15212, n183_adj_5643, n15211, n15210, 
        n15209, n15208, n15207, n15206, n15205, n15204, n15203, 
        n15202, n15201, n15200, n15199, n15198, n15197, n15196, 
        n15195, n15194, n15193, n15192, n15191, n15190, n15189, 
        n15188, n15187, n15186, n15185, n15184, n15183, n15182, 
        n15181, n15180, n15179, n15178, n15177, n15176, n15175, 
        n15174, n15173, n15172, n15171, n15170, n15169, n15168, 
        n15167, n15166, n15165, n15164, n15163, n15162, n15161, 
        n15160, n15159, n15158, n15157, n15156, n15155, n15154, 
        n15153, n15152, n15151, n15150, n15149, n15148, n15147, 
        n15146, n15145, n15144, n15143, n15142, n15141, n15140, 
        n15139, n15138, n15137, n15136, n15135, n15134, n15133, 
        n15132, n15131, n15130, n15129, n15128, n15127, n15126, 
        n15125, n15124, n15123, n15122, n15121, n15120, n15119, 
        n15118, n15117, n15116, n15115, n15114, n15113, n15112, 
        n15111, n15110, n15109, n15108, n15107, n15106, n15105, 
        n15104, n15103, n15101, n15100, n15099, n15098, n15097, 
        cout_adj_5644, n15096, n15095, n15094, n15093, n15092, n15091, 
        n15090, n15089, n15088, n15087, n15086, n15085, n15084, 
        n15083, n15082, n15081, n15080, n15079, n15078, n15077, 
        n15076, n15075, n15074, n15073, n15072, n15071, n15070, 
        n15069, n15068, n15067, n15066, n15064, n15063, n15062, 
        n15061, n15060, n15059, n15058, n15057, n15056, n15055, 
        n15054, n15053, n15052, n15051, n15050, n15049, n15048, 
        n15047, n15046, n15045, n15044, n15043, n15042, n15041, 
        n15040, n15039, n15038, n15037, n15036, n15035, n15034, 
        n15033, n15032, n15031, n15030, n15029, n15028, n15027, 
        n15026, n15025, n15024, n15023, n78_adj_5645, n81_adj_5646, 
        n84_adj_5647, n87_adj_5648, n90_adj_5649, n93_adj_5650, n96_adj_5651, 
        n99_adj_5652, n102_adj_5653, n105_adj_5654, n108_adj_5655, n111_adj_5656, 
        n114_adj_5657, n117_adj_5658, n120_adj_5659, n123_adj_5660, 
        n126_adj_5661, n129_adj_5662, n132_adj_5663, n135_adj_5664, 
        n138_adj_5665, n141_adj_5666, n144_adj_5667, n147_adj_5668, 
        n150_adj_5669, n153_adj_5670, n156_adj_5671, n159_adj_5672, 
        n162_adj_5673, n165_adj_5674, n168_adj_5675, n171_adj_5676, 
        n174_adj_5677, n177_adj_5678, n180_adj_5679, n183_adj_5680, 
        n17778, n37_adj_5681, n40, n43, n46, n49, n17325, n52, 
        n55, n58, n61, n64, n67, n70, n15013, n15012, n15011, 
        n15010, n15009, n15008, n15007, n15006, n15005, n15003, 
        n14998, n14997, n14967, n15000, n15001, n14993, n14996, 
        n45_adj_5682, n14995, n48_adj_5683, n14994, n51_adj_5684, 
        n54_adj_5685, n57_adj_5686, n15004, n60_adj_5687, n63_adj_5688, 
        n66_adj_5689, n69_adj_5690, n72_adj_5691, n75_adj_5692, n78_adj_5693, 
        n17828, n81_adj_5694, n84_adj_5695, n17827, n87_adj_5696, 
        n90_adj_5697, n17826, n17825, n16869, n8_adj_5698, n17823, 
        n17822, n16837, n17081, n17820, n17075, n17073, n17817, 
        n17022, n17815, n8_adj_5699, clk_80mhz_enable_1411, n18096, 
        n17069, n16944, n17032, cout_adj_5700, n16842, n17302, n15002, 
        n17814, n17813, n14999;
    
    VHI i2 (.Z(VCC_net));
    \uart_rx(CLKS_PER_BIT=87)  uart_rx_inst (.clk_80mhz(clk_80mhz), .i_Rx_Serial_c(i_Rx_Serial_c), 
            .o_Rx_Byte1({o_Rx_Byte1}), .o_Rx_DV1(o_Rx_DV1), .GND_net(GND_net), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(179[33] 184[5])
    CCU2C _add_1_1490_add_4_8 (.A0(d_d7[5]), .B0(d7[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[6]), .B1(d7[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16115), .COUT(n16116), .S0(d8_71__N_1603[5]), .S1(d8_71__N_1603[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_19 (.A0(d6_adj_5715[52]), .B0(cout_adj_5464), 
          .C0(n135_adj_4897), .D0(n21_adj_4577), .A1(d6_adj_5715[53]), 
          .B1(cout_adj_5464), .C1(n132_adj_4896), .D1(n20_adj_4578), .CIN(n16182), 
          .COUT(n16183), .S0(d7_71__N_1531_adj_5743[52]), .S1(d7_71__N_1531_adj_5743[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_6 (.A0(d_d7[3]), .B0(d7[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[4]), .B1(d7[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16114), .COUT(n16115), .S0(d8_71__N_1603[3]), .S1(d8_71__N_1603[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_34 (.A0(d2_adj_5711[67]), .B0(d1_adj_5710[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[68]), .B1(d1_adj_5710[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16038), .COUT(n16039), .S0(n90_adj_5612), 
          .S1(n87_adj_5611));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_34.INJECT1_1 = "NO";
    OB led_pad_6 (.I(led_c_6), .O(led[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(44[22:25])
    CCU2C _add_1_1418_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5464), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16174));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1418_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1418_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_1.INJECT1_1 = "NO";
    FD1S3AX o_Rx_DV_40 (.D(o_Rx_DV1), .CK(clk_80mhz), .Q(o_Rx_DV));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam o_Rx_DV_40.GSR = "ENABLED";
    CCU2C _add_1_1490_add_4_4 (.A0(d_d7[1]), .B0(d7[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[2]), .B1(d7[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16113), .COUT(n16114), .S0(d8_71__N_1603[1]), .S1(d8_71__N_1603[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_4.INJECT1_1 = "NO";
    Mixer Mixer_inst (.MixerOutSin({MixerOutSin}), .clk_80mhz(clk_80mhz), 
          .DiffOut_c(DiffOut_c), .MixerOutCos({MixerOutCos}), .RFIn_c(RFIn_c), 
          .\LOSine[1] (LOSine[1]), .MixerOutSin_11__N_236({MixerOutSin_11__N_236}), 
          .\LOCosine[1] (LOCosine[1]), .MixerOutCos_11__N_250({MixerOutCos_11__N_250}), 
          .\LOSine[6] (LOSine[6]), .\LOSine[11] (LOSine[11]), .\LOSine[10] (LOSine[10]), 
          .\LOSine[9] (LOSine[9]), .\LOSine[5] (LOSine[5]), .\LOSine[4] (LOSine[4]), 
          .\LOSine[8] (LOSine[8]), .\LOSine[7] (LOSine[7]), .\LOSine[3] (LOSine[3]), 
          .\LOSine[2] (LOSine[2]), .\LOCosine[12] (LOCosine[12]), .\LOCosine[11] (LOCosine[11]), 
          .\LOCosine[10] (LOCosine[10]), .\LOCosine[9] (LOCosine[9]), .\LOCosine[8] (LOCosine[8]), 
          .\LOCosine[7] (LOCosine[7]), .\LOCosine[6] (LOCosine[6]), .\LOCosine[5] (LOCosine[5]), 
          .\LOCosine[4] (LOCosine[4]), .\LOCosine[3] (LOCosine[3]), .\LOCosine[2] (LOCosine[2]), 
          .\LOSine[12] (LOSine[12])) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(122[10] 130[5])
    CCU2C _add_1_1544_add_4_32 (.A0(d2_adj_5711[65]), .B0(d1_adj_5710[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[66]), .B1(d1_adj_5710[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16037), .COUT(n16038), .S0(n96_adj_5614), 
          .S1(n93_adj_5613));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_32.INJECT1_1 = "NO";
    CCU2C add_3659_5 (.A0(n50), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(n17826), .C1(n47), .D1(VCC_net), 
          .CIN(n16371), .COUT(n16372), .S0(n57), .S1(n54));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3659_5.INIT0 = 16'haaa0;
    defparam add_3659_5.INIT1 = 16'h6969;
    defparam add_3659_5.INJECT1_0 = "NO";
    defparam add_3659_5.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_36 (.A0(d_d_tmp[33]), .B0(d_tmp[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[34]), .B1(d_tmp[34]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15621), .COUT(n15622), .S0(d6_71__N_1459[33]), 
          .S1(d6_71__N_1459[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_12 (.A0(d5_adj_5714[45]), .B0(d4_adj_5713[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[46]), .B1(d4_adj_5713[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16157), .COUT(n16158), .S0(n156_adj_5564), 
          .S1(n153_adj_5563));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_8 (.A0(d5_adj_5714[41]), .B0(d4_adj_5713[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[42]), .B1(d4_adj_5713[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16155), .COUT(n16156), .S0(n168_adj_5568), 
          .S1(n165_adj_5567));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_23 (.A0(d4[56]), .B0(cout_adj_2810), .C0(n123_adj_5300), 
          .D0(d5[56]), .A1(d4[57]), .B1(cout_adj_2810), .C1(n120_adj_5299), 
          .D1(d5[57]), .CIN(n16054), .COUT(n16055), .S0(d5_71__N_706[56]), 
          .S1(d5_71__N_706[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_17 (.A0(d6_adj_5715[50]), .B0(cout_adj_5464), 
          .C0(n141_adj_4899), .D0(n23_adj_4557), .A1(d6_adj_5715[51]), 
          .B1(cout_adj_5464), .C1(n138_adj_4898), .D1(n22_adj_4576), .CIN(n16181), 
          .COUT(n16182), .S0(d7_71__N_1531_adj_5743[50]), .S1(d7_71__N_1531_adj_5743[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[0]), .B1(d7[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16113), .S1(d8_71__N_1603[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1490_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_12 (.A0(counter[9]), .B0(DataInReg[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16112), .S1(cout_adj_5576));
    defparam _add_1_1565_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1565_add_4_12.INIT1 = 16'h0000;
    defparam _add_1_1565_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_12.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i0 (.D(phase_inc_carrGen[0]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i0.GSR = "ENABLED";
    CCU2C _add_1_1565_add_4_10 (.A0(counter[7]), .B0(DataInReg[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[8]), .B1(DataInReg[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16111), .COUT(n16112));
    defparam _add_1_1565_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1565_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1565_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_8 (.A0(counter[5]), .B0(DataInReg[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[6]), .B1(DataInReg[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16110), .COUT(n16111));
    defparam _add_1_1565_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1565_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1565_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_8.INJECT1_1 = "NO";
    PWM PWM_inst (.\DataInReg[0] (DataInReg[0]), .clk_80mhz(clk_80mhz), 
        .\DataInReg_11__N_1856[0] (DataInReg_11__N_1856[0]), .counter({counter}), 
        .GND_net(GND_net), .VCC_net(VCC_net), .\DataInReg[1] (DataInReg[1]), 
        .\DataInReg_11__N_1856[1] (DataInReg_11__N_1856[1]), .\DataInReg[2] (DataInReg[2]), 
        .\DataInReg_11__N_1856[2] (DataInReg_11__N_1856[2]), .\DataInReg[3] (DataInReg[3]), 
        .\DataInReg_11__N_1856[3] (DataInReg_11__N_1856[3]), .\DataInReg[4] (DataInReg[4]), 
        .\DataInReg_11__N_1856[4] (DataInReg_11__N_1856[4]), .\DataInReg[5] (DataInReg[5]), 
        .\DataInReg_11__N_1856[5] (DataInReg_11__N_1856[5]), .\DataInReg[6] (DataInReg[6]), 
        .\DataInReg_11__N_1856[6] (DataInReg_11__N_1856[6]), .\DataInReg[7] (DataInReg[7]), 
        .\DataInReg_11__N_1856[7] (DataInReg_11__N_1856[7]), .\DataInReg[8] (DataInReg[8]), 
        .\DataInReg_11__N_1856[8] (DataInReg_11__N_1856[8]), .\DataInReg[9] (DataInReg[9]), 
        .\DemodOut[9] (DemodOut[9])) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(156[8] 160[5])
    CCU2C _add_1_1565_add_4_6 (.A0(counter[3]), .B0(DataInReg[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[4]), .B1(DataInReg[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16109), .COUT(n16110));
    defparam _add_1_1565_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1565_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1565_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_30 (.A0(d2_adj_5711[63]), .B0(d1_adj_5710[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[64]), .B1(d1_adj_5710[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16036), .COUT(n16037), .S0(n102_adj_5616), 
          .S1(n99_adj_5615));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_4 (.A0(counter[1]), .B0(DataInReg[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[2]), .B1(DataInReg[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16108), .COUT(n16109));
    defparam _add_1_1565_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1565_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1565_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1565_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[0]), .B1(DataInReg[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16108));
    defparam _add_1_1565_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1565_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1565_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1565_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_28 (.A0(d2_adj_5711[61]), .B0(d1_adj_5710[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[62]), .B1(d1_adj_5710[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16035), .COUT(n16036), .S0(n108_adj_5618), 
          .S1(n105_adj_5617));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_37 (.A0(d_d9_adj_5722[71]), .B0(d9_adj_5721[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16107), .S0(n76_adj_5577));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_37.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_37.INIT1 = 16'h0000;
    defparam _add_1_1409_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_10 (.A0(d2_adj_5711[43]), .B0(d1_adj_5710[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[44]), .B1(d1_adj_5710[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16026), .COUT(n16027), .S0(n162_adj_5636), 
          .S1(n159_adj_5635));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_35 (.A0(d_d9_adj_5722[69]), .B0(d9_adj_5721[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[70]), .B1(d9_adj_5721[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16106), .COUT(n16107), .S0(n82_adj_5579), 
          .S1(n79_adj_5578));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_35.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_35.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_33 (.A0(d_d9_adj_5722[67]), .B0(d9_adj_5721[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[68]), .B1(d9_adj_5721[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16105), .COUT(n16106), .S0(n88_adj_5581), 
          .S1(n85_adj_5580));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_33.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_33.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_31 (.A0(d_d9_adj_5722[65]), .B0(d9_adj_5721[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[66]), .B1(d9_adj_5721[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16104), .COUT(n16105), .S0(n94_adj_5583), 
          .S1(n91_adj_5582));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_31.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_31.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_29 (.A0(d_d9_adj_5722[63]), .B0(d9_adj_5721[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[64]), .B1(d9_adj_5721[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16103), .COUT(n16104), .S0(n100_adj_5585), 
          .S1(n97_adj_5584));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_29.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_29.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_8 (.A0(d2_adj_5711[41]), .B0(d1_adj_5710[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[42]), .B1(d1_adj_5710[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16025), .COUT(n16026), .S0(n168_adj_5638), 
          .S1(n165_adj_5637));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_15 (.A0(d6_adj_5715[48]), .B0(cout_adj_5464), 
          .C0(n147_adj_4901), .D0(n25_adj_2798), .A1(d6_adj_5715[49]), 
          .B1(cout_adj_5464), .C1(n144_adj_4900), .D1(n24_adj_4556), .CIN(n16180), 
          .COUT(n16181), .S0(d7_71__N_1531_adj_5743[48]), .S1(d7_71__N_1531_adj_5743[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_27 (.A0(d_d9_adj_5722[61]), .B0(d9_adj_5721[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[62]), .B1(d9_adj_5721[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16102), .COUT(n16103), .S0(n106_adj_5587), 
          .S1(n103_adj_5586));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_27.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_27.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_25 (.A0(d_d9_adj_5722[59]), .B0(d9_adj_5721[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[60]), .B1(d9_adj_5721[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16101), .COUT(n16102), .S0(n112_adj_5589), 
          .S1(n109_adj_5588));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_25.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_25.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_23 (.A0(d_d9_adj_5722[57]), .B0(d9_adj_5721[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[58]), .B1(d9_adj_5721[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16100), .COUT(n16101), .S0(n118_adj_5591), 
          .S1(n115_adj_5590));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_23.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_23.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_21 (.A0(d_d9_adj_5722[55]), .B0(d9_adj_5721[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[56]), .B1(d9_adj_5721[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16099), .COUT(n16100));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_21.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_21.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_19 (.A0(d_d9_adj_5722[53]), .B0(d9_adj_5721[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[54]), .B1(d9_adj_5721[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16098), .COUT(n16099));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_19.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_19.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_19.INJECT1_1 = "NO";
    CCU2C add_3659_3 (.A0(d_out_d_11__N_1874[17]), .B0(ISquare[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16370), .COUT(n16371), .S1(n60));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3659_3.INIT0 = 16'h666a;
    defparam add_3659_3.INIT1 = 16'h555f;
    defparam add_3659_3.INJECT1_0 = "NO";
    defparam add_3659_3.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_17 (.A0(d_d9_adj_5722[51]), .B0(d9_adj_5721[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[52]), .B1(d9_adj_5721[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16097), .COUT(n16098));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_17.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_17.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_15 (.A0(d_d9_adj_5722[49]), .B0(d9_adj_5721[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[50]), .B1(d9_adj_5721[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16096), .COUT(n16097));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_15.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_15.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_26 (.A0(d2_adj_5711[59]), .B0(d1_adj_5710[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[60]), .B1(d1_adj_5710[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16034), .COUT(n16035), .S0(n114_adj_5620), 
          .S1(n111_adj_5619));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_13 (.A0(d_d9_adj_5722[47]), .B0(d9_adj_5721[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[48]), .B1(d9_adj_5721[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16095), .COUT(n16096));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_13.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_13.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_11 (.A0(d_d9_adj_5722[45]), .B0(d9_adj_5721[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[46]), .B1(d9_adj_5721[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16094), .COUT(n16095));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_13 (.A0(d6_adj_5715[46]), .B0(cout_adj_5464), 
          .C0(n153_adj_4903), .D0(n27_adj_4750), .A1(d6_adj_5715[47]), 
          .B1(cout_adj_5464), .C1(n150_adj_4902), .D1(n26_adj_2797), .CIN(n16179), 
          .COUT(n16180), .S0(d7_71__N_1531_adj_5743[46]), .S1(d7_71__N_1531_adj_5743[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_13.INJECT1_1 = "NO";
    FD1S3AX phase_accum_e3_i0_i0 (.D(n321), .CK(clk_80mhz), .Q(phase_accum_adj_5702[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i0.GSR = "ENABLED";
    CCU2C add_3659_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16370));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3659_1.INIT0 = 16'h0000;
    defparam add_3659_1.INIT1 = 16'haaaf;
    defparam add_3659_1.INJECT1_0 = "NO";
    defparam add_3659_1.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_9 (.A0(d_d9_adj_5722[43]), .B0(d9_adj_5721[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[44]), .B1(d9_adj_5721[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16093), .COUT(n16094));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_11 (.A0(d6_adj_5715[44]), .B0(cout_adj_5464), 
          .C0(n159_adj_4905), .D0(n29_adj_4748), .A1(d6_adj_5715[45]), 
          .B1(cout_adj_5464), .C1(n156_adj_4904), .D1(n28_adj_4749), .CIN(n16178), 
          .COUT(n16179), .S0(d7_71__N_1531_adj_5743[44]), .S1(d7_71__N_1531_adj_5743[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_7 (.A0(d_d9_adj_5722[41]), .B0(d9_adj_5721[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[42]), .B1(d9_adj_5721[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16092), .COUT(n16093));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_5 (.A0(d_d9_adj_5722[39]), .B0(d9_adj_5721[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[40]), .B1(d9_adj_5721[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16091), .COUT(n16092));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_3 (.A0(d_d9_adj_5722[37]), .B0(d9_adj_5721[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[38]), .B1(d9_adj_5721[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16090), .COUT(n16091));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_1409_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1409_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9_adj_5722[36]), .B1(d9_adj_5721[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16090));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1409_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1409_add_4_1.INIT1 = 16'h9995;
    defparam _add_1_1409_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1409_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_31 (.A0(d6_adj_5715[64]), .B0(cout_adj_5464), 
          .C0(n99_adj_4885), .D0(n9_adj_4755), .A1(d6_adj_5715[65]), .B1(cout_adj_5464), 
          .C1(n96_adj_4884), .D1(n8_adj_4756), .CIN(n16188), .COUT(n16189), 
          .S0(d7_71__N_1531_adj_5743[64]), .S1(d7_71__N_1531_adj_5743[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_29 (.A0(d6_adj_5715[62]), .B0(cout_adj_5464), 
          .C0(n105_adj_4887), .D0(n11_adj_4753), .A1(d6_adj_5715[63]), 
          .B1(cout_adj_5464), .C1(n102_adj_4886), .D1(n10_adj_4754), .CIN(n16187), 
          .COUT(n16188), .S0(d7_71__N_1531_adj_5743[62]), .S1(d7_71__N_1531_adj_5743[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_27 (.A0(d6_adj_5715[60]), .B0(cout_adj_5464), 
          .C0(n111_adj_4889), .D0(n13_adj_4744), .A1(d6_adj_5715[61]), 
          .B1(cout_adj_5464), .C1(n108_adj_4888), .D1(n12_adj_4751), .CIN(n16186), 
          .COUT(n16187), .S0(d7_71__N_1531_adj_5743[60]), .S1(d7_71__N_1531_adj_5743[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_27.INJECT1_1 = "NO";
    IB RFIn_pad (.I(RFIn), .O(RFIn_c));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(42[22:26])
    IB i_Rx_Serial_pad (.I(i_Rx_Serial), .O(i_Rx_Serial_c));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(41[22:33])
    CCU2C _add_1_1418_add_4_25 (.A0(d6_adj_5715[58]), .B0(cout_adj_5464), 
          .C0(n117_adj_4891), .D0(n15_adj_2794), .A1(d6_adj_5715[59]), 
          .B1(cout_adj_5464), .C1(n114_adj_4890), .D1(n14_adj_4732), .CIN(n16185), 
          .COUT(n16186), .S0(d7_71__N_1531_adj_5743[58]), .S1(d7_71__N_1531_adj_5743[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_25.INJECT1_1 = "NO";
    IB clk_25mhz_pad (.I(clk_25mhz), .O(clk_25mhz_c));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(40[22:31])
    OB CIC_out_clkSin_pad (.I(GND_net), .O(CIC_out_clkSin));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(58[22:36])
    OB sin_out_pad (.I(GND_net), .O(sin_out));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(57[22:29])
    CCU2C _add_1_1418_add_4_23 (.A0(d6_adj_5715[56]), .B0(cout_adj_5464), 
          .C0(n123_adj_4893), .D0(n17_adj_4595), .A1(d6_adj_5715[57]), 
          .B1(cout_adj_5464), .C1(n120_adj_4892), .D1(n16_adj_4731), .CIN(n16184), 
          .COUT(n16185), .S0(d7_71__N_1531_adj_5743[56]), .S1(d7_71__N_1531_adj_5743[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_23.INJECT1_1 = "NO";
    OB sinGen_pad (.I(sinGen_c), .O(sinGen));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(56[22:28])
    OB PWMOutN4_pad (.I(PWMOutN4_c), .O(PWMOutN4));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(55[22:30])
    CCU2C _add_1_1544_add_4_24 (.A0(d2_adj_5711[57]), .B0(d1_adj_5710[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[58]), .B1(d1_adj_5710[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16033), .COUT(n16034), .S0(n120_adj_5622), 
          .S1(n117_adj_5621));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_24.INJECT1_1 = "NO";
    OB PWMOutN3_pad (.I(PWMOutN4_c), .O(PWMOutN3));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(54[22:30])
    OB PWMOutN2_pad (.I(PWMOutN4_c), .O(PWMOutN2));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(53[22:30])
    CCU2C _add_1_1544_add_4_22 (.A0(d2_adj_5711[55]), .B0(d1_adj_5710[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[56]), .B1(d1_adj_5710[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16032), .COUT(n16033), .S0(n126_adj_5624), 
          .S1(n123_adj_5623));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_4 (.A0(d5_adj_5714[37]), .B0(d4_adj_5713[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[38]), .B1(d4_adj_5713[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16153), .COUT(n16154), .S0(n180_adj_5572), 
          .S1(n177_adj_5571));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_4.INJECT1_1 = "NO";
    OB PWMOutN1_pad (.I(PWMOutN4_c), .O(PWMOutN1));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(52[22:30])
    CCU2C add_3661_11 (.A0(ISquare[31]), .B0(n17828), .C0(n17826), .D0(VCC_net), 
          .A1(ISquare[31]), .B1(n17828), .C1(n17826), .D1(VCC_net), 
          .CIN(n16364), .S0(n29_adj_4752), .S1(d_out_d_11__N_1874[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3661_11.INIT0 = 16'he1e1;
    defparam add_3661_11.INIT1 = 16'he1e1;
    defparam add_3661_11.INJECT1_0 = "NO";
    defparam add_3661_11.INJECT1_1 = "NO";
    CCU2C add_3661_9 (.A0(n17826), .B0(ISquare[31]), .C0(ISquare[23]), 
          .D0(ISquare[22]), .A1(n23_adj_5022), .B1(n14967), .C1(n213), 
          .D1(ISquare[31]), .CIN(n16363), .COUT(n16364), .S0(n35_adj_4742), 
          .S1(n32_adj_4743));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3661_9.INIT0 = 16'h6665;
    defparam add_3661_9.INIT1 = 16'h556a;
    defparam add_3661_9.INJECT1_0 = "NO";
    defparam add_3661_9.INJECT1_1 = "NO";
    CCU2C add_3661_7 (.A0(n32_adj_5023), .B0(ISquare[31]), .C0(ISquare[23]), 
          .D0(ISquare[22]), .A1(n17828), .B1(ISquare[31]), .C1(ISquare[23]), 
          .D1(ISquare[22]), .CIN(n16362), .COUT(n16363), .S0(n41), .S1(n38));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3661_7.INIT0 = 16'h999a;
    defparam add_3661_7.INIT1 = 16'haaa9;
    defparam add_3661_7.INJECT1_0 = "NO";
    defparam add_3661_7.INJECT1_1 = "NO";
    CCU2C add_3661_5 (.A0(ISquare[22]), .B0(ISquare[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[23]), .B1(ISquare[22]), .C1(ISquare[31]), 
          .D1(n14967), .CIN(n16361), .COUT(n16362), .S0(n47), .S1(n44));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3661_5.INIT0 = 16'h9999;
    defparam add_3661_5.INIT1 = 16'heee1;
    defparam add_3661_5.INJECT1_0 = "NO";
    defparam add_3661_5.INJECT1_1 = "NO";
    CCU2C add_3661_3 (.A0(ISquare[31]), .B0(n17828), .C0(ISquare[20]), 
          .D0(VCC_net), .A1(ISquare[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16360), .COUT(n16361), .S1(n50));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3661_3.INIT0 = 16'he1e1;
    defparam add_3661_3.INIT1 = 16'h555f;
    defparam add_3661_3.INJECT1_0 = "NO";
    defparam add_3661_3.INJECT1_1 = "NO";
    CCU2C add_3661_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(ISquare[22]), .B1(ISquare[23]), .C1(n213), .D1(ISquare[31]), 
          .COUT(n16360));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3661_1.INIT0 = 16'h0000;
    defparam add_3661_1.INIT1 = 16'h001f;
    defparam add_3661_1.INJECT1_0 = "NO";
    defparam add_3661_1.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_37 (.A0(d3[70]), .B0(cout_adj_4267), .C0(n81_adj_5250), 
          .D0(d4[70]), .A1(d3[71]), .B1(cout_adj_4267), .C1(n78_adj_5249), 
          .D1(d4[71]), .CIN(n16083), .S0(d4_71__N_634[70]), .S1(d4_71__N_634[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_6 (.A0(d5_adj_5714[39]), .B0(d4_adj_5713[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[40]), .B1(d4_adj_5713[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16154), .COUT(n16155), .S0(n174_adj_5570), 
          .S1(n171_adj_5569));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_6.INJECT1_1 = "NO";
    OB PWMOutP4_pad (.I(PWMOutP4_c), .O(PWMOutP4));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(51[22:30])
    CCU2C add_3662_17 (.A0(ISquare[31]), .B0(n917), .C0(GND_net), .D0(VCC_net), 
          .A1(n916), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16354), 
          .S1(d_out_d_11__N_2401[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3662_17.INIT0 = 16'h666a;
    defparam add_3662_17.INIT1 = 16'haaa0;
    defparam add_3662_17.INJECT1_0 = "NO";
    defparam add_3662_17.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_36 (.A0(d5_adj_5714[69]), .B0(d4_adj_5713[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[70]), .B1(d4_adj_5713[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16169), .COUT(n16170), .S0(n84_adj_5540), 
          .S1(n81_adj_5539));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_10 (.A0(d5_adj_5714[43]), .B0(d4_adj_5713[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[44]), .B1(d4_adj_5713[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16156), .COUT(n16157), .S0(n162_adj_5566), 
          .S1(n159_adj_5565));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_10.INJECT1_1 = "NO";
    CCU2C add_3662_15 (.A0(ISquare[31]), .B0(n919), .C0(GND_net), .D0(VCC_net), 
          .A1(ISquare[31]), .B1(n918), .C1(GND_net), .D1(VCC_net), .CIN(n16353), 
          .COUT(n16354));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3662_15.INIT0 = 16'h666a;
    defparam add_3662_15.INIT1 = 16'h666a;
    defparam add_3662_15.INJECT1_0 = "NO";
    defparam add_3662_15.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_20 (.A0(d2_adj_5711[53]), .B0(d1_adj_5710[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[54]), .B1(d1_adj_5710[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16031), .COUT(n16032), .S0(n132_adj_5626), 
          .S1(n129_adj_5625));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_18 (.A0(d2_adj_5711[51]), .B0(d1_adj_5710[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[52]), .B1(d1_adj_5710[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16030), .COUT(n16031), .S0(n138_adj_5628), 
          .S1(n135_adj_5627));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_21 (.A0(d4[54]), .B0(cout_adj_2810), .C0(n129_adj_5302), 
          .D0(d5[54]), .A1(d4[55]), .B1(cout_adj_2810), .C1(n126_adj_5301), 
          .D1(d5[55]), .CIN(n16053), .COUT(n16054), .S0(d5_71__N_706[54]), 
          .S1(d5_71__N_706[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_21 (.A0(d6_adj_5715[54]), .B0(cout_adj_5464), 
          .C0(n129_adj_4895), .D0(n19_adj_4579), .A1(d6_adj_5715[55]), 
          .B1(cout_adj_5464), .C1(n126_adj_4894), .D1(n18_adj_4580), .CIN(n16183), 
          .COUT(n16184), .S0(d7_71__N_1531_adj_5743[54]), .S1(d7_71__N_1531_adj_5743[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_35 (.A0(d3[68]), .B0(cout_adj_4267), .C0(n87_adj_5252), 
          .D0(d4[68]), .A1(d3[69]), .B1(cout_adj_4267), .C1(n84_adj_5251), 
          .D1(d4[69]), .CIN(n16082), .COUT(n16083), .S0(d4_71__N_634[68]), 
          .S1(d4_71__N_634[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_19 (.A0(d4[52]), .B0(cout_adj_2810), .C0(n135_adj_5304), 
          .D0(d5[52]), .A1(d4[53]), .B1(cout_adj_2810), .C1(n132_adj_5303), 
          .D1(d5[53]), .CIN(n16052), .COUT(n16053), .S0(d5_71__N_706[52]), 
          .S1(d5_71__N_706[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_17 (.A0(d4[50]), .B0(cout_adj_2810), .C0(n141_adj_5306), 
          .D0(d5[50]), .A1(d4[51]), .B1(cout_adj_2810), .C1(n138_adj_5305), 
          .D1(d5[51]), .CIN(n16051), .COUT(n16052), .S0(d5_71__N_706[50]), 
          .S1(d5_71__N_706[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d5_adj_5714[36]), .B1(d4_adj_5713[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16153), .S1(n183_adj_5573));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1553_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_16 (.A0(d2_adj_5711[49]), .B0(d1_adj_5710[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[50]), .B1(d1_adj_5710[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16029), .COUT(n16030), .S0(n144_adj_5630), 
          .S1(n141_adj_5629));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_33 (.A0(d2[66]), .B0(cout), .C0(n93_adj_5159), 
          .D0(d3[66]), .A1(d2[67]), .B1(cout), .C1(n90_adj_5158), .D1(d3[67]), 
          .CIN(n16149), .COUT(n16150), .S0(d3_71__N_562[66]), .S1(d3_71__N_562[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_27 (.A0(d2[60]), .B0(cout), .C0(n111_adj_5165), 
          .D0(d3[60]), .A1(d2[61]), .B1(cout), .C1(n108_adj_5164), .D1(d3[61]), 
          .CIN(n16146), .COUT(n16147), .S0(d3_71__N_562[60]), .S1(d3_71__N_562[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_33 (.A0(d3[66]), .B0(cout_adj_4267), .C0(n93_adj_5254), 
          .D0(d4[66]), .A1(d3[67]), .B1(cout_adj_4267), .C1(n90_adj_5253), 
          .D1(d4[67]), .CIN(n16081), .COUT(n16082), .S0(d4_71__N_634[66]), 
          .S1(d4_71__N_634[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_31 (.A0(d2[64]), .B0(cout), .C0(n99_adj_5161), 
          .D0(d3[64]), .A1(d2[65]), .B1(cout), .C1(n96_adj_5160), .D1(d3[65]), 
          .CIN(n16148), .COUT(n16149), .S0(d3_71__N_562[64]), .S1(d3_71__N_562[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_37 (.A0(d2[70]), .B0(cout), .C0(n81_adj_5155), 
          .D0(d3[70]), .A1(d2[71]), .B1(cout), .C1(n78_adj_5154), .D1(d3[71]), 
          .CIN(n16151), .S0(d3_71__N_562[70]), .S1(d3_71__N_562[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_29 (.A0(d2[62]), .B0(cout), .C0(n105_adj_5163), 
          .D0(d3[62]), .A1(d2[63]), .B1(cout), .C1(n102_adj_5162), .D1(d3[63]), 
          .CIN(n16147), .COUT(n16148), .S0(d3_71__N_562[62]), .S1(d3_71__N_562[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_25 (.A0(d2[58]), .B0(cout), .C0(n117_adj_5167), 
          .D0(d3[58]), .A1(d2[59]), .B1(cout), .C1(n114_adj_5166), .D1(d3[59]), 
          .CIN(n16145), .COUT(n16146), .S0(d3_71__N_562[58]), .S1(d3_71__N_562[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_35 (.A0(d2[68]), .B0(cout), .C0(n87_adj_5157), 
          .D0(d3[68]), .A1(d2[69]), .B1(cout), .C1(n84_adj_5156), .D1(d3[69]), 
          .CIN(n16150), .COUT(n16151), .S0(d3_71__N_562[68]), .S1(d3_71__N_562[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_34 (.A0(d_d_tmp[31]), .B0(d_tmp[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[32]), .B1(d_tmp[32]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15620), .COUT(n15621), .S0(d6_71__N_1459[31]), 
          .S1(d6_71__N_1459[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_32 (.A0(d_d_tmp[29]), .B0(d_tmp[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[30]), .B1(d_tmp[30]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15619), .COUT(n15620), .S0(d6_71__N_1459[29]), 
          .S1(d6_71__N_1459[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_30 (.A0(d_d_tmp[27]), .B0(d_tmp[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[28]), .B1(d_tmp[28]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15618), .COUT(n15619), .S0(d6_71__N_1459[27]), 
          .S1(d6_71__N_1459[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_28 (.A0(d_d_tmp[25]), .B0(d_tmp[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[26]), .B1(d_tmp[26]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15617), .COUT(n15618), .S0(d6_71__N_1459[25]), 
          .S1(d6_71__N_1459[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_31 (.A0(d3[64]), .B0(cout_adj_4267), .C0(n99_adj_5256), 
          .D0(d4[64]), .A1(d3[65]), .B1(cout_adj_4267), .C1(n96_adj_5255), 
          .D1(d4[65]), .CIN(n16080), .COUT(n16081), .S0(d4_71__N_634[64]), 
          .S1(d4_71__N_634[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_26 (.A0(d_d_tmp[23]), .B0(d_tmp[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[24]), .B1(d_tmp[24]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15616), .COUT(n15617), .S0(d6_71__N_1459[23]), 
          .S1(d6_71__N_1459[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_26.INJECT1_1 = "NO";
    PFUMX i2666 (.BLUT(n11980), .ALUT(n12253), .C0(n17389), .Z(n12571));
    CCU2C _add_1_1457_add_4_29 (.A0(d3[62]), .B0(cout_adj_4267), .C0(n105_adj_5258), 
          .D0(d4[62]), .A1(d3[63]), .B1(cout_adj_4267), .C1(n102_adj_5257), 
          .D1(d4[63]), .CIN(n16079), .COUT(n16080), .S0(d4_71__N_634[62]), 
          .S1(d4_71__N_634[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_27 (.A0(d3[60]), .B0(cout_adj_4267), .C0(n111_adj_5260), 
          .D0(d4[60]), .A1(d3[61]), .B1(cout_adj_4267), .C1(n108_adj_5259), 
          .D1(d4[61]), .CIN(n16078), .COUT(n16079), .S0(d4_71__N_634[60]), 
          .S1(d4_71__N_634[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_15 (.A0(d4[48]), .B0(cout_adj_2810), .C0(n147_adj_5308), 
          .D0(d5[48]), .A1(d4[49]), .B1(cout_adj_2810), .C1(n144_adj_5307), 
          .D1(d5[49]), .CIN(n16050), .COUT(n16051), .S0(d5_71__N_706[48]), 
          .S1(d5_71__N_706[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_25 (.A0(d3[58]), .B0(cout_adj_4267), .C0(n117_adj_5262), 
          .D0(d4[58]), .A1(d3[59]), .B1(cout_adj_4267), .C1(n114_adj_5261), 
          .D1(d4[59]), .CIN(n16077), .COUT(n16078), .S0(d4_71__N_634[58]), 
          .S1(d4_71__N_634[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_23 (.A0(d2[56]), .B0(cout), .C0(n123_adj_5169), 
          .D0(d3[56]), .A1(d2[57]), .B1(cout), .C1(n120_adj_5168), .D1(d3[57]), 
          .CIN(n16144), .COUT(n16145), .S0(d3_71__N_562[56]), .S1(d3_71__N_562[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_21 (.A0(d2[54]), .B0(cout), .C0(n129_adj_5171), 
          .D0(d3[54]), .A1(d2[55]), .B1(cout), .C1(n126_adj_5170), .D1(d3[55]), 
          .CIN(n16143), .COUT(n16144), .S0(d3_71__N_562[54]), .S1(d3_71__N_562[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_19 (.A0(d2[52]), .B0(cout), .C0(n135_adj_5173), 
          .D0(d3[52]), .A1(d2[53]), .B1(cout), .C1(n132_adj_5172), .D1(d3[53]), 
          .CIN(n16142), .COUT(n16143), .S0(d3_71__N_562[52]), .S1(d3_71__N_562[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_13 (.A0(d4[46]), .B0(cout_adj_2810), .C0(n153_adj_5310), 
          .D0(d5[46]), .A1(d4[47]), .B1(cout_adj_2810), .C1(n150_adj_5309), 
          .D1(d5[47]), .CIN(n16049), .COUT(n16050), .S0(d5_71__N_706[46]), 
          .S1(d5_71__N_706[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_17 (.A0(d2[50]), .B0(cout), .C0(n141_adj_5175), 
          .D0(d3[50]), .A1(d2[51]), .B1(cout), .C1(n138_adj_5174), .D1(d3[51]), 
          .CIN(n16141), .COUT(n16142), .S0(d3_71__N_562[50]), .S1(d3_71__N_562[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_13 (.A0(d2[46]), .B0(cout), .C0(n153_adj_5179), 
          .D0(d3[46]), .A1(d2[47]), .B1(cout), .C1(n150_adj_5178), .D1(d3[47]), 
          .CIN(n16139), .COUT(n16140), .S0(d3_71__N_562[46]), .S1(d3_71__N_562[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_13.INJECT1_1 = "NO";
    PFUMX i2662 (.BLUT(n11978), .ALUT(n12251), .C0(n17389), .Z(n12567));
    CCU2C _add_1_1601_add_4_24 (.A0(d_d_tmp[21]), .B0(d_tmp[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[22]), .B1(d_tmp[22]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15615), .COUT(n15616), .S0(d6_71__N_1459[21]), 
          .S1(d6_71__N_1459[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_24.INJECT1_1 = "NO";
    FD1P3AX phase_inc_carrGen_i0_i0 (.D(n1994), .SP(clk_80mhz_enable_23), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i0.GSR = "ENABLED";
    CCU2C _add_1_1553_add_4_20 (.A0(d5_adj_5714[53]), .B0(d4_adj_5713[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[54]), .B1(d4_adj_5713[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16161), .COUT(n16162), .S0(n132_adj_5556), 
          .S1(n129_adj_5555));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_14 (.A0(d2_adj_5711[47]), .B0(d1_adj_5710[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[48]), .B1(d1_adj_5710[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16028), .COUT(n16029), .S0(n150_adj_5632), 
          .S1(n147_adj_5631));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_14.INJECT1_1 = "NO";
    OB PWMOutP3_pad (.I(PWMOutP4_c), .O(PWMOutP3));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(50[22:30])
    OB PWMOutP2_pad (.I(PWMOutP4_c), .O(PWMOutP2));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(49[22:30])
    OB PWMOutP1_pad (.I(PWMOutP4_c), .O(PWMOutP1));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(48[22:30])
    OB PWMOut_pad (.I(PWMOutP4_c), .O(PWMOut));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(47[22:28])
    OB DiffOut_pad (.I(DiffOut_c), .O(DiffOut));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(46[22:29])
    OB XOut_pad (.I(GND_net), .O(XOut));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(45[22:26])
    OB led_pad_0 (.I(led_c_0), .O(led[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(44[22:25])
    OB led_pad_1 (.I(led_c_1), .O(led[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(44[22:25])
    OB led_pad_2 (.I(led_c_2), .O(led[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(44[22:25])
    OB led_pad_3 (.I(led_c_3), .O(led[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(44[22:25])
    CCU2C _add_1_1553_add_4_30 (.A0(d5_adj_5714[63]), .B0(d4_adj_5713[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[64]), .B1(d4_adj_5713[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16166), .COUT(n16167), .S0(n102_adj_5546), 
          .S1(n99_adj_5545));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_16 (.A0(d5_adj_5714[49]), .B0(d4_adj_5713[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[50]), .B1(d4_adj_5713[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16159), .COUT(n16160), .S0(n144_adj_5560), 
          .S1(n141_adj_5559));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_16.INJECT1_1 = "NO";
    OB led_pad_4 (.I(led_c_4), .O(led[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(44[22:25])
    FD1P3IX phase_inc_carrGen_i0_i58 (.D(n12615), .SP(o_Rx_DV), .CD(n17822), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[58]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i58.GSR = "ENABLED";
    CCU2C add_3662_13 (.A0(n921), .B0(n14967), .C0(n213), .D0(ISquare[31]), 
          .A1(n920), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16352), 
          .COUT(n16353));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3662_13.INIT0 = 16'h556a;
    defparam add_3662_13.INIT1 = 16'haaa0;
    defparam add_3662_13.INJECT1_0 = "NO";
    defparam add_3662_13.INJECT1_1 = "NO";
    FD1P3IX phase_inc_carrGen_i0_i56 (.D(n12613), .SP(o_Rx_DV), .CD(n17822), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[56]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i56.GSR = "ENABLED";
    CCU2C add_3662_11 (.A0(d_out_d_11__N_1876[17]), .B0(n923), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), .B1(n922), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16351), .COUT(n16352));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3662_11.INIT0 = 16'h9995;
    defparam add_3662_11.INIT1 = 16'h9995;
    defparam add_3662_11.INJECT1_0 = "NO";
    defparam add_3662_11.INJECT1_1 = "NO";
    CCU2C add_3662_9 (.A0(d_out_d_11__N_1880[17]), .B0(n925), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n924), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16350), .COUT(n16351));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3662_9.INIT0 = 16'h9995;
    defparam add_3662_9.INIT1 = 16'h9995;
    defparam add_3662_9.INJECT1_0 = "NO";
    defparam add_3662_9.INJECT1_1 = "NO";
    CCU2C add_3662_7 (.A0(d_out_d_11__N_1884[17]), .B0(n927), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n926), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16349), .COUT(n16350));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3662_7.INIT0 = 16'h9995;
    defparam add_3662_7.INIT1 = 16'h9995;
    defparam add_3662_7.INJECT1_0 = "NO";
    defparam add_3662_7.INJECT1_1 = "NO";
    CCU2C add_3662_5 (.A0(d_out_d_11__N_1888[17]), .B0(n929), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), .B1(n928), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16348), .COUT(n16349));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3662_5.INIT0 = 16'h9995;
    defparam add_3662_5.INIT1 = 16'h9995;
    defparam add_3662_5.INJECT1_0 = "NO";
    defparam add_3662_5.INJECT1_1 = "NO";
    CCU2C add_3662_3 (.A0(d_out_d_11__N_1892[17]), .B0(n931), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1890[17]), .B1(n930), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16347), .COUT(n16348));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3662_3.INIT0 = 16'h9995;
    defparam add_3662_3.INIT1 = 16'h9995;
    defparam add_3662_3.INJECT1_0 = "NO";
    defparam add_3662_3.INJECT1_1 = "NO";
    CCU2C add_3662_1 (.A0(ISquare[0]), .B0(GND_net), .C0(GND_net), .D0(ISquare[0]), 
          .A1(d_out_d_11__N_1892[17]), .B1(ISquare[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16347));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3662_1.INIT0 = 16'h000A;
    defparam add_3662_1.INIT1 = 16'h666a;
    defparam add_3662_1.INJECT1_0 = "NO";
    defparam add_3662_1.INJECT1_1 = "NO";
    CCU2C add_3663_19 (.A0(d_out_d_11__N_1879), .B0(d_out_d_11__N_1880[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1879), .B1(d_out_d_11__N_1880[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16345), .S0(n45_adj_5190), 
          .S1(d_out_d_11__N_1882[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3663_19.INIT0 = 16'h666a;
    defparam add_3663_19.INIT1 = 16'h666a;
    defparam add_3663_19.INJECT1_0 = "NO";
    defparam add_3663_19.INJECT1_1 = "NO";
    CCU2C add_3663_17 (.A0(d_out_d_11__N_1880[17]), .B0(n44_adj_4838), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n41_adj_4837), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16344), .COUT(n16345), .S0(n51_adj_5192), 
          .S1(n48_adj_5191));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3663_17.INIT0 = 16'h9995;
    defparam add_3663_17.INIT1 = 16'h9995;
    defparam add_3663_17.INJECT1_0 = "NO";
    defparam add_3663_17.INJECT1_1 = "NO";
    CCU2C add_3663_15 (.A0(d_out_d_11__N_1880[17]), .B0(n50_adj_4840), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n47_adj_4839), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16343), .COUT(n16344), .S0(n57_adj_5194), 
          .S1(n54_adj_5193));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3663_15.INIT0 = 16'h9995;
    defparam add_3663_15.INIT1 = 16'h9995;
    defparam add_3663_15.INJECT1_0 = "NO";
    defparam add_3663_15.INJECT1_1 = "NO";
    CCU2C add_3663_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1880[17]), .C0(n56), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n53), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16342), .COUT(n16343), .S0(n63_adj_5196), 
          .S1(n60_adj_5195));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3663_13.INIT0 = 16'h6969;
    defparam add_3663_13.INIT1 = 16'h9995;
    defparam add_3663_13.INJECT1_0 = "NO";
    defparam add_3663_13.INJECT1_1 = "NO";
    CCU2C add_3663_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1880[17]), .C0(n62), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1880[17]), 
          .C1(n59), .D1(VCC_net), .CIN(n16341), .COUT(n16342), .S0(n69_adj_5198), 
          .S1(n66_adj_5197));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3663_11.INIT0 = 16'h6969;
    defparam add_3663_11.INIT1 = 16'h6969;
    defparam add_3663_11.INJECT1_0 = "NO";
    defparam add_3663_11.INJECT1_1 = "NO";
    CCU2C add_3663_9 (.A0(d_out_d_11__N_1880[17]), .B0(n17826), .C0(n68), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n65_adj_4841), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16340), .COUT(n16341), .S0(n75_adj_5200), 
          .S1(n72_adj_5199));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3663_9.INIT0 = 16'h6969;
    defparam add_3663_9.INIT1 = 16'h9995;
    defparam add_3663_9.INJECT1_0 = "NO";
    defparam add_3663_9.INJECT1_1 = "NO";
    FD1P3IX phase_inc_carrGen_i0_i55 (.D(n12611), .SP(o_Rx_DV), .CD(n17822), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i55.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i54 (.D(n12609), .SP(o_Rx_DV), .CD(n17822), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[54]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i54.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i53 (.D(n12607), .SP(o_Rx_DV), .CD(n17822), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i53.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i51 (.D(n12605), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i51.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i50 (.D(n12603), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[50]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i50.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i49 (.D(n12601), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i49.GSR = "ENABLED";
    CCU2C _add_1_1544_add_4_6 (.A0(d2_adj_5711[39]), .B0(d1_adj_5710[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[40]), .B1(d1_adj_5710[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16024), .COUT(n16025), .S0(n174_adj_5640), 
          .S1(n171_adj_5639));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_6.INJECT1_1 = "NO";
    FD1P3IX phase_inc_carrGen_i0_i48 (.D(n12599), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[48]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i48.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i46 (.D(n12597), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[46]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i46.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i40 (.D(n12593), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[40]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i40.GSR = "ENABLED";
    CCU2C add_3663_7 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1880[17]), 
          .C0(n74), .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), .B1(d_out_d_11__N_1880[17]), 
          .C1(n71), .D1(VCC_net), .CIN(n16339), .COUT(n16340), .S0(n81_adj_5202), 
          .S1(n78_adj_5201));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3663_7.INIT0 = 16'h9696;
    defparam add_3663_7.INIT1 = 16'h9696;
    defparam add_3663_7.INJECT1_0 = "NO";
    defparam add_3663_7.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i63 (.D(phase_inc_carrGen[63]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i63.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i62 (.D(phase_inc_carrGen[62]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[62]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i62.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i61 (.D(phase_inc_carrGen[61]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i61.GSR = "ENABLED";
    CCU2C _add_1_1601_add_4_22 (.A0(d_d_tmp[19]), .B0(d_tmp[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[20]), .B1(d_tmp[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15614), .COUT(n15615), .S0(d6_71__N_1459[19]), 
          .S1(d6_71__N_1459[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_22.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i60 (.D(phase_inc_carrGen[60]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[60]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i60.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i59 (.D(phase_inc_carrGen[59]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i59.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i58 (.D(phase_inc_carrGen[58]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[58]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i58.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i57 (.D(phase_inc_carrGen[57]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i57.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i56 (.D(phase_inc_carrGen[56]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[56]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i56.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i55 (.D(phase_inc_carrGen[55]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i55.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i54 (.D(phase_inc_carrGen[54]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[54]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i54.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i53 (.D(phase_inc_carrGen[53]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i53.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i52 (.D(phase_inc_carrGen[52]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[52]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i52.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i51 (.D(phase_inc_carrGen[51]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i51.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i50 (.D(phase_inc_carrGen[50]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[50]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i50.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i49 (.D(phase_inc_carrGen[49]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i49.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i48 (.D(phase_inc_carrGen[48]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[48]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i48.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i47 (.D(phase_inc_carrGen[47]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i47.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i46 (.D(phase_inc_carrGen[46]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[46]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i46.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i45 (.D(phase_inc_carrGen[45]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i45.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i44 (.D(phase_inc_carrGen[44]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[44]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i44.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i43 (.D(phase_inc_carrGen[43]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i43.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i42 (.D(phase_inc_carrGen[42]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[42]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i42.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i41 (.D(phase_inc_carrGen[41]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i41.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i40 (.D(phase_inc_carrGen[40]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[40]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i40.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i39 (.D(phase_inc_carrGen[39]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i39.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i38 (.D(phase_inc_carrGen[38]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[38]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i38.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i37 (.D(phase_inc_carrGen[37]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i37.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i36 (.D(phase_inc_carrGen[36]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[36]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i36.GSR = "ENABLED";
    CCU2C _add_1_1553_add_4_18 (.A0(d5_adj_5714[51]), .B0(d4_adj_5713[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[52]), .B1(d4_adj_5713[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16160), .COUT(n16161), .S0(n138_adj_5558), 
          .S1(n135_adj_5557));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_18.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i35 (.D(phase_inc_carrGen[35]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i35.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i34 (.D(phase_inc_carrGen[34]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i34.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i33 (.D(phase_inc_carrGen[33]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i33.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i32 (.D(phase_inc_carrGen[32]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i32.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i31 (.D(phase_inc_carrGen[31]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i31.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i30 (.D(phase_inc_carrGen[30]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i30.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i29 (.D(phase_inc_carrGen[29]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i29.GSR = "ENABLED";
    CCU2C _add_1_1601_add_4_20 (.A0(d_d_tmp[17]), .B0(d_tmp[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[18]), .B1(d_tmp[18]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15613), .COUT(n15614), .S0(d6_71__N_1459[17]), 
          .S1(d6_71__N_1459[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_20.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i28 (.D(phase_inc_carrGen[28]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i28.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i27 (.D(phase_inc_carrGen[27]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i27.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i26 (.D(phase_inc_carrGen[26]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i26.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i25 (.D(phase_inc_carrGen[25]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i25.GSR = "ENABLED";
    CCU2C _add_1_1460_add_4_11 (.A0(d2[44]), .B0(cout), .C0(n159_adj_5181), 
          .D0(d3[44]), .A1(d2[45]), .B1(cout), .C1(n156_adj_5180), .D1(d3[45]), 
          .CIN(n16138), .COUT(n16139), .S0(d3_71__N_562[44]), .S1(d3_71__N_562[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_11.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i24 (.D(phase_inc_carrGen[24]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i24.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i23 (.D(phase_inc_carrGen[23]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i23.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i22 (.D(phase_inc_carrGen[22]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i22.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i21 (.D(phase_inc_carrGen[21]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i21.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i20 (.D(phase_inc_carrGen[20]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i20.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i19 (.D(phase_inc_carrGen[19]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i19.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i18 (.D(phase_inc_carrGen[18]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i18.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i17 (.D(phase_inc_carrGen[17]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i17.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i16 (.D(phase_inc_carrGen[16]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i16.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i15 (.D(phase_inc_carrGen[15]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i15.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i14 (.D(phase_inc_carrGen[14]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i14.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i13 (.D(phase_inc_carrGen[13]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i13.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i12 (.D(phase_inc_carrGen[12]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i12.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i11 (.D(phase_inc_carrGen[11]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i11.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i10 (.D(phase_inc_carrGen[10]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i10.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i9 (.D(phase_inc_carrGen[9]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i9.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i8 (.D(phase_inc_carrGen[8]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i8.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i7 (.D(phase_inc_carrGen[7]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i7.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i6 (.D(phase_inc_carrGen[6]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i6.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i5 (.D(phase_inc_carrGen[5]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i5.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i4 (.D(phase_inc_carrGen[4]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i4.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i3 (.D(phase_inc_carrGen[3]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i3.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i2 (.D(phase_inc_carrGen[2]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i2.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i1 (.D(phase_inc_carrGen[1]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen1_i1.GSR = "ENABLED";
    CCU2C _add_1_1457_add_4_23 (.A0(d3[56]), .B0(cout_adj_4267), .C0(n123_adj_5264), 
          .D0(d4[56]), .A1(d3[57]), .B1(cout_adj_4267), .C1(n120_adj_5263), 
          .D1(d4[57]), .CIN(n16076), .COUT(n16077), .S0(d4_71__N_634[56]), 
          .S1(d4_71__N_634[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_18 (.A0(d_d_tmp[15]), .B0(d_tmp[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[16]), .B1(d_tmp[16]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15612), .COUT(n15613), .S0(d6_71__N_1459[15]), 
          .S1(d6_71__N_1459[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_16 (.A0(d_d_tmp[13]), .B0(d_tmp[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[14]), .B1(d_tmp[14]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15611), .COUT(n15612), .S0(d6_71__N_1459[13]), 
          .S1(d6_71__N_1459[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_3 (.A0(d2[36]), .B0(cout), .C0(n183_adj_5189), 
          .D0(d3[36]), .A1(d2[37]), .B1(cout), .C1(n180_adj_5188), .D1(d3[37]), 
          .CIN(n16134), .COUT(n16135), .S0(d3_71__N_562[36]), .S1(d3_71__N_562[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_14 (.A0(d_d_tmp[11]), .B0(d_tmp[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[12]), .B1(d_tmp[12]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15610), .COUT(n15611), .S0(d6_71__N_1459[11]), 
          .S1(d6_71__N_1459[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_32 (.A0(d_d7[29]), .B0(d7[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[30]), .B1(d7[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16127), .COUT(n16128), .S0(d8_71__N_1603[29]), .S1(d8_71__N_1603[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_12 (.A0(d_d_tmp[9]), .B0(d_tmp[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[10]), .B1(d_tmp[10]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15609), .COUT(n15610), .S0(d6_71__N_1459[9]), 
          .S1(d6_71__N_1459[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_10 (.A0(d_d_tmp[7]), .B0(d_tmp[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[8]), .B1(d_tmp[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15608), .COUT(n15609), .S0(d6_71__N_1459[7]), 
          .S1(d6_71__N_1459[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_21 (.A0(d3[54]), .B0(cout_adj_4267), .C0(n129_adj_5266), 
          .D0(d4[54]), .A1(d3[55]), .B1(cout_adj_4267), .C1(n126_adj_5265), 
          .D1(d4[55]), .CIN(n16075), .COUT(n16076), .S0(d4_71__N_634[54]), 
          .S1(d4_71__N_634[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_8 (.A0(d_d_tmp[5]), .B0(d_tmp[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[6]), .B1(d_tmp[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15607), .COUT(n15608), .S0(d6_71__N_1459[5]), 
          .S1(d6_71__N_1459[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_6 (.A0(d_d_tmp[3]), .B0(d_tmp[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[4]), .B1(d_tmp[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15606), .COUT(n15607), .S0(d6_71__N_1459[3]), 
          .S1(d6_71__N_1459[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_4 (.A0(d_d_tmp[1]), .B0(d_tmp[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[2]), .B1(d_tmp[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15605), .COUT(n15606), .S0(d6_71__N_1459[1]), 
          .S1(d6_71__N_1459[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_30 (.A0(d_d7[27]), .B0(d7[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[28]), .B1(d7[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16126), .COUT(n16127), .S0(d8_71__N_1603[27]), .S1(d8_71__N_1603[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_11 (.A0(d4[44]), .B0(cout_adj_2810), .C0(n159_adj_5312), 
          .D0(d5[44]), .A1(d4[45]), .B1(cout_adj_2810), .C1(n156_adj_5311), 
          .D1(d5[45]), .CIN(n16048), .COUT(n16049), .S0(d5_71__N_706[44]), 
          .S1(d5_71__N_706[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[0]), .B1(d_tmp[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15605), .S1(d6_71__N_1459[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1601_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1601_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15604), .S0(cout_adj_4835));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1380_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1380_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16134));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1460_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1460_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_36 (.A0(d2_adj_5711[34]), .B0(d1_adj_5710[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[35]), .B1(d1_adj_5710[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15603), .COUT(n15604), .S0(d2_71__N_490_adj_5727[34]), 
          .S1(d2_71__N_490_adj_5727[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_28 (.A0(d_d7[25]), .B0(d7[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[26]), .B1(d7[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16125), .COUT(n16126), .S0(d8_71__N_1603[25]), .S1(d8_71__N_1603[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_9 (.A0(d2[42]), .B0(cout), .C0(n165_adj_5183), 
          .D0(d3[42]), .A1(d2[43]), .B1(cout), .C1(n162_adj_5182), .D1(d3[43]), 
          .CIN(n16137), .COUT(n16138), .S0(d3_71__N_562[42]), .S1(d3_71__N_562[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_34 (.A0(d2_adj_5711[32]), .B0(d1_adj_5710[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[33]), .B1(d1_adj_5710[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15602), .COUT(n15603), .S0(d2_71__N_490_adj_5727[32]), 
          .S1(d2_71__N_490_adj_5727[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_38 (.A0(d_d7[35]), .B0(d7[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16130), .S0(d8_71__N_1603[35]), .S1(cout_adj_5575));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1490_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_38.INJECT1_1 = "NO";
    FD1S3AX ISquare_e3__i1 (.D(n126_adj_5248), .CK(CIC1_out_clkSin), .Q(ISquare[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i1.GSR = "ENABLED";
    CCU2C _add_1_1380_add_4_32 (.A0(d2_adj_5711[30]), .B0(d1_adj_5710[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[31]), .B1(d1_adj_5710[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15601), .COUT(n15602), .S0(d2_71__N_490_adj_5727[30]), 
          .S1(d2_71__N_490_adj_5727[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_4 (.A0(d2_adj_5711[37]), .B0(d1_adj_5710[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[38]), .B1(d1_adj_5710[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16023), .COUT(n16024), .S0(n180_adj_5642), 
          .S1(n177_adj_5641));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_26 (.A0(d_d7[23]), .B0(d7[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[24]), .B1(d7[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16124), .COUT(n16125), .S0(d8_71__N_1603[23]), .S1(d8_71__N_1603[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_26.INJECT1_1 = "NO";
    PFUMX i2652 (.BLUT(n11972), .ALUT(n12249), .C0(n17389), .Z(n12557));
    CCU2C _add_1_1460_add_4_15 (.A0(d2[48]), .B0(cout), .C0(n147_adj_5177), 
          .D0(d3[48]), .A1(d2[49]), .B1(cout), .C1(n144_adj_5176), .D1(d3[49]), 
          .CIN(n16140), .COUT(n16141), .S0(d3_71__N_562[48]), .S1(d3_71__N_562[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_19 (.A0(d3[52]), .B0(cout_adj_4267), .C0(n135_adj_5268), 
          .D0(d4[52]), .A1(d3[53]), .B1(cout_adj_4267), .C1(n132_adj_5267), 
          .D1(d4[53]), .CIN(n16074), .COUT(n16075), .S0(d4_71__N_634[52]), 
          .S1(d4_71__N_634[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_36 (.A0(d_d7[33]), .B0(d7[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[34]), .B1(d7[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16129), .COUT(n16130), .S0(d8_71__N_1603[33]), .S1(d8_71__N_1603[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_7 (.A0(d2[40]), .B0(cout), .C0(n171_adj_5185), 
          .D0(d3[40]), .A1(d2[41]), .B1(cout), .C1(n168_adj_5184), .D1(d3[41]), 
          .CIN(n16136), .COUT(n16137), .S0(d3_71__N_562[40]), .S1(d3_71__N_562[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_34 (.A0(d_d7[31]), .B0(d7[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[32]), .B1(d7[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16128), .COUT(n16129), .S0(d8_71__N_1603[31]), .S1(d8_71__N_1603[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_24 (.A0(d_d7[21]), .B0(d7[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[22]), .B1(d7[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16123), .COUT(n16124), .S0(d8_71__N_1603[21]), .S1(d8_71__N_1603[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1460_add_4_5 (.A0(d2[38]), .B0(cout), .C0(n177_adj_5187), 
          .D0(d3[38]), .A1(d2[39]), .B1(cout), .C1(n174_adj_5186), .D1(d3[39]), 
          .CIN(n16135), .COUT(n16136), .S0(d3_71__N_562[38]), .S1(d3_71__N_562[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1460_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1460_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1460_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1460_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_22 (.A0(d_d7[19]), .B0(d7[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[20]), .B1(d7[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16122), .COUT(n16123), .S0(d8_71__N_1603[19]), .S1(d8_71__N_1603[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_9 (.A0(d4[42]), .B0(cout_adj_2810), .C0(n165_adj_5314), 
          .D0(d5[42]), .A1(d4[43]), .B1(cout_adj_2810), .C1(n162_adj_5313), 
          .D1(d5[43]), .CIN(n16047), .COUT(n16048), .S0(d5_71__N_706[42]), 
          .S1(d5_71__N_706[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_17 (.A0(d3[50]), .B0(cout_adj_4267), .C0(n141_adj_5270), 
          .D0(d4[50]), .A1(d3[51]), .B1(cout_adj_4267), .C1(n138_adj_5269), 
          .D1(d4[51]), .CIN(n16073), .COUT(n16074), .S0(d4_71__N_634[50]), 
          .S1(d4_71__N_634[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_20 (.A0(d_d7[17]), .B0(d7[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[18]), .B1(d7[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16121), .COUT(n16122), .S0(d8_71__N_1603[17]), .S1(d8_71__N_1603[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_18 (.A0(d_d7[15]), .B0(d7[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[16]), .B1(d7[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16120), .COUT(n16121), .S0(d8_71__N_1603[15]), .S1(d8_71__N_1603[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_30 (.A0(d2_adj_5711[28]), .B0(d1_adj_5710[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[29]), .B1(d1_adj_5710[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15600), .COUT(n15601), .S0(d2_71__N_490_adj_5727[28]), 
          .S1(d2_71__N_490_adj_5727[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_30.INJECT1_1 = "NO";
    PFUMX i2642 (.BLUT(n11966), .ALUT(n12247), .C0(n17389), .Z(n12547));
    CCU2C _add_1_1380_add_4_28 (.A0(d2_adj_5711[26]), .B0(d1_adj_5710[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[27]), .B1(d1_adj_5710[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15599), .COUT(n15600), .S0(d2_71__N_490_adj_5727[26]), 
          .S1(d2_71__N_490_adj_5727[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_26 (.A0(d2_adj_5711[24]), .B0(d1_adj_5710[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[25]), .B1(d1_adj_5710[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15598), .COUT(n15599), .S0(d2_71__N_490_adj_5727[24]), 
          .S1(d2_71__N_490_adj_5727[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_26.INJECT1_1 = "NO";
    OB led_pad_7 (.I(led_c_7), .O(led[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(44[22:25])
    CCU2C _add_1_1490_add_4_10 (.A0(d_d7[7]), .B0(d7[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[8]), .B1(d7[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16116), .COUT(n16117), .S0(d8_71__N_1603[7]), .S1(d8_71__N_1603[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_24 (.A0(d2_adj_5711[22]), .B0(d1_adj_5710[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[23]), .B1(d1_adj_5710[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15597), .COUT(n15598), .S0(d2_71__N_490_adj_5727[22]), 
          .S1(d2_71__N_490_adj_5727[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_5 (.A0(d4[38]), .B0(cout_adj_2810), .C0(n177_adj_5318), 
          .D0(d5[38]), .A1(d4[39]), .B1(cout_adj_2810), .C1(n174_adj_5317), 
          .D1(d5[39]), .CIN(n16045), .COUT(n16046), .S0(d5_71__N_706[38]), 
          .S1(d5_71__N_706[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_9 (.A0(d6_adj_5715[42]), .B0(cout_adj_5464), 
          .C0(n165_adj_4907), .D0(n31_adj_4746), .A1(d6_adj_5715[43]), 
          .B1(cout_adj_5464), .C1(n162_adj_4906), .D1(n30_adj_4747), .CIN(n16177), 
          .COUT(n16178), .S0(d7_71__N_1531_adj_5743[42]), .S1(d7_71__N_1531_adj_5743[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_7 (.A0(d6_adj_5715[40]), .B0(cout_adj_5464), 
          .C0(n171_adj_4909), .D0(n33_adj_4733), .A1(d6_adj_5715[41]), 
          .B1(cout_adj_5464), .C1(n168_adj_4908), .D1(n32_adj_4745), .CIN(n16176), 
          .COUT(n16177), .S0(d7_71__N_1531_adj_5743[40]), .S1(d7_71__N_1531_adj_5743[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d2_adj_5711[36]), .B1(d1_adj_5710[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16023), .S1(n183_adj_5643));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1544_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_38 (.A0(d_d6[35]), .B0(d6[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16022), .S0(d7_71__N_1531[35]), .S1(cout_adj_5644));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1493_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_16 (.A0(d_d7[13]), .B0(d7[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[14]), .B1(d7[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16119), .COUT(n16120), .S0(d8_71__N_1603[13]), .S1(d8_71__N_1603[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_14 (.A0(d_d7[11]), .B0(d7[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[12]), .B1(d7[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16118), .COUT(n16119), .S0(d8_71__N_1603[11]), .S1(d8_71__N_1603[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1490_add_4_12 (.A0(d_d7[9]), .B0(d7[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[10]), .B1(d7[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16117), .COUT(n16118), .S0(d8_71__N_1603[9]), .S1(d8_71__N_1603[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1490_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1490_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1490_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1490_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_22 (.A0(d2_adj_5711[20]), .B0(d1_adj_5710[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[21]), .B1(d1_adj_5710[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15596), .COUT(n15597), .S0(d2_71__N_490_adj_5727[20]), 
          .S1(d2_71__N_490_adj_5727[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_5 (.A0(d6_adj_5715[38]), .B0(cout_adj_5464), 
          .C0(n177_adj_4911), .D0(n35_adj_4735), .A1(d6_adj_5715[39]), 
          .B1(cout_adj_5464), .C1(n174_adj_4910), .D1(n34_adj_4734), .CIN(n16175), 
          .COUT(n16176), .S0(d7_71__N_1531_adj_5743[38]), .S1(d7_71__N_1531_adj_5743[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_5.INJECT1_1 = "NO";
    LUT4 mux_305_i42_4_lut_4_lut (.A(n17822), .B(n12538), .C(n8_adj_4739), 
         .D(n200), .Z(n1953)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam mux_305_i42_4_lut_4_lut.init = 16'h5410;
    LUT4 mux_305_i2_4_lut (.A(n320), .B(n11959), .C(n17815), .D(n17809), 
         .Z(n1993)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i2_4_lut.init = 16'h0aca;
    LUT4 i2065_3_lut (.A(led_c_0), .B(n316), .C(led_c_4), .Z(n11959)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2065_3_lut.init = 16'hcaca;
    CCU2C _add_1_1493_add_4_36 (.A0(d_d6[33]), .B0(d6[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[34]), .B1(d6[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16021), .COUT(n16022), .S0(d7_71__N_1531[33]), .S1(d7_71__N_1531[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_15 (.A0(d3[48]), .B0(cout_adj_4267), .C0(n147_adj_5272), 
          .D0(d4[48]), .A1(d3[49]), .B1(cout_adj_4267), .C1(n144_adj_5271), 
          .D1(d4[49]), .CIN(n16072), .COUT(n16073), .S0(d4_71__N_634[48]), 
          .S1(d4_71__N_634[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_15.INJECT1_1 = "NO";
    OB led_pad_5 (.I(led_c_5), .O(led[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(44[22:25])
    CCU2C _add_1_1418_add_4_3 (.A0(d6_adj_5715[36]), .B0(cout_adj_5464), 
          .C0(n183_adj_4913), .D0(n37_adj_4737), .A1(d6_adj_5715[37]), 
          .B1(cout_adj_5464), .C1(n180_adj_4912), .D1(n36_adj_4736), .CIN(n16174), 
          .COUT(n16175), .S0(d7_71__N_1531_adj_5743[36]), .S1(d7_71__N_1531_adj_5743[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_3.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n12538), .B(n18096), .C(n16837), .D(n17081), .Z(clk_80mhz_enable_1388)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C))) */ ;
    defparam i1_4_lut.init = 16'hcc8c;
    CCU2C _add_1_1457_add_4_13 (.A0(d3[46]), .B0(cout_adj_4267), .C0(n153_adj_5274), 
          .D0(d4[46]), .A1(d3[47]), .B1(cout_adj_4267), .C1(n150_adj_5273), 
          .D1(d4[47]), .CIN(n16071), .COUT(n16072), .S0(d4_71__N_634[46]), 
          .S1(d4_71__N_634[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_13.INJECT1_1 = "NO";
    CCU2C add_3663_5 (.A0(n80), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1878[17]), .B1(d_out_d_11__N_1880[17]), .C1(n77), 
          .D1(VCC_net), .CIN(n16338), .COUT(n16339), .S0(n87_adj_5204), 
          .S1(n84_adj_5203));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3663_5.INIT0 = 16'haaa0;
    defparam add_3663_5.INIT1 = 16'h9696;
    defparam add_3663_5.INJECT1_0 = "NO";
    defparam add_3663_5.INJECT1_1 = "NO";
    LUT4 i3263_4_lut (.A(n314), .B(n17822), .C(n12245), .D(n12538), 
         .Z(n12542)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i3263_4_lut.init = 16'h2230;
    CCU2C add_3663_3 (.A0(d_out_d_11__N_1880[17]), .B0(ISquare[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[13]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16337), .COUT(n16338), .S1(n90_adj_5205));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3663_3.INIT0 = 16'h666a;
    defparam add_3663_3.INIT1 = 16'h555f;
    defparam add_3663_3.INJECT1_0 = "NO";
    defparam add_3663_3.INJECT1_1 = "NO";
    OB o_Tx_Serial_pad (.I(GND_net), .O(o_Tx_Serial));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(43[22:33])
    LUT4 i1280_1_lut (.A(led_c_2), .Z(n3674)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1280_1_lut.init = 16'h5555;
    CCU2C add_3663_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1880[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16337));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3663_1.INIT0 = 16'h0000;
    defparam add_3663_1.INIT1 = 16'haaaf;
    defparam add_3663_1.INJECT1_0 = "NO";
    defparam add_3663_1.INJECT1_1 = "NO";
    LUT4 i2342_3_lut (.A(n12701), .B(n310), .C(led_c_4), .Z(n12245)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2342_3_lut.init = 16'hc5c5;
    FD1P3IX phase_inc_carrGen_i0_i16 (.D(n12559), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i16.GSR = "ENABLED";
    CCU2C _add_1_1493_add_4_34 (.A0(d_d6[31]), .B0(d6[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[32]), .B1(d6[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16020), .COUT(n16021), .S0(d7_71__N_1531[31]), .S1(d7_71__N_1531[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_32 (.A0(d_d6[29]), .B0(d6[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[30]), .B1(d6[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16019), .COUT(n16020), .S0(d7_71__N_1531[29]), .S1(d7_71__N_1531[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_32.INJECT1_1 = "NO";
    LUT4 mux_305_i22_4_lut_4_lut (.A(n17822), .B(n12538), .C(n8_adj_5699), 
         .D(n260), .Z(n1973)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam mux_305_i22_4_lut_4_lut.init = 16'h5410;
    CCU2C _add_1_1380_add_4_20 (.A0(d2_adj_5711[18]), .B0(d1_adj_5710[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[19]), .B1(d1_adj_5710[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15595), .COUT(n15596), .S0(d2_71__N_490_adj_5727[18]), 
          .S1(d2_71__N_490_adj_5727[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_18 (.A0(d2_adj_5711[16]), .B0(d1_adj_5710[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[17]), .B1(d1_adj_5710[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15594), .COUT(n15595), .S0(d2_71__N_490_adj_5727[16]), 
          .S1(d2_71__N_490_adj_5727[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_16 (.A0(d2_adj_5711[14]), .B0(d1_adj_5710[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[15]), .B1(d1_adj_5710[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15593), .COUT(n15594), .S0(d2_71__N_490_adj_5727[14]), 
          .S1(d2_71__N_490_adj_5727[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_14 (.A0(d2_adj_5711[12]), .B0(d1_adj_5710[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[13]), .B1(d1_adj_5710[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15592), .COUT(n15593), .S0(d2_71__N_490_adj_5727[12]), 
          .S1(d2_71__N_490_adj_5727[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_14.INJECT1_1 = "NO";
    LUT4 mux_745_i3_3_lut_4_lut (.A(n12424), .B(n17825), .C(led_c_4), 
         .D(led_c_2), .Z(n3728)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam mux_745_i3_3_lut_4_lut.init = 16'hf780;
    FD1S3AX o_Rx_Byte_i8 (.D(o_Rx_Byte1[7]), .CK(clk_80mhz), .Q(led_c_7));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam o_Rx_Byte_i8.GSR = "ENABLED";
    LUT4 i365_2_lut_rep_200 (.A(n18096), .B(n16837), .Z(n17822)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i365_2_lut_rep_200.init = 16'h2222;
    FD1S3AX o_Rx_Byte_i7 (.D(o_Rx_Byte1[6]), .CK(clk_80mhz), .Q(led_c_6));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    LUT4 i5986_4_lut_4_lut (.A(n18096), .B(n16837), .C(n17069), .D(n17813), 
         .Z(clk_80mhz_enable_1408)) /* synthesis lut_function=(A (((D)+!C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i5986_4_lut_4_lut.init = 16'haa2a;
    FD1S3AX o_Rx_Byte_i6 (.D(o_Rx_Byte1[5]), .CK(clk_80mhz), .Q(led_c_5));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i5 (.D(o_Rx_Byte1[4]), .CK(clk_80mhz), .Q(led_c_4));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    CCU2C _add_1_1493_add_4_30 (.A0(d_d6[27]), .B0(d6[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[28]), .B1(d6[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16018), .COUT(n16019), .S0(d7_71__N_1531[27]), .S1(d7_71__N_1531[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_30.INJECT1_1 = "NO";
    FD1S3AX _add_1_1565_i7 (.D(cout_adj_5576), .CK(clk_80mhz), .Q(PWMOutP4_c));
    defparam _add_1_1565_i7.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i4 (.D(o_Rx_Byte1[3]), .CK(clk_80mhz), .Q(led_c_3));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i3 (.D(o_Rx_Byte1[2]), .CK(clk_80mhz), .Q(led_c_2));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i2 (.D(o_Rx_Byte1[1]), .CK(clk_80mhz), .Q(led_c_1));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    CCU2C _add_1_1493_add_4_28 (.A0(d_d6[25]), .B0(d6[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[26]), .B1(d6[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16017), .COUT(n16018), .S0(d7_71__N_1531[25]), .S1(d7_71__N_1531[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_26 (.A0(d_d6[23]), .B0(d6[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[24]), .B1(d6[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16016), .COUT(n16017), .S0(d7_71__N_1531[23]), .S1(d7_71__N_1531[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_26.INJECT1_1 = "NO";
    LUT4 i4_2_lut_rep_193_3_lut (.A(n18096), .B(n16837), .C(n12538), .Z(n17815)) /* synthesis lut_function=(!(A (B (C))+!A (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i4_2_lut_rep_193_3_lut.init = 16'h2f2f;
    CCU2C _add_1_1493_add_4_24 (.A0(d_d6[21]), .B0(d6[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[22]), .B1(d6[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16015), .COUT(n16016), .S0(d7_71__N_1531[21]), .S1(d7_71__N_1531[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_22 (.A0(d_d6[19]), .B0(d6[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[20]), .B1(d6[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16014), .COUT(n16015), .S0(d7_71__N_1531[19]), .S1(d7_71__N_1531[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_22.INJECT1_1 = "NO";
    LUT4 i2354_3_lut (.A(n12256), .B(n203), .C(n12538), .Z(n12257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2354_3_lut.init = 16'hcaca;
    CCU2C _add_1_1493_add_4_20 (.A0(d_d6[17]), .B0(d6[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[18]), .B1(d6[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16013), .COUT(n16014), .S0(d7_71__N_1531[17]), .S1(d7_71__N_1531[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_18 (.A0(d_d6[15]), .B0(d6[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[16]), .B1(d6[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16012), .COUT(n16013), .S0(d7_71__N_1531[15]), .S1(d7_71__N_1531[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_16 (.A0(d_d6[13]), .B0(d6[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[14]), .B1(d6[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16011), .COUT(n16012), .S0(d7_71__N_1531[13]), .S1(d7_71__N_1531[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_14 (.A0(d_d6[11]), .B0(d6[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[12]), .B1(d6[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16010), .COUT(n16011), .S0(d7_71__N_1531[11]), .S1(d7_71__N_1531[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_12 (.A0(d_d6[9]), .B0(d6[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[10]), .B1(d6[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16009), .COUT(n16010), .S0(d7_71__N_1531[9]), .S1(d7_71__N_1531[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_10 (.A0(d_d6[7]), .B0(d6[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[8]), .B1(d6[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16008), .COUT(n16009), .S0(d7_71__N_1531[7]), .S1(d7_71__N_1531[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_10.INJECT1_1 = "NO";
    LUT4 i5068_2_lut (.A(MultResult2[0]), .B(MultResult1[0]), .Z(n126_adj_5248)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5068_2_lut.init = 16'h6666;
    CCU2C _add_1_1493_add_4_8 (.A0(d_d6[5]), .B0(d6[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[6]), .B1(d6[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16007), .COUT(n16008), .S0(d7_71__N_1531[5]), .S1(d7_71__N_1531[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1493_add_4_6 (.A0(d_d6[3]), .B0(d6[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[4]), .B1(d6[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16006), .COUT(n16007), .S0(d7_71__N_1531[3]), .S1(d7_71__N_1531[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_6.INJECT1_1 = "NO";
    LUT4 i5512_3_lut_rep_192_4_lut (.A(n17825), .B(led_c_3), .C(n17834), 
         .D(n16869), .Z(n17814)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i5512_3_lut_rep_192_4_lut.init = 16'h2220;
    LUT4 mux_305_i6_4_lut (.A(n308), .B(n11963), .C(n17815), .D(n17809), 
         .Z(n1989)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i6_4_lut.init = 16'h0aca;
    LUT4 i2069_3_lut (.A(n11962), .B(n304), .C(n18053), .Z(n11963)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2069_3_lut.init = 16'hcaca;
    LUT4 mux_305_i20_4_lut_4_lut (.A(n17822), .B(n12538), .C(n8_adj_5698), 
         .D(n266), .Z(n1975)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam mux_305_i20_4_lut_4_lut.init = 16'h5410;
    CCU2C _add_1_1493_add_4_4 (.A0(d_d6[1]), .B0(d6[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[2]), .B1(d6[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16005), .COUT(n16006), .S0(d7_71__N_1531[1]), .S1(d7_71__N_1531[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1493_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_4.INJECT1_1 = "NO";
    LUT4 i2356_3_lut (.A(n12258), .B(n179), .C(n12538), .Z(n12259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2356_3_lut.init = 16'hcaca;
    CCU2C _add_1_1493_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[0]), .B1(d6[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16005), .S1(d7_71__N_1531[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1493_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1493_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1493_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1493_add_4_2.INJECT1_1 = "NO";
    CCU2C add_3664_19 (.A0(d_out_d_11__N_1890[17]), .B0(n48_adj_5446), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1890[17]), .B1(n45_adj_5445), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16331), .S0(n916), .S1(d_out_d_11__N_1892[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3664_19.INIT0 = 16'h9995;
    defparam add_3664_19.INIT1 = 16'h9995;
    defparam add_3664_19.INJECT1_0 = "NO";
    defparam add_3664_19.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_38 (.A0(d_d7[71]), .B0(d7[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16004), .S0(n78_adj_5645));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1562_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_38.INJECT1_1 = "NO";
    LUT4 i2358_3_lut (.A(n12260), .B(n164), .C(n12538), .Z(n12261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2358_3_lut.init = 16'hcaca;
    CCU2C _add_1_1457_add_4_11 (.A0(d3[44]), .B0(cout_adj_4267), .C0(n159_adj_5276), 
          .D0(d4[44]), .A1(d3[45]), .B1(cout_adj_4267), .C1(n156_adj_5275), 
          .D1(d4[45]), .CIN(n16070), .COUT(n16071), .S0(d4_71__N_634[44]), 
          .S1(d4_71__N_634[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_38 (.A0(d5_adj_5714[71]), .B0(d4_adj_5713[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16170), .S0(n78_adj_5538));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1553_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_34 (.A0(d5_adj_5714[67]), .B0(d4_adj_5713[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[68]), .B1(d4_adj_5713[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16168), .COUT(n16169), .S0(n90_adj_5542), 
          .S1(n87_adj_5541));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_9 (.A0(d3[42]), .B0(cout_adj_4267), .C0(n165_adj_5278), 
          .D0(d4[42]), .A1(d3[43]), .B1(cout_adj_4267), .C1(n162_adj_5277), 
          .D1(d4[43]), .CIN(n16069), .COUT(n16070), .S0(d4_71__N_634[42]), 
          .S1(d4_71__N_634[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_32 (.A0(d5_adj_5714[65]), .B0(d4_adj_5713[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[66]), .B1(d4_adj_5713[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16167), .COUT(n16168), .S0(n96_adj_5544), 
          .S1(n93_adj_5543));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_36 (.A0(d_d7[69]), .B0(d7[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[70]), .B1(d7[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16003), .COUT(n16004), .S0(n84_adj_5647), .S1(n81_adj_5646));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_34 (.A0(d_d7[67]), .B0(d7[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[68]), .B1(d7[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16002), .COUT(n16003), .S0(n90_adj_5649), .S1(n87_adj_5648));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_32 (.A0(d_d7[65]), .B0(d7[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[66]), .B1(d7[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16001), .COUT(n16002), .S0(n96_adj_5651), .S1(n93_adj_5650));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_32.INJECT1_1 = "NO";
    SinCos SinCos_inst (.clk_80mhz(clk_80mhz), .VCC_net(VCC_net), .GND_net(GND_net), 
           .\phase_accum[57] (phase_accum[57]), .\phase_accum[58] (phase_accum[58]), 
           .\phase_accum[59] (phase_accum[59]), .\phase_accum[60] (phase_accum[60]), 
           .\phase_accum[61] (phase_accum[61]), .\phase_accum[62] (phase_accum[62]), 
           .\phase_accum[63] (phase_accum[63]), .\LOSine[1] (LOSine[1]), 
           .\LOSine[2] (LOSine[2]), .\LOSine[3] (LOSine[3]), .\LOSine[4] (LOSine[4]), 
           .\LOSine[5] (LOSine[5]), .\LOSine[6] (LOSine[6]), .\LOSine[7] (LOSine[7]), 
           .\LOSine[8] (LOSine[8]), .\LOSine[9] (LOSine[9]), .\LOSine[10] (LOSine[10]), 
           .\LOSine[11] (LOSine[11]), .\LOSine[12] (LOSine[12]), .\LOCosine[1] (LOCosine[1]), 
           .\LOCosine[2] (LOCosine[2]), .\LOCosine[3] (LOCosine[3]), .\LOCosine[4] (LOCosine[4]), 
           .\LOCosine[5] (LOCosine[5]), .\LOCosine[6] (LOCosine[6]), .\LOCosine[7] (LOCosine[7]), 
           .\LOCosine[8] (LOCosine[8]), .\LOCosine[9] (LOCosine[9]), .\LOCosine[10] (LOCosine[10]), 
           .\LOCosine[11] (LOCosine[11]), .\LOCosine[12] (LOCosine[12]), 
           .\phase_accum[56] (phase_accum[56])) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    CCU2C _add_1_1562_add_4_30 (.A0(d_d7[63]), .B0(d7[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[64]), .B1(d7[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16000), .COUT(n16001), .S0(n102_adj_5653), .S1(n99_adj_5652));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_30.INJECT1_1 = "NO";
    LUT4 PWMOut_I_0_1_lut (.A(PWMOutP4_c), .Z(PWMOutN4_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(92[22:29])
    defparam PWMOut_I_0_1_lut.init = 16'h5555;
    CCU2C _add_1_1562_add_4_28 (.A0(d_d7[61]), .B0(d7[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[62]), .B1(d7[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15999), .COUT(n16000), .S0(n108_adj_5655), .S1(n105_adj_5654));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_26 (.A0(d_d7[59]), .B0(d7[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[60]), .B1(d7[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15998), .COUT(n15999), .S0(n114_adj_5657), .S1(n111_adj_5656));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_26.INJECT1_1 = "NO";
    LUT4 i354_2_lut_rep_191_3_lut_4_lut (.A(n17825), .B(led_c_3), .C(led_c_4), 
         .D(n17834), .Z(n17813)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i354_2_lut_rep_191_3_lut_4_lut.init = 16'h0200;
    CCU2C _add_1_1562_add_4_24 (.A0(d_d7[57]), .B0(d7[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[58]), .B1(d7[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15997), .COUT(n15998), .S0(n120_adj_5659), .S1(n117_adj_5658));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_7 (.A0(d3[40]), .B0(cout_adj_4267), .C0(n171_adj_5280), 
          .D0(d4[40]), .A1(d3[41]), .B1(cout_adj_4267), .C1(n168_adj_5279), 
          .D1(d4[41]), .CIN(n16068), .COUT(n16069), .S0(d4_71__N_634[40]), 
          .S1(d4_71__N_634[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_5 (.A0(d3[38]), .B0(cout_adj_4267), .C0(n177_adj_5282), 
          .D0(d4[38]), .A1(d3[39]), .B1(cout_adj_4267), .C1(n174_adj_5281), 
          .D1(d4[39]), .CIN(n16067), .COUT(n16068), .S0(d4_71__N_634[38]), 
          .S1(d4_71__N_634[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1457_add_4_3 (.A0(d3[36]), .B0(cout_adj_4267), .C0(n183_adj_5284), 
          .D0(d4[36]), .A1(d3[37]), .B1(cout_adj_4267), .C1(n180_adj_5283), 
          .D1(d4[37]), .CIN(n16066), .COUT(n16067), .S0(d4_71__N_634[36]), 
          .S1(d4_71__N_634[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1457_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1457_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_3.INJECT1_1 = "NO";
    LUT4 mux_305_i8_4_lut (.A(n302), .B(n11965), .C(n17815), .D(n17809), 
         .Z(n1987)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i8_4_lut.init = 16'h0aca;
    CCU2C _add_1_1457_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_4267), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16066));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1457_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1457_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1457_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1457_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_37 (.A0(d4[70]), .B0(cout_adj_2810), .C0(n81_adj_5286), 
          .D0(d5[70]), .A1(d4[71]), .B1(cout_adj_2810), .C1(n78_adj_5285), 
          .D1(d5[71]), .CIN(n16061), .S0(d5_71__N_706[70]), .S1(d5_71__N_706[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_35 (.A0(d4[68]), .B0(cout_adj_2810), .C0(n87_adj_5288), 
          .D0(d5[68]), .A1(d4[69]), .B1(cout_adj_2810), .C1(n84_adj_5287), 
          .D1(d5[69]), .CIN(n16060), .COUT(n16061), .S0(d5_71__N_706[68]), 
          .S1(d5_71__N_706[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_33 (.A0(d4[66]), .B0(cout_adj_2810), .C0(n93_adj_5290), 
          .D0(d5[66]), .A1(d4[67]), .B1(cout_adj_2810), .C1(n90_adj_5289), 
          .D1(d5[67]), .CIN(n16059), .COUT(n16060), .S0(d5_71__N_706[66]), 
          .S1(d5_71__N_706[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_31 (.A0(d4[64]), .B0(cout_adj_2810), .C0(n99_adj_5292), 
          .D0(d5[64]), .A1(d4[65]), .B1(cout_adj_2810), .C1(n96_adj_5291), 
          .D1(d5[65]), .CIN(n16058), .COUT(n16059), .S0(d5_71__N_706[64]), 
          .S1(d5_71__N_706[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_31.INJECT1_1 = "NO";
    LUT4 i364_2_lut_rep_190_3_lut_4_lut (.A(n17825), .B(led_c_3), .C(n18053), 
         .D(n16869), .Z(n17812)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i364_2_lut_rep_190_3_lut_4_lut.init = 16'h0200;
    CCU2C _add_1_1562_add_4_22 (.A0(d_d7[55]), .B0(d7[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[56]), .B1(d7[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15996), .COUT(n15997), .S0(n126_adj_5661), .S1(n123_adj_5660));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_20 (.A0(d_d7[53]), .B0(d7[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[54]), .B1(d7[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15995), .COUT(n15996), .S0(n132_adj_5663), .S1(n129_adj_5662));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_18 (.A0(d_d7[51]), .B0(d7[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[52]), .B1(d7[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15994), .COUT(n15995), .S0(n138_adj_5665), .S1(n135_adj_5664));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_16 (.A0(d_d7[49]), .B0(d7[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[50]), .B1(d7[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15993), .COUT(n15994), .S0(n144_adj_5667), .S1(n141_adj_5666));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_14 (.A0(d_d7[47]), .B0(d7[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[48]), .B1(d7[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15992), .COUT(n15993), .S0(n150_adj_5669), .S1(n147_adj_5668));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_12 (.A0(d_d7[45]), .B0(d7[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[46]), .B1(d7[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15991), .COUT(n15992), .S0(n156_adj_5671), .S1(n153_adj_5670));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_10 (.A0(d_d7[43]), .B0(d7[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[44]), .B1(d7[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15990), .COUT(n15991), .S0(n162_adj_5673), .S1(n159_adj_5672));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_8 (.A0(d_d7[41]), .B0(d7[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[42]), .B1(d7[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15989), .COUT(n15990), .S0(n168_adj_5675), .S1(n165_adj_5674));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_6 (.A0(d_d7[39]), .B0(d7[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[40]), .B1(d7[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15988), .COUT(n15989), .S0(n174_adj_5677), .S1(n171_adj_5676));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_4 (.A0(d_d7[37]), .B0(d7[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[38]), .B1(d7[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15987), .COUT(n15988), .S0(n180_adj_5679), .S1(n177_adj_5678));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1562_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1562_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[36]), .B1(d7[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15987), .S1(n183_adj_5680));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1562_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1562_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1562_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1562_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_37 (.A0(d7_adj_5717[70]), .B0(cout_adj_5501), 
          .C0(n81_adj_4915), .D0(n3_adj_4764), .A1(d7_adj_5717[71]), .B1(cout_adj_5501), 
          .C1(n78_adj_4914), .D1(n2_adj_4763), .CIN(n15985), .S0(d8_71__N_1603_adj_5744[70]), 
          .S1(d8_71__N_1603_adj_5744[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_35 (.A0(d7_adj_5717[68]), .B0(cout_adj_5501), 
          .C0(n87_adj_4917), .D0(n5_adj_4766), .A1(d7_adj_5717[69]), .B1(cout_adj_5501), 
          .C1(n84_adj_4916), .D1(n4_adj_4765), .CIN(n15984), .COUT(n15985), 
          .S0(d8_71__N_1603_adj_5744[68]), .S1(d8_71__N_1603_adj_5744[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_33 (.A0(d7_adj_5717[66]), .B0(cout_adj_5501), 
          .C0(n93_adj_4919), .D0(n7_adj_4768), .A1(d7_adj_5717[67]), .B1(cout_adj_5501), 
          .C1(n90_adj_4918), .D1(n6_adj_4767), .CIN(n15983), .COUT(n15984), 
          .S0(d8_71__N_1603_adj_5744[66]), .S1(d8_71__N_1603_adj_5744[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_31 (.A0(d7_adj_5717[64]), .B0(cout_adj_5501), 
          .C0(n99_adj_4921), .D0(n9_adj_4770), .A1(d7_adj_5717[65]), .B1(cout_adj_5501), 
          .C1(n96_adj_4920), .D1(n8_adj_4769), .CIN(n15982), .COUT(n15983), 
          .S0(d8_71__N_1603_adj_5744[64]), .S1(d8_71__N_1603_adj_5744[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_29 (.A0(d7_adj_5717[62]), .B0(cout_adj_5501), 
          .C0(n105_adj_4923), .D0(n11_adj_4772), .A1(d7_adj_5717[63]), 
          .B1(cout_adj_5501), .C1(n102_adj_4922), .D1(n10_adj_4771), .CIN(n15981), 
          .COUT(n15982), .S0(d8_71__N_1603_adj_5744[62]), .S1(d8_71__N_1603_adj_5744[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_27 (.A0(d7_adj_5717[60]), .B0(cout_adj_5501), 
          .C0(n111_adj_4925), .D0(n13_adj_4774), .A1(d7_adj_5717[61]), 
          .B1(cout_adj_5501), .C1(n108_adj_4924), .D1(n12_adj_4773), .CIN(n15980), 
          .COUT(n15981), .S0(d8_71__N_1603_adj_5744[60]), .S1(d8_71__N_1603_adj_5744[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_25 (.A0(d7_adj_5717[58]), .B0(cout_adj_5501), 
          .C0(n117_adj_4927), .D0(n15_adj_4776), .A1(d7_adj_5717[59]), 
          .B1(cout_adj_5501), .C1(n114_adj_4926), .D1(n14_adj_4775), .CIN(n15979), 
          .COUT(n15980), .S0(d8_71__N_1603_adj_5744[58]), .S1(d8_71__N_1603_adj_5744[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_23 (.A0(d7_adj_5717[56]), .B0(cout_adj_5501), 
          .C0(n123_adj_4929), .D0(n17_adj_4778), .A1(d7_adj_5717[57]), 
          .B1(cout_adj_5501), .C1(n120_adj_4928), .D1(n16_adj_4777), .CIN(n15978), 
          .COUT(n15979), .S0(d8_71__N_1603_adj_5744[56]), .S1(d8_71__N_1603_adj_5744[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_21 (.A0(d7_adj_5717[54]), .B0(cout_adj_5501), 
          .C0(n129_adj_4931), .D0(n19_adj_4780), .A1(d7_adj_5717[55]), 
          .B1(cout_adj_5501), .C1(n126_adj_4930), .D1(n18_adj_4779), .CIN(n15977), 
          .COUT(n15978), .S0(d8_71__N_1603_adj_5744[54]), .S1(d8_71__N_1603_adj_5744[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_19 (.A0(d7_adj_5717[52]), .B0(cout_adj_5501), 
          .C0(n135_adj_4933), .D0(n21_adj_4782), .A1(d7_adj_5717[53]), 
          .B1(cout_adj_5501), .C1(n132_adj_4932), .D1(n20_adj_4781), .CIN(n15976), 
          .COUT(n15977), .S0(d8_71__N_1603_adj_5744[52]), .S1(d8_71__N_1603_adj_5744[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_17 (.A0(d7_adj_5717[50]), .B0(cout_adj_5501), 
          .C0(n141_adj_4935), .D0(n23_adj_4784), .A1(d7_adj_5717[51]), 
          .B1(cout_adj_5501), .C1(n138_adj_4934), .D1(n22_adj_4783), .CIN(n15975), 
          .COUT(n15976), .S0(d8_71__N_1603_adj_5744[50]), .S1(d8_71__N_1603_adj_5744[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_15 (.A0(d7_adj_5717[48]), .B0(cout_adj_5501), 
          .C0(n147_adj_4937), .D0(n25_adj_4786), .A1(d7_adj_5717[49]), 
          .B1(cout_adj_5501), .C1(n144_adj_4936), .D1(n24_adj_4785), .CIN(n15974), 
          .COUT(n15975), .S0(d8_71__N_1603_adj_5744[48]), .S1(d8_71__N_1603_adj_5744[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_13 (.A0(d7_adj_5717[46]), .B0(cout_adj_5501), 
          .C0(n153_adj_4939), .D0(n27_adj_4788), .A1(d7_adj_5717[47]), 
          .B1(cout_adj_5501), .C1(n150_adj_4938), .D1(n26_adj_4787), .CIN(n15973), 
          .COUT(n15974), .S0(d8_71__N_1603_adj_5744[46]), .S1(d8_71__N_1603_adj_5744[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_11 (.A0(d7_adj_5717[44]), .B0(cout_adj_5501), 
          .C0(n159_adj_4941), .D0(n29_adj_4790), .A1(d7_adj_5717[45]), 
          .B1(cout_adj_5501), .C1(n156_adj_4940), .D1(n28_adj_4789), .CIN(n15972), 
          .COUT(n15973), .S0(d8_71__N_1603_adj_5744[44]), .S1(d8_71__N_1603_adj_5744[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_9 (.A0(d7_adj_5717[42]), .B0(cout_adj_5501), 
          .C0(n165_adj_4943), .D0(n31_adj_4792), .A1(d7_adj_5717[43]), 
          .B1(cout_adj_5501), .C1(n162_adj_4942), .D1(n30_adj_4791), .CIN(n15971), 
          .COUT(n15972), .S0(d8_71__N_1603_adj_5744[42]), .S1(d8_71__N_1603_adj_5744[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_7 (.A0(d7_adj_5717[40]), .B0(cout_adj_5501), 
          .C0(n171_adj_4945), .D0(n33_adj_4794), .A1(d7_adj_5717[41]), 
          .B1(cout_adj_5501), .C1(n168_adj_4944), .D1(n32_adj_4793), .CIN(n15970), 
          .COUT(n15971), .S0(d8_71__N_1603_adj_5744[40]), .S1(d8_71__N_1603_adj_5744[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_5 (.A0(d7_adj_5717[38]), .B0(cout_adj_5501), 
          .C0(n177_adj_4947), .D0(n35_adj_4796), .A1(d7_adj_5717[39]), 
          .B1(cout_adj_5501), .C1(n174_adj_4946), .D1(n34_adj_4795), .CIN(n15969), 
          .COUT(n15970), .S0(d8_71__N_1603_adj_5744[38]), .S1(d8_71__N_1603_adj_5744[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_3 (.A0(d7_adj_5717[36]), .B0(cout_adj_5501), 
          .C0(n183_adj_4949), .D0(n37_adj_4798), .A1(d7_adj_5717[37]), 
          .B1(cout_adj_5501), .C1(n180_adj_4948), .D1(n36_adj_4797), .CIN(n15968), 
          .COUT(n15969), .S0(d8_71__N_1603_adj_5744[36]), .S1(d8_71__N_1603_adj_5744[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1415_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1415_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5501), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15968));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1415_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1415_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1415_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_37 (.A0(d8_adj_5719[70]), .B0(cout_adj_5700), 
          .C0(n81_adj_4951), .D0(n3_adj_4800), .A1(d8_adj_5719[71]), .B1(cout_adj_5700), 
          .C1(n78_adj_4950), .D1(n2_adj_4799), .CIN(n15963), .S0(d9_71__N_1675_adj_5745[70]), 
          .S1(d9_71__N_1675_adj_5745[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_35 (.A0(d8_adj_5719[68]), .B0(cout_adj_5700), 
          .C0(n87_adj_4953), .D0(n5_adj_4802), .A1(d8_adj_5719[69]), .B1(cout_adj_5700), 
          .C1(n84_adj_4952), .D1(n4_adj_4801), .CIN(n15962), .COUT(n15963), 
          .S0(d9_71__N_1675_adj_5745[68]), .S1(d9_71__N_1675_adj_5745[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_33 (.A0(d8_adj_5719[66]), .B0(cout_adj_5700), 
          .C0(n93_adj_4955), .D0(n7_adj_4804), .A1(d8_adj_5719[67]), .B1(cout_adj_5700), 
          .C1(n90_adj_4954), .D1(n6_adj_4803), .CIN(n15961), .COUT(n15962), 
          .S0(d9_71__N_1675_adj_5745[66]), .S1(d9_71__N_1675_adj_5745[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_31 (.A0(d8_adj_5719[64]), .B0(cout_adj_5700), 
          .C0(n99_adj_4957), .D0(n9_adj_4806), .A1(d8_adj_5719[65]), .B1(cout_adj_5700), 
          .C1(n96_adj_4956), .D1(n8_adj_4805), .CIN(n15960), .COUT(n15961), 
          .S0(d9_71__N_1675_adj_5745[64]), .S1(d9_71__N_1675_adj_5745[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_29 (.A0(d8_adj_5719[62]), .B0(cout_adj_5700), 
          .C0(n105_adj_4959), .D0(n11_adj_4808), .A1(d8_adj_5719[63]), 
          .B1(cout_adj_5700), .C1(n102_adj_4958), .D1(n10_adj_4807), .CIN(n15959), 
          .COUT(n15960), .S0(d9_71__N_1675_adj_5745[62]), .S1(d9_71__N_1675_adj_5745[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_27 (.A0(d8_adj_5719[60]), .B0(cout_adj_5700), 
          .C0(n111_adj_4961), .D0(n13_adj_4810), .A1(d8_adj_5719[61]), 
          .B1(cout_adj_5700), .C1(n108_adj_4960), .D1(n12_adj_4809), .CIN(n15958), 
          .COUT(n15959), .S0(d9_71__N_1675_adj_5745[60]), .S1(d9_71__N_1675_adj_5745[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_25 (.A0(d8_adj_5719[58]), .B0(cout_adj_5700), 
          .C0(n117_adj_4963), .D0(n15_adj_4812), .A1(d8_adj_5719[59]), 
          .B1(cout_adj_5700), .C1(n114_adj_4962), .D1(n14_adj_4811), .CIN(n15957), 
          .COUT(n15958), .S0(d9_71__N_1675_adj_5745[58]), .S1(d9_71__N_1675_adj_5745[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_23 (.A0(d8_adj_5719[56]), .B0(cout_adj_5700), 
          .C0(n123_adj_4965), .D0(n17_adj_4814), .A1(d8_adj_5719[57]), 
          .B1(cout_adj_5700), .C1(n120_adj_4964), .D1(n16_adj_4813), .CIN(n15956), 
          .COUT(n15957), .S0(d9_71__N_1675_adj_5745[56]), .S1(d9_71__N_1675_adj_5745[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_21 (.A0(d8_adj_5719[54]), .B0(cout_adj_5700), 
          .C0(n129_adj_4967), .D0(n19_adj_4816), .A1(d8_adj_5719[55]), 
          .B1(cout_adj_5700), .C1(n126_adj_4966), .D1(n18_adj_4815), .CIN(n15955), 
          .COUT(n15956), .S0(d9_71__N_1675_adj_5745[54]), .S1(d9_71__N_1675_adj_5745[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_19 (.A0(d8_adj_5719[52]), .B0(cout_adj_5700), 
          .C0(n135_adj_4969), .D0(n21_adj_4818), .A1(d8_adj_5719[53]), 
          .B1(cout_adj_5700), .C1(n132_adj_4968), .D1(n20_adj_4817), .CIN(n15954), 
          .COUT(n15955), .S0(d9_71__N_1675_adj_5745[52]), .S1(d9_71__N_1675_adj_5745[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_17 (.A0(d8_adj_5719[50]), .B0(cout_adj_5700), 
          .C0(n141_adj_4971), .D0(n23_adj_4820), .A1(d8_adj_5719[51]), 
          .B1(cout_adj_5700), .C1(n138_adj_4970), .D1(n22_adj_4819), .CIN(n15953), 
          .COUT(n15954), .S0(d9_71__N_1675_adj_5745[50]), .S1(d9_71__N_1675_adj_5745[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_15 (.A0(d8_adj_5719[48]), .B0(cout_adj_5700), 
          .C0(n147_adj_4973), .D0(n25_adj_4822), .A1(d8_adj_5719[49]), 
          .B1(cout_adj_5700), .C1(n144_adj_4972), .D1(n24_adj_4821), .CIN(n15952), 
          .COUT(n15953), .S0(d9_71__N_1675_adj_5745[48]), .S1(d9_71__N_1675_adj_5745[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_13 (.A0(d8_adj_5719[46]), .B0(cout_adj_5700), 
          .C0(n153_adj_4975), .D0(n27_adj_4824), .A1(d8_adj_5719[47]), 
          .B1(cout_adj_5700), .C1(n150_adj_4974), .D1(n26_adj_4823), .CIN(n15951), 
          .COUT(n15952), .S0(d9_71__N_1675_adj_5745[46]), .S1(d9_71__N_1675_adj_5745[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_11 (.A0(d8_adj_5719[44]), .B0(cout_adj_5700), 
          .C0(n159_adj_4977), .D0(n29_adj_4826), .A1(d8_adj_5719[45]), 
          .B1(cout_adj_5700), .C1(n156_adj_4976), .D1(n28_adj_4825), .CIN(n15950), 
          .COUT(n15951), .S0(d9_71__N_1675_adj_5745[44]), .S1(d9_71__N_1675_adj_5745[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_9 (.A0(d8_adj_5719[42]), .B0(cout_adj_5700), 
          .C0(n165_adj_4979), .D0(n31_adj_4828), .A1(d8_adj_5719[43]), 
          .B1(cout_adj_5700), .C1(n162_adj_4978), .D1(n30_adj_4827), .CIN(n15949), 
          .COUT(n15950), .S0(d9_71__N_1675_adj_5745[42]), .S1(d9_71__N_1675_adj_5745[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_7 (.A0(d8_adj_5719[40]), .B0(cout_adj_5700), 
          .C0(n171_adj_4981), .D0(n33_adj_4830), .A1(d8_adj_5719[41]), 
          .B1(cout_adj_5700), .C1(n168_adj_4980), .D1(n32_adj_4829), .CIN(n15948), 
          .COUT(n15949), .S0(d9_71__N_1675_adj_5745[40]), .S1(d9_71__N_1675_adj_5745[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_5 (.A0(d8_adj_5719[38]), .B0(cout_adj_5700), 
          .C0(n177_adj_4983), .D0(n35_adj_4832), .A1(d8_adj_5719[39]), 
          .B1(cout_adj_5700), .C1(n174_adj_4982), .D1(n34_adj_4831), .CIN(n15947), 
          .COUT(n15948), .S0(d9_71__N_1675_adj_5745[38]), .S1(d9_71__N_1675_adj_5745[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_3 (.A0(d8_adj_5719[36]), .B0(cout_adj_5700), 
          .C0(n183_adj_4985), .D0(n37_adj_4834), .A1(d8_adj_5719[37]), 
          .B1(cout_adj_5700), .C1(n180_adj_4984), .D1(n36_adj_4833), .CIN(n15946), 
          .COUT(n15947), .S0(d9_71__N_1675_adj_5745[36]), .S1(d9_71__N_1675_adj_5745[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1412_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1412_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5700), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15946));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1412_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1412_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1412_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_37 (.A0(d_tmp_adj_5708[70]), .B0(cout_adj_5463), 
          .C0(n81_adj_4843), .D0(n3), .A1(d_tmp_adj_5708[71]), .B1(cout_adj_5463), 
          .C1(n78_adj_4842), .D1(n2), .CIN(n15941), .S0(d6_71__N_1459_adj_5742[70]), 
          .S1(d6_71__N_1459_adj_5742[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_35 (.A0(d_tmp_adj_5708[68]), .B0(cout_adj_5463), 
          .C0(n87_adj_4845), .D0(n5), .A1(d_tmp_adj_5708[69]), .B1(cout_adj_5463), 
          .C1(n84_adj_4844), .D1(n4), .CIN(n15940), .COUT(n15941), .S0(d6_71__N_1459_adj_5742[68]), 
          .S1(d6_71__N_1459_adj_5742[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_33 (.A0(d_tmp_adj_5708[66]), .B0(cout_adj_5463), 
          .C0(n93_adj_4847), .D0(n7), .A1(d_tmp_adj_5708[67]), .B1(cout_adj_5463), 
          .C1(n90_adj_4846), .D1(n6), .CIN(n15939), .COUT(n15940), .S0(d6_71__N_1459_adj_5742[66]), 
          .S1(d6_71__N_1459_adj_5742[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_31 (.A0(d_tmp_adj_5708[64]), .B0(cout_adj_5463), 
          .C0(n99_adj_4849), .D0(n9), .A1(d_tmp_adj_5708[65]), .B1(cout_adj_5463), 
          .C1(n96_adj_4848), .D1(n8), .CIN(n15938), .COUT(n15939), .S0(d6_71__N_1459_adj_5742[64]), 
          .S1(d6_71__N_1459_adj_5742[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_29 (.A0(d_tmp_adj_5708[62]), .B0(cout_adj_5463), 
          .C0(n105_adj_4851), .D0(n11), .A1(d_tmp_adj_5708[63]), .B1(cout_adj_5463), 
          .C1(n102_adj_4850), .D1(n10), .CIN(n15937), .COUT(n15938), 
          .S0(d6_71__N_1459_adj_5742[62]), .S1(d6_71__N_1459_adj_5742[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_27 (.A0(d_tmp_adj_5708[60]), .B0(cout_adj_5463), 
          .C0(n111_adj_4853), .D0(n13), .A1(d_tmp_adj_5708[61]), .B1(cout_adj_5463), 
          .C1(n108_adj_4852), .D1(n12), .CIN(n15936), .COUT(n15937), 
          .S0(d6_71__N_1459_adj_5742[60]), .S1(d6_71__N_1459_adj_5742[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_25 (.A0(d_tmp_adj_5708[58]), .B0(cout_adj_5463), 
          .C0(n117_adj_4855), .D0(n15), .A1(d_tmp_adj_5708[59]), .B1(cout_adj_5463), 
          .C1(n114_adj_4854), .D1(n14), .CIN(n15935), .COUT(n15936), 
          .S0(d6_71__N_1459_adj_5742[58]), .S1(d6_71__N_1459_adj_5742[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_23 (.A0(d_tmp_adj_5708[56]), .B0(cout_adj_5463), 
          .C0(n123_adj_4857), .D0(n17), .A1(d_tmp_adj_5708[57]), .B1(cout_adj_5463), 
          .C1(n120_adj_4856), .D1(n16), .CIN(n15934), .COUT(n15935), 
          .S0(d6_71__N_1459_adj_5742[56]), .S1(d6_71__N_1459_adj_5742[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_21 (.A0(d_tmp_adj_5708[54]), .B0(cout_adj_5463), 
          .C0(n129_adj_4859), .D0(n19), .A1(d_tmp_adj_5708[55]), .B1(cout_adj_5463), 
          .C1(n126_adj_4858), .D1(n18), .CIN(n15933), .COUT(n15934), 
          .S0(d6_71__N_1459_adj_5742[54]), .S1(d6_71__N_1459_adj_5742[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_19 (.A0(d_tmp_adj_5708[52]), .B0(cout_adj_5463), 
          .C0(n135_adj_4861), .D0(n21), .A1(d_tmp_adj_5708[53]), .B1(cout_adj_5463), 
          .C1(n132_adj_4860), .D1(n20), .CIN(n15932), .COUT(n15933), 
          .S0(d6_71__N_1459_adj_5742[52]), .S1(d6_71__N_1459_adj_5742[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_17 (.A0(d_tmp_adj_5708[50]), .B0(cout_adj_5463), 
          .C0(n141_adj_4863), .D0(n23), .A1(d_tmp_adj_5708[51]), .B1(cout_adj_5463), 
          .C1(n138_adj_4862), .D1(n22), .CIN(n15931), .COUT(n15932), 
          .S0(d6_71__N_1459_adj_5742[50]), .S1(d6_71__N_1459_adj_5742[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_15 (.A0(d_tmp_adj_5708[48]), .B0(cout_adj_5463), 
          .C0(n147_adj_4865), .D0(n25), .A1(d_tmp_adj_5708[49]), .B1(cout_adj_5463), 
          .C1(n144_adj_4864), .D1(n24), .CIN(n15930), .COUT(n15931), 
          .S0(d6_71__N_1459_adj_5742[48]), .S1(d6_71__N_1459_adj_5742[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_13 (.A0(d_tmp_adj_5708[46]), .B0(cout_adj_5463), 
          .C0(n153_adj_4867), .D0(n27), .A1(d_tmp_adj_5708[47]), .B1(cout_adj_5463), 
          .C1(n150_adj_4866), .D1(n26), .CIN(n15929), .COUT(n15930), 
          .S0(d6_71__N_1459_adj_5742[46]), .S1(d6_71__N_1459_adj_5742[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_11 (.A0(d_tmp_adj_5708[44]), .B0(cout_adj_5463), 
          .C0(n159_adj_4869), .D0(n29), .A1(d_tmp_adj_5708[45]), .B1(cout_adj_5463), 
          .C1(n156_adj_4868), .D1(n28), .CIN(n15928), .COUT(n15929), 
          .S0(d6_71__N_1459_adj_5742[44]), .S1(d6_71__N_1459_adj_5742[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_9 (.A0(d_tmp_adj_5708[42]), .B0(cout_adj_5463), 
          .C0(n165_adj_4871), .D0(n31), .A1(d_tmp_adj_5708[43]), .B1(cout_adj_5463), 
          .C1(n162_adj_4870), .D1(n30), .CIN(n15927), .COUT(n15928), 
          .S0(d6_71__N_1459_adj_5742[42]), .S1(d6_71__N_1459_adj_5742[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_7 (.A0(d_tmp_adj_5708[40]), .B0(cout_adj_5463), 
          .C0(n171_adj_4873), .D0(n33), .A1(d_tmp_adj_5708[41]), .B1(cout_adj_5463), 
          .C1(n168_adj_4872), .D1(n32), .CIN(n15926), .COUT(n15927), 
          .S0(d6_71__N_1459_adj_5742[40]), .S1(d6_71__N_1459_adj_5742[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_5 (.A0(d_tmp_adj_5708[38]), .B0(cout_adj_5463), 
          .C0(n177_adj_4875), .D0(n35), .A1(d_tmp_adj_5708[39]), .B1(cout_adj_5463), 
          .C1(n174_adj_4874), .D1(n34), .CIN(n15925), .COUT(n15926), 
          .S0(d6_71__N_1459_adj_5742[38]), .S1(d6_71__N_1459_adj_5742[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_5.INJECT1_1 = "NO";
    CCU2C add_3664_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1890[17]), .C0(n54_adj_5448), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1890[17]), 
          .C1(n51_adj_5447), .D1(VCC_net), .CIN(n16330), .COUT(n16331), 
          .S0(n918), .S1(n917));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3664_17.INIT0 = 16'h6969;
    defparam add_3664_17.INIT1 = 16'h6969;
    defparam add_3664_17.INJECT1_0 = "NO";
    defparam add_3664_17.INJECT1_1 = "NO";
    CCU2C add_3664_15 (.A0(d_out_d_11__N_1890[17]), .B0(n60_adj_5450), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1890[17]), 
          .C1(n57_adj_5449), .D1(VCC_net), .CIN(n16329), .COUT(n16330), 
          .S0(n920), .S1(n919));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3664_15.INIT0 = 16'h9995;
    defparam add_3664_15.INIT1 = 16'h6969;
    defparam add_3664_15.INJECT1_0 = "NO";
    defparam add_3664_15.INJECT1_1 = "NO";
    CCU2C add_3664_13 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n66_adj_5452), .D0(VCC_net), .A1(d_out_d_11__N_1890[17]), 
          .B1(n17826), .C1(n63_adj_5451), .D1(VCC_net), .CIN(n16328), 
          .COUT(n16329), .S0(n922), .S1(n921));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3664_13.INIT0 = 16'h9696;
    defparam add_3664_13.INIT1 = 16'h6969;
    defparam add_3664_13.INJECT1_0 = "NO";
    defparam add_3664_13.INJECT1_1 = "NO";
    CCU2C add_3664_11 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n72_adj_5454), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(n69_adj_5453), .D1(VCC_net), 
          .CIN(n16327), .COUT(n16328), .S0(n924), .S1(n923));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3664_11.INIT0 = 16'h9696;
    defparam add_3664_11.INIT1 = 16'h9696;
    defparam add_3664_11.INJECT1_0 = "NO";
    defparam add_3664_11.INJECT1_1 = "NO";
    CCU2C add_3664_9 (.A0(d_out_d_11__N_1882[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n78_adj_5456), .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(n75_adj_5455), .D1(VCC_net), 
          .CIN(n16326), .COUT(n16327), .S0(n926), .S1(n925));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3664_9.INIT0 = 16'h9696;
    defparam add_3664_9.INIT1 = 16'h9696;
    defparam add_3664_9.INJECT1_0 = "NO";
    defparam add_3664_9.INJECT1_1 = "NO";
    CCU2C add_3664_7 (.A0(d_out_d_11__N_1886[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n84_adj_5458), .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(n81_adj_5457), .D1(VCC_net), 
          .CIN(n16325), .COUT(n16326), .S0(n928), .S1(n927));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3664_7.INIT0 = 16'h9696;
    defparam add_3664_7.INIT1 = 16'h9696;
    defparam add_3664_7.INJECT1_0 = "NO";
    defparam add_3664_7.INJECT1_1 = "NO";
    CCU2C add_3664_5 (.A0(n90_adj_5460), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1888[17]), .B1(d_out_d_11__N_1890[17]), .C1(n87_adj_5459), 
          .D1(VCC_net), .CIN(n16324), .COUT(n16325), .S0(n930), .S1(n929));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3664_5.INIT0 = 16'haaa0;
    defparam add_3664_5.INIT1 = 16'h9696;
    defparam add_3664_5.INJECT1_0 = "NO";
    defparam add_3664_5.INJECT1_1 = "NO";
    CCU2C add_3664_3 (.A0(d_out_d_11__N_1890[17]), .B0(ISquare[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16323), .COUT(n16324), .S1(n931));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3664_3.INIT0 = 16'h666a;
    defparam add_3664_3.INIT1 = 16'h555f;
    defparam add_3664_3.INJECT1_0 = "NO";
    defparam add_3664_3.INJECT1_1 = "NO";
    CCU2C add_3664_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1890[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16323));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3664_1.INIT0 = 16'h0000;
    defparam add_3664_1.INIT1 = 16'haaaf;
    defparam add_3664_1.INJECT1_0 = "NO";
    defparam add_3664_1.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_38 (.A0(d_d9[35]), .B0(d9[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16318), .S1(cout_adj_5462));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1484_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_36 (.A0(d_d9[33]), .B0(d9[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[34]), .B1(d9[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16317), .COUT(n16318));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_34 (.A0(d_d9[31]), .B0(d9[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[32]), .B1(d9[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16316), .COUT(n16317));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_32 (.A0(d_d9[29]), .B0(d9[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[30]), .B1(d9[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16315), .COUT(n16316));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_32.INJECT1_1 = "NO";
    FD1S3AX phase_accum_e3_i0_i1 (.D(n318), .CK(clk_80mhz), .Q(phase_accum_adj_5702[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i1.GSR = "ENABLED";
    CCU2C _add_1_1484_add_4_30 (.A0(d_d9[27]), .B0(d9[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[28]), .B1(d9[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16314), .COUT(n16315));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_30.INJECT1_1 = "NO";
    LUT4 i2071_3_lut (.A(n11964), .B(n298), .C(n18053), .Z(n11965)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2071_3_lut.init = 16'hcaca;
    CCU2C _add_1_1484_add_4_28 (.A0(d_d9[25]), .B0(d9[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[26]), .B1(d9[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16313), .COUT(n16314));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_26 (.A0(d_d9[23]), .B0(d9[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[24]), .B1(d9[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16312), .COUT(n16313));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_24 (.A0(d_d9[21]), .B0(d9[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[22]), .B1(d9[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16311), .COUT(n16312));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_22 (.A0(d_d9[19]), .B0(d9[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[20]), .B1(d9[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16310), .COUT(n16311));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_22.INJECT1_1 = "NO";
    LUT4 i5871_2_lut_rep_188_3_lut_4_lut (.A(n17825), .B(led_c_3), .C(n18053), 
         .D(n16869), .Z(n17810)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i5871_2_lut_rep_188_3_lut_4_lut.init = 16'hf2f0;
    CCU2C _add_1_1484_add_4_20 (.A0(d_d9[17]), .B0(d9[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[18]), .B1(d9[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16309), .COUT(n16310));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_18 (.A0(d_d9[15]), .B0(d9[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[16]), .B1(d9[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16308), .COUT(n16309));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_16 (.A0(d_d9[13]), .B0(d9[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[14]), .B1(d9[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16307), .COUT(n16308));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_16.INJECT1_1 = "NO";
    LUT4 mux_305_i12_4_lut_4_lut (.A(n17822), .B(n12538), .C(n8_adj_5574), 
         .D(n290), .Z(n1983)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam mux_305_i12_4_lut_4_lut.init = 16'h5410;
    CCU2C _add_1_1484_add_4_14 (.A0(d_d9[11]), .B0(d9[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[12]), .B1(d9[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16306), .COUT(n16307));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_12 (.A0(d_d9[9]), .B0(d9[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[10]), .B1(d9[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16305), .COUT(n16306));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_12.INJECT1_1 = "NO";
    LUT4 i19_4_lut (.A(n280_adj_5074), .B(n286), .C(n18053), .D(n17814), 
         .Z(n8_adj_5574)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i19_4_lut.init = 16'hc0ca;
    LUT4 mux_305_i16_4_lut (.A(n278), .B(n11975), .C(n17815), .D(n17809), 
         .Z(n1979)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i16_4_lut.init = 16'h0aca;
    CCU2C _add_1_1484_add_4_10 (.A0(d_d9[7]), .B0(d9[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[8]), .B1(d9[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16304), .COUT(n16305));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_8 (.A0(d_d9[5]), .B0(d9[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[6]), .B1(d9[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16303), .COUT(n16304));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1484_add_4_6 (.A0(d_d9[3]), .B0(d9[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[4]), .B1(d9[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16302), .COUT(n16303));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_6.INJECT1_1 = "NO";
    LUT4 i2081_3_lut (.A(n11974), .B(n274), .C(n18053), .Z(n11975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2081_3_lut.init = 16'hcaca;
    CCU2C _add_1_1484_add_4_4 (.A0(d_d9[1]), .B0(d9[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[2]), .B1(d9[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16301), .COUT(n16302));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1484_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_4.INJECT1_1 = "NO";
    LUT4 i1989_2_lut_rep_187_3_lut_4_lut (.A(n17823), .B(n17834), .C(n17822), 
         .D(led_c_4), .Z(n17809)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i1989_2_lut_rep_187_3_lut_4_lut.init = 16'hf0f8;
    CCU2C _add_1_1484_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[0]), .B1(d9[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16301));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1484_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1484_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1484_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1484_add_4_2.INJECT1_1 = "NO";
    LUT4 i19_4_lut_adj_68 (.A(n256_adj_5066), .B(n262), .C(led_c_4), .D(n17814), 
         .Z(n8_adj_5698)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i19_4_lut_adj_68.init = 16'hc0ca;
    CCU2C _add_1_1550_add_4_38 (.A0(d4_adj_5713[71]), .B0(d3_adj_5712[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16300), .S0(n78_adj_5409));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1550_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_38.INJECT1_1 = "NO";
    LUT4 i5947_3_lut_4_lut (.A(n17823), .B(n17834), .C(led_c_4), .D(n12538), 
         .Z(n17389)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i5947_3_lut_4_lut.init = 16'hfff8;
    LUT4 i19_4_lut_adj_69 (.A(n250_adj_5064), .B(n256), .C(n18053), .D(n17814), 
         .Z(n8_adj_5699)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i19_4_lut_adj_69.init = 16'hc0ca;
    CCU2C _add_1_1550_add_4_36 (.A0(d4_adj_5713[69]), .B0(d3_adj_5712[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[70]), .B1(d3_adj_5712[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16299), .COUT(n16300), .S0(n84_adj_5411), 
          .S1(n81_adj_5410));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_34 (.A0(d4_adj_5713[67]), .B0(d3_adj_5712[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[68]), .B1(d3_adj_5712[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16298), .COUT(n16299), .S0(n90_adj_5413), 
          .S1(n87_adj_5412));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_34.INJECT1_1 = "NO";
    LUT4 mux_305_i25_4_lut (.A(n251), .B(n2621), .C(n17815), .D(n17809), 
         .Z(n1970)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i25_4_lut.init = 16'h0aca;
    CCU2C _add_1_1550_add_4_32 (.A0(d4_adj_5713[65]), .B0(d3_adj_5712[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[66]), .B1(d3_adj_5712[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16297), .COUT(n16298), .S0(n96_adj_5415), 
          .S1(n93_adj_5414));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_30 (.A0(d4_adj_5713[63]), .B0(d3_adj_5712[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[64]), .B1(d3_adj_5712[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16296), .COUT(n16297), .S0(n102_adj_5417), 
          .S1(n99_adj_5416));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_30.INJECT1_1 = "NO";
    LUT4 mux_305_i27_4_lut (.A(n245), .B(n11983), .C(n17815), .D(n17809), 
         .Z(n1968)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i27_4_lut.init = 16'h0aca;
    CCU2C _add_1_1550_add_4_28 (.A0(d4_adj_5713[61]), .B0(d3_adj_5712[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[62]), .B1(d3_adj_5712[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16295), .COUT(n16296), .S0(n108_adj_5419), 
          .S1(n105_adj_5418));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_26 (.A0(d4_adj_5713[59]), .B0(d3_adj_5712[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[60]), .B1(d3_adj_5712[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16294), .COUT(n16295), .S0(n114_adj_5421), 
          .S1(n111_adj_5420));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_26.INJECT1_1 = "NO";
    LUT4 i2089_3_lut (.A(n11982), .B(n241), .C(led_c_4), .Z(n11983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2089_3_lut.init = 16'hcaca;
    CCU2C _add_1_1550_add_4_24 (.A0(d4_adj_5713[57]), .B0(d3_adj_5712[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[58]), .B1(d3_adj_5712[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16293), .COUT(n16294), .S0(n120_adj_5423), 
          .S1(n117_adj_5422));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_22 (.A0(d4_adj_5713[55]), .B0(d3_adj_5712[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[56]), .B1(d3_adj_5712[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16292), .COUT(n16293), .S0(n126_adj_5425), 
          .S1(n123_adj_5424));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_22.INJECT1_1 = "NO";
    LUT4 mux_305_i31_4_lut (.A(n233), .B(n11987), .C(n17815), .D(n17809), 
         .Z(n1964)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i31_4_lut.init = 16'h0aca;
    LUT4 i2093_3_lut (.A(n11986), .B(n229), .C(led_c_4), .Z(n11987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2093_3_lut.init = 16'hcaca;
    CCU2C _add_1_1550_add_4_20 (.A0(d4_adj_5713[53]), .B0(d3_adj_5712[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[54]), .B1(d3_adj_5712[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16291), .COUT(n16292), .S0(n132_adj_5427), 
          .S1(n129_adj_5426));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_20.INJECT1_1 = "NO";
    FD1S3AX phase_accum_e3_i0_i2 (.D(n315), .CK(clk_80mhz), .Q(phase_accum_adj_5702[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i2.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i3 (.D(n312), .CK(clk_80mhz), .Q(phase_accum_adj_5702[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i3.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i4 (.D(n309), .CK(clk_80mhz), .Q(phase_accum_adj_5702[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i4.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i5 (.D(n306), .CK(clk_80mhz), .Q(phase_accum_adj_5702[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i5.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i6 (.D(n303), .CK(clk_80mhz), .Q(phase_accum_adj_5702[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i6.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i7 (.D(n300), .CK(clk_80mhz), .Q(phase_accum_adj_5702[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i7.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i8 (.D(n297), .CK(clk_80mhz), .Q(phase_accum_adj_5702[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i8.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i9 (.D(n294), .CK(clk_80mhz), .Q(phase_accum_adj_5702[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i9.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i10 (.D(n291), .CK(clk_80mhz), .Q(phase_accum_adj_5702[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i10.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i11 (.D(n288), .CK(clk_80mhz), .Q(phase_accum_adj_5702[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i11.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i12 (.D(n285), .CK(clk_80mhz), .Q(phase_accum_adj_5702[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i12.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i13 (.D(n282), .CK(clk_80mhz), .Q(phase_accum_adj_5702[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i13.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i14 (.D(n279), .CK(clk_80mhz), .Q(phase_accum_adj_5702[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i14.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i15 (.D(n276), .CK(clk_80mhz), .Q(phase_accum_adj_5702[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i15.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i16 (.D(n273), .CK(clk_80mhz), .Q(phase_accum_adj_5702[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i16.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i17 (.D(n270), .CK(clk_80mhz), .Q(phase_accum_adj_5702[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i17.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i18 (.D(n267), .CK(clk_80mhz), .Q(phase_accum_adj_5702[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i18.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i19 (.D(n264), .CK(clk_80mhz), .Q(phase_accum_adj_5702[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i19.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i20 (.D(n261), .CK(clk_80mhz), .Q(phase_accum_adj_5702[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i20.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i21 (.D(n258), .CK(clk_80mhz), .Q(phase_accum_adj_5702[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i21.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i22 (.D(n255), .CK(clk_80mhz), .Q(phase_accum_adj_5702[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i22.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i23 (.D(n252), .CK(clk_80mhz), .Q(phase_accum_adj_5702[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i23.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i24 (.D(n249), .CK(clk_80mhz), .Q(phase_accum_adj_5702[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i24.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i25 (.D(n246), .CK(clk_80mhz), .Q(phase_accum_adj_5702[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i25.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i26 (.D(n243), .CK(clk_80mhz), .Q(phase_accum_adj_5702[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i26.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i27 (.D(n240), .CK(clk_80mhz), .Q(phase_accum_adj_5702[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i27.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i28 (.D(n237), .CK(clk_80mhz), .Q(phase_accum_adj_5702[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i28.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i29 (.D(n234), .CK(clk_80mhz), .Q(phase_accum_adj_5702[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i29.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i30 (.D(n231), .CK(clk_80mhz), .Q(phase_accum_adj_5702[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i30.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i31 (.D(n228), .CK(clk_80mhz), .Q(phase_accum_adj_5702[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i31.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i32 (.D(n225), .CK(clk_80mhz), .Q(phase_accum_adj_5702[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i32.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i33 (.D(n222), .CK(clk_80mhz), .Q(phase_accum_adj_5702[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i33.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i34 (.D(n219), .CK(clk_80mhz), .Q(phase_accum_adj_5702[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i34.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i35 (.D(n216), .CK(clk_80mhz), .Q(phase_accum_adj_5702[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i35.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i36 (.D(n213_adj_5020), .CK(clk_80mhz), .Q(phase_accum_adj_5702[36]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i36.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i37 (.D(n210), .CK(clk_80mhz), .Q(phase_accum_adj_5702[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i37.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i38 (.D(n207), .CK(clk_80mhz), .Q(phase_accum_adj_5702[38]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i38.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i39 (.D(n204), .CK(clk_80mhz), .Q(phase_accum_adj_5702[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i39.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i40 (.D(n201), .CK(clk_80mhz), .Q(phase_accum_adj_5702[40]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i40.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i41 (.D(n198), .CK(clk_80mhz), .Q(phase_accum_adj_5702[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i41.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i42 (.D(n195), .CK(clk_80mhz), .Q(phase_accum_adj_5702[42]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i42.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i43 (.D(n192), .CK(clk_80mhz), .Q(phase_accum_adj_5702[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i43.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i44 (.D(n189), .CK(clk_80mhz), .Q(phase_accum_adj_5702[44]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i44.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i45 (.D(n186), .CK(clk_80mhz), .Q(phase_accum_adj_5702[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i45.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i46 (.D(n183_adj_5019), .CK(clk_80mhz), .Q(phase_accum_adj_5702[46]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i46.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i47 (.D(n180_adj_5018), .CK(clk_80mhz), .Q(phase_accum_adj_5702[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i47.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i48 (.D(n177_adj_5017), .CK(clk_80mhz), .Q(phase_accum_adj_5702[48]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i48.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i49 (.D(n174_adj_5016), .CK(clk_80mhz), .Q(phase_accum_adj_5702[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i49.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i50 (.D(n171_adj_5015), .CK(clk_80mhz), .Q(phase_accum_adj_5702[50]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i50.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i51 (.D(n168_adj_5014), .CK(clk_80mhz), .Q(phase_accum_adj_5702[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i51.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i52 (.D(n165_adj_5013), .CK(clk_80mhz), .Q(phase_accum_adj_5702[52]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i52.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i53 (.D(n162_adj_5012), .CK(clk_80mhz), .Q(phase_accum_adj_5702[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i53.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i54 (.D(n159_adj_5011), .CK(clk_80mhz), .Q(phase_accum_adj_5702[54]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i54.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i55 (.D(n156_adj_5010), .CK(clk_80mhz), .Q(phase_accum_adj_5702[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i55.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i56 (.D(n153_adj_5009), .CK(clk_80mhz), .Q(phase_accum[56]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i56.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i57 (.D(n150_adj_5008), .CK(clk_80mhz), .Q(phase_accum[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i57.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i58 (.D(n147_adj_5007), .CK(clk_80mhz), .Q(phase_accum[58]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i58.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i59 (.D(n144_adj_5006), .CK(clk_80mhz), .Q(phase_accum[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i59.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i60 (.D(n141_adj_5005), .CK(clk_80mhz), .Q(phase_accum[60]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i60.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i61 (.D(n138_adj_5004), .CK(clk_80mhz), .Q(phase_accum[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i61.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i62 (.D(n135_adj_5003), .CK(clk_80mhz), .Q(phase_accum[62]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i62.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i63 (.D(n132_adj_5002), .CK(clk_80mhz), .Q(phase_accum[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i63.GSR = "ENABLED";
    LUT4 mux_305_i33_4_lut (.A(n227), .B(n2613), .C(n17815), .D(n17809), 
         .Z(n1962)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i33_4_lut.init = 16'h0aca;
    CCU2C _add_1_1421_add_4_3 (.A0(d_tmp_adj_5708[36]), .B0(cout_adj_5463), 
          .C0(n183_adj_4877), .D0(n37), .A1(d_tmp_adj_5708[37]), .B1(cout_adj_5463), 
          .C1(n180_adj_4876), .D1(n36), .CIN(n15924), .COUT(n15925), 
          .S0(d6_71__N_1459_adj_5742[36]), .S1(d6_71__N_1459_adj_5742[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1421_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1421_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_3.INJECT1_1 = "NO";
    FD1P3IX phase_inc_carrGen_i0_i39 (.D(n12591), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i39.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i38 (.D(n12589), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[38]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i38.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i37 (.D(n12587), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i37.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i36 (.D(n12585), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[36]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i36.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i35 (.D(n12583), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i35.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i33 (.D(n12581), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i33.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i31 (.D(n12579), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i31.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i29 (.D(n12577), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i29.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i28 (.D(n12575), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i28.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i27 (.D(n12573), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i27.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i25 (.D(n12571), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i25.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i23 (.D(n12569), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i23.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i22 (.D(n12567), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i22.GSR = "ENABLED";
    LUT4 i2345_3_lut (.A(led_c_1), .B(n277), .C(led_c_4), .Z(n12248)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2345_3_lut.init = 16'hc5c5;
    FD1P3IX phase_inc_carrGen_i0_i20 (.D(n12565), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i20.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i18 (.D(n12563), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i18.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i17 (.D(n12561), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i17.GSR = "ENABLED";
    LUT4 i2098_3_lut_4_lut (.A(n17823), .B(n16869), .C(led_c_0), .D(n193_adj_5045), 
         .Z(n11992)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i2098_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_305_i35_4_lut (.A(n221), .B(n11989), .C(n17815), .D(n17809), 
         .Z(n1960)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i35_4_lut.init = 16'h0aca;
    LUT4 i2095_3_lut (.A(n11988), .B(n217), .C(led_c_4), .Z(n11989)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2095_3_lut.init = 16'hcaca;
    FD1P3IX phase_inc_carrGen_i0_i14 (.D(n12557), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i14.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut_4_lut (.A(led_c_0), .B(led_c_3), .C(led_c_1), 
         .D(led_c_2), .Z(n39_adj_4738)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'hf814;
    FD1P3IX phase_inc_carrGen_i0_i13 (.D(n12555), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i13.GSR = "ENABLED";
    CCU2C _add_1_1421_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5463), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15924));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1421_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1421_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1421_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_195_3_lut_4_lut (.A(n18096), .B(n17827), .C(n16869), 
         .D(led_c_3), .Z(n17817)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i1_2_lut_rep_195_3_lut_4_lut.init = 16'h0080;
    FD1P3IX phase_inc_carrGen_i0_i12 (.D(n12553), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i12.GSR = "ENABLED";
    LUT4 i2343_3_lut (.A(led_c_1), .B(n295), .C(led_c_4), .Z(n12246)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2343_3_lut.init = 16'hc5c5;
    CCU2C _add_1_1550_add_4_18 (.A0(d4_adj_5713[51]), .B0(d3_adj_5712[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[52]), .B1(d3_adj_5712[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16290), .COUT(n16291), .S0(n138_adj_5429), 
          .S1(n135_adj_5428));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_16 (.A0(d4_adj_5713[49]), .B0(d3_adj_5712[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[50]), .B1(d3_adj_5712[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16289), .COUT(n16290), .S0(n144_adj_5431), 
          .S1(n141_adj_5430));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_14 (.A0(d4_adj_5713[47]), .B0(d3_adj_5712[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[48]), .B1(d3_adj_5712[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16288), .COUT(n16289), .S0(n150_adj_5433), 
          .S1(n147_adj_5432));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_12 (.A0(d4_adj_5713[45]), .B0(d3_adj_5712[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[46]), .B1(d3_adj_5712[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16287), .COUT(n16288), .S0(n156_adj_5435), 
          .S1(n153_adj_5434));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_10 (.A0(d4_adj_5713[43]), .B0(d3_adj_5712[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[44]), .B1(d3_adj_5712[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16286), .COUT(n16287), .S0(n162_adj_5437), 
          .S1(n159_adj_5436));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_8 (.A0(d4_adj_5713[41]), .B0(d3_adj_5712[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[42]), .B1(d3_adj_5712[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16285), .COUT(n16286), .S0(n168_adj_5439), 
          .S1(n165_adj_5438));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_6 (.A0(d4_adj_5713[39]), .B0(d3_adj_5712[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[40]), .B1(d3_adj_5712[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16284), .COUT(n16285), .S0(n174_adj_5441), 
          .S1(n171_adj_5440));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_4 (.A0(d4_adj_5713[37]), .B0(d3_adj_5712[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[38]), .B1(d3_adj_5712[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16283), .COUT(n16284), .S0(n180_adj_5443), 
          .S1(n177_adj_5442));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1550_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1550_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d4_adj_5713[36]), .B1(d3_adj_5712[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16283), .S1(n183_adj_5444));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1550_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1550_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1550_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1550_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_38 (.A0(d_d_tmp_adj_5709[35]), .B0(d_tmp_adj_5708[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16282), .S0(d6_71__N_1459_adj_5742[35]), 
          .S1(cout_adj_5463));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1481_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_38 (.A0(d_d8_adj_5720[35]), .B0(d8_adj_5719[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15920), .S0(d9_71__N_1675_adj_5745[35]), 
          .S1(cout_adj_5700));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1472_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_36 (.A0(d_d_tmp_adj_5709[33]), .B0(d_tmp_adj_5708[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[34]), .B1(d_tmp_adj_5708[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16281), .COUT(n16282), .S0(d6_71__N_1459_adj_5742[33]), 
          .S1(d6_71__N_1459_adj_5742[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_36.INJECT1_1 = "NO";
    FD1P3IX phase_inc_carrGen_i0_i10 (.D(n12551), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i10.GSR = "ENABLED";
    CCU2C _add_1_1481_add_4_34 (.A0(d_d_tmp_adj_5709[31]), .B0(d_tmp_adj_5708[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[32]), .B1(d_tmp_adj_5708[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16280), .COUT(n16281), .S0(d6_71__N_1459_adj_5742[31]), 
          .S1(d6_71__N_1459_adj_5742[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_32 (.A0(d_d_tmp_adj_5709[29]), .B0(d_tmp_adj_5708[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[30]), .B1(d_tmp_adj_5708[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16279), .COUT(n16280), .S0(d6_71__N_1459_adj_5742[29]), 
          .S1(d6_71__N_1459_adj_5742[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_32.INJECT1_1 = "NO";
    FD1P3IX phase_inc_carrGen_i0_i9 (.D(n12549), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i9.GSR = "ENABLED";
    CCU2C _add_1_1481_add_4_30 (.A0(d_d_tmp_adj_5709[27]), .B0(d_tmp_adj_5708[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[28]), .B1(d_tmp_adj_5708[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16278), .COUT(n16279), .S0(d6_71__N_1459_adj_5742[27]), 
          .S1(d6_71__N_1459_adj_5742[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_36 (.A0(d_d8_adj_5720[33]), .B0(d8_adj_5719[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[34]), .B1(d8_adj_5719[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15919), .COUT(n15920), .S0(d9_71__N_1675_adj_5745[33]), 
          .S1(d9_71__N_1675_adj_5745[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_34 (.A0(d_d8_adj_5720[31]), .B0(d8_adj_5719[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[32]), .B1(d8_adj_5719[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15918), .COUT(n15919), .S0(d9_71__N_1675_adj_5745[31]), 
          .S1(d9_71__N_1675_adj_5745[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_32 (.A0(d_d8_adj_5720[29]), .B0(d8_adj_5719[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[30]), .B1(d8_adj_5719[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15917), .COUT(n15918), .S0(d9_71__N_1675_adj_5745[29]), 
          .S1(d9_71__N_1675_adj_5745[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_32.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_198_3_lut_4_lut (.A(led_c_5), .B(n17835), .C(n12424), 
         .D(n18096), .Z(n17820)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i1_2_lut_rep_198_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_201_3_lut_4_lut (.A(led_c_5), .B(n17835), .C(led_c_3), 
         .D(n18096), .Z(n17823)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i1_2_lut_rep_201_3_lut_4_lut.init = 16'h0800;
    LUT4 i4990_2_lut_rep_206 (.A(ISquare[23]), .B(ISquare[22]), .Z(n17828)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam i4990_2_lut_rep_206.init = 16'heeee;
    CCU2C _add_1_1380_add_4_12 (.A0(d2_adj_5711[10]), .B0(d1_adj_5710[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[11]), .B1(d1_adj_5710[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15591), .COUT(n15592), .S0(d2_71__N_490_adj_5727[10]), 
          .S1(d2_71__N_490_adj_5727[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_10 (.A0(d2_adj_5711[8]), .B0(d1_adj_5710[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[9]), .B1(d1_adj_5710[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15590), .COUT(n15591), .S0(d2_71__N_490_adj_5727[8]), 
          .S1(d2_71__N_490_adj_5727[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_8 (.A0(d2_adj_5711[6]), .B0(d1_adj_5710[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[7]), .B1(d1_adj_5710[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15589), .COUT(n15590), .S0(d2_71__N_490_adj_5727[6]), 
          .S1(d2_71__N_490_adj_5727[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_6 (.A0(d2_adj_5711[4]), .B0(d1_adj_5710[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[5]), .B1(d1_adj_5710[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15588), .COUT(n15589), .S0(d2_71__N_490_adj_5727[4]), 
          .S1(d2_71__N_490_adj_5727[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_4 (.A0(d2_adj_5711[2]), .B0(d1_adj_5710[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[3]), .B1(d1_adj_5710[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15587), .COUT(n15588), .S0(d2_71__N_490_adj_5727[2]), 
          .S1(d2_71__N_490_adj_5727[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1380_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1380_add_4_2 (.A0(d2_adj_5711[0]), .B0(d1_adj_5710[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[1]), .B1(d1_adj_5710[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15587), .S1(d2_71__N_490_adj_5727[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1380_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1380_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1380_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1380_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15585), .S0(cout_adj_4836));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1383_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1383_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_36 (.A0(d3_adj_5712[34]), .B0(d2_adj_5711[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[35]), .B1(d2_adj_5711[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15584), .COUT(n15585), .S0(d3_71__N_562_adj_5728[34]), 
          .S1(d3_71__N_562_adj_5728[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_34 (.A0(d3_adj_5712[32]), .B0(d2_adj_5711[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[33]), .B1(d2_adj_5711[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15583), .COUT(n15584), .S0(d3_71__N_562_adj_5728[32]), 
          .S1(d3_71__N_562_adj_5728[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_32 (.A0(d3_adj_5712[30]), .B0(d2_adj_5711[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[31]), .B1(d2_adj_5711[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15582), .COUT(n15583), .S0(d3_71__N_562_adj_5728[30]), 
          .S1(d3_71__N_562_adj_5728[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_30 (.A0(d3_adj_5712[28]), .B0(d2_adj_5711[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[29]), .B1(d2_adj_5711[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15581), .COUT(n15582), .S0(d3_71__N_562_adj_5728[28]), 
          .S1(d3_71__N_562_adj_5728[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_28 (.A0(d3_adj_5712[26]), .B0(d2_adj_5711[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[27]), .B1(d2_adj_5711[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15580), .COUT(n15581), .S0(d3_71__N_562_adj_5728[26]), 
          .S1(d3_71__N_562_adj_5728[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_26 (.A0(d3_adj_5712[24]), .B0(d2_adj_5711[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[25]), .B1(d2_adj_5711[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15579), .COUT(n15580), .S0(d3_71__N_562_adj_5728[24]), 
          .S1(d3_71__N_562_adj_5728[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_24 (.A0(d3_adj_5712[22]), .B0(d2_adj_5711[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[23]), .B1(d2_adj_5711[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15578), .COUT(n15579), .S0(d3_71__N_562_adj_5728[22]), 
          .S1(d3_71__N_562_adj_5728[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_22 (.A0(d3_adj_5712[20]), .B0(d2_adj_5711[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[21]), .B1(d2_adj_5711[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15577), .COUT(n15578), .S0(d3_71__N_562_adj_5728[20]), 
          .S1(d3_71__N_562_adj_5728[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_20 (.A0(d3_adj_5712[18]), .B0(d2_adj_5711[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[19]), .B1(d2_adj_5711[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15576), .COUT(n15577), .S0(d3_71__N_562_adj_5728[18]), 
          .S1(d3_71__N_562_adj_5728[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_18 (.A0(d3_adj_5712[16]), .B0(d2_adj_5711[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[17]), .B1(d2_adj_5711[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15575), .COUT(n15576), .S0(d3_71__N_562_adj_5728[16]), 
          .S1(d3_71__N_562_adj_5728[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_16 (.A0(d3_adj_5712[14]), .B0(d2_adj_5711[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[15]), .B1(d2_adj_5711[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15574), .COUT(n15575), .S0(d3_71__N_562_adj_5728[14]), 
          .S1(d3_71__N_562_adj_5728[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_14 (.A0(d3_adj_5712[12]), .B0(d2_adj_5711[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[13]), .B1(d2_adj_5711[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15573), .COUT(n15574), .S0(d3_71__N_562_adj_5728[12]), 
          .S1(d3_71__N_562_adj_5728[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_12 (.A0(d3_adj_5712[10]), .B0(d2_adj_5711[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[11]), .B1(d2_adj_5711[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15572), .COUT(n15573), .S0(d3_71__N_562_adj_5728[10]), 
          .S1(d3_71__N_562_adj_5728[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_10 (.A0(d3_adj_5712[8]), .B0(d2_adj_5711[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[9]), .B1(d2_adj_5711[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15571), .COUT(n15572), .S0(d3_71__N_562_adj_5728[8]), 
          .S1(d3_71__N_562_adj_5728[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_8 (.A0(d3_adj_5712[6]), .B0(d2_adj_5711[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[7]), .B1(d2_adj_5711[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15570), .COUT(n15571), .S0(d3_71__N_562_adj_5728[6]), 
          .S1(d3_71__N_562_adj_5728[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_6 (.A0(d3_adj_5712[4]), .B0(d2_adj_5711[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[5]), .B1(d2_adj_5711[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15569), .COUT(n15570), .S0(d3_71__N_562_adj_5728[4]), 
          .S1(d3_71__N_562_adj_5728[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_4 (.A0(d3_adj_5712[2]), .B0(d2_adj_5711[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[3]), .B1(d2_adj_5711[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15568), .COUT(n15569), .S0(d3_71__N_562_adj_5728[2]), 
          .S1(d3_71__N_562_adj_5728[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1383_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1383_add_4_2 (.A0(d3_adj_5712[0]), .B0(d2_adj_5711[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[1]), .B1(d2_adj_5711[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15568), .S1(d3_71__N_562_adj_5728[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1383_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1383_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1383_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1383_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15566), .S0(cout_adj_4558));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1362_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1362_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_36 (.A0(d2[34]), .B0(d1[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[35]), .B1(d1[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15565), .COUT(n15566), .S0(d2_71__N_490[34]), .S1(d2_71__N_490[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_34 (.A0(d2[32]), .B0(d1[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[33]), .B1(d1[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15564), .COUT(n15565), .S0(d2_71__N_490[32]), .S1(d2_71__N_490[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_32 (.A0(d2[30]), .B0(d1[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[31]), .B1(d1[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15563), .COUT(n15564), .S0(d2_71__N_490[30]), .S1(d2_71__N_490[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_30 (.A0(d2[28]), .B0(d1[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[29]), .B1(d1[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15562), .COUT(n15563), .S0(d2_71__N_490[28]), .S1(d2_71__N_490[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_28 (.A0(d2[26]), .B0(d1[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[27]), .B1(d1[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15561), .COUT(n15562), .S0(d2_71__N_490[26]), .S1(d2_71__N_490[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_26 (.A0(d2[24]), .B0(d1[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[25]), .B1(d1[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15560), .COUT(n15561), .S0(d2_71__N_490[24]), .S1(d2_71__N_490[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_24 (.A0(d2[22]), .B0(d1[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[23]), .B1(d1[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15559), .COUT(n15560), .S0(d2_71__N_490[22]), .S1(d2_71__N_490[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_22 (.A0(d2[20]), .B0(d1[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[21]), .B1(d1[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15558), .COUT(n15559), .S0(d2_71__N_490[20]), .S1(d2_71__N_490[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_20 (.A0(d2[18]), .B0(d1[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[19]), .B1(d1[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15557), .COUT(n15558), .S0(d2_71__N_490[18]), .S1(d2_71__N_490[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_18 (.A0(d2[16]), .B0(d1[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[17]), .B1(d1[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15556), .COUT(n15557), .S0(d2_71__N_490[16]), .S1(d2_71__N_490[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_16 (.A0(d2[14]), .B0(d1[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[15]), .B1(d1[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15555), .COUT(n15556), .S0(d2_71__N_490[14]), .S1(d2_71__N_490[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_14 (.A0(d2[12]), .B0(d1[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[13]), .B1(d1[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15554), .COUT(n15555), .S0(d2_71__N_490[12]), .S1(d2_71__N_490[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_12 (.A0(d2[10]), .B0(d1[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[11]), .B1(d1[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15553), .COUT(n15554), .S0(d2_71__N_490[10]), .S1(d2_71__N_490[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_10 (.A0(d2[8]), .B0(d1[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[9]), .B1(d1[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15552), .COUT(n15553), .S0(d2_71__N_490[8]), .S1(d2_71__N_490[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_8 (.A0(d2[6]), .B0(d1[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[7]), .B1(d1[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15551), 
          .COUT(n15552), .S0(d2_71__N_490[6]), .S1(d2_71__N_490[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_6 (.A0(d2[4]), .B0(d1[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[5]), .B1(d1[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15550), 
          .COUT(n15551), .S0(d2_71__N_490[4]), .S1(d2_71__N_490[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_4 (.A0(d2[2]), .B0(d1[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[3]), .B1(d1[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15549), 
          .COUT(n15550), .S0(d2_71__N_490[2]), .S1(d2_71__N_490[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1362_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1362_add_4_2 (.A0(d2[0]), .B0(d1[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[1]), .B1(d1[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15549), 
          .S1(d2_71__N_490[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1362_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1362_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1362_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1362_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15547), .S0(cout));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1365_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1365_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_36 (.A0(d3[34]), .B0(d2[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[35]), .B1(d2[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15546), .COUT(n15547), .S0(d3_71__N_562[34]), .S1(d3_71__N_562[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_34 (.A0(d3[32]), .B0(d2[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[33]), .B1(d2[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15545), .COUT(n15546), .S0(d3_71__N_562[32]), .S1(d3_71__N_562[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_32 (.A0(d3[30]), .B0(d2[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[31]), .B1(d2[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15544), .COUT(n15545), .S0(d3_71__N_562[30]), .S1(d3_71__N_562[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_30 (.A0(d3[28]), .B0(d2[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[29]), .B1(d2[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15543), .COUT(n15544), .S0(d3_71__N_562[28]), .S1(d3_71__N_562[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_28 (.A0(d3[26]), .B0(d2[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[27]), .B1(d2[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15542), .COUT(n15543), .S0(d3_71__N_562[26]), .S1(d3_71__N_562[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_26 (.A0(d3[24]), .B0(d2[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[25]), .B1(d2[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15541), .COUT(n15542), .S0(d3_71__N_562[24]), .S1(d3_71__N_562[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_24 (.A0(d3[22]), .B0(d2[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[23]), .B1(d2[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15540), .COUT(n15541), .S0(d3_71__N_562[22]), .S1(d3_71__N_562[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_22 (.A0(d3[20]), .B0(d2[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[21]), .B1(d2[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15539), .COUT(n15540), .S0(d3_71__N_562[20]), .S1(d3_71__N_562[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_20 (.A0(d3[18]), .B0(d2[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[19]), .B1(d2[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15538), .COUT(n15539), .S0(d3_71__N_562[18]), .S1(d3_71__N_562[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_18 (.A0(d3[16]), .B0(d2[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[17]), .B1(d2[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15537), .COUT(n15538), .S0(d3_71__N_562[16]), .S1(d3_71__N_562[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_16 (.A0(d3[14]), .B0(d2[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[15]), .B1(d2[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15536), .COUT(n15537), .S0(d3_71__N_562[14]), .S1(d3_71__N_562[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_14 (.A0(d3[12]), .B0(d2[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[13]), .B1(d2[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15535), .COUT(n15536), .S0(d3_71__N_562[12]), .S1(d3_71__N_562[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_12 (.A0(d3[10]), .B0(d2[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[11]), .B1(d2[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15534), .COUT(n15535), .S0(d3_71__N_562[10]), .S1(d3_71__N_562[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_10 (.A0(d3[8]), .B0(d2[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[9]), .B1(d2[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15533), .COUT(n15534), .S0(d3_71__N_562[8]), .S1(d3_71__N_562[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_8 (.A0(d3[6]), .B0(d2[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[7]), .B1(d2[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15532), 
          .COUT(n15533), .S0(d3_71__N_562[6]), .S1(d3_71__N_562[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_6 (.A0(d3[4]), .B0(d2[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[5]), .B1(d2[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15531), 
          .COUT(n15532), .S0(d3_71__N_562[4]), .S1(d3_71__N_562[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_4 (.A0(d3[2]), .B0(d2[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[3]), .B1(d2[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15530), 
          .COUT(n15531), .S0(d3_71__N_562[2]), .S1(d3_71__N_562[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1365_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1365_add_4_2 (.A0(d3[0]), .B0(d2[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[1]), .B1(d2[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15530), 
          .S1(d3_71__N_562[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1365_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1365_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1365_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1365_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1403_add_4_13 (.A0(LOSine[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15528), .S0(MixerOutSin_11__N_236[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1403_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_1403_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_1403_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1403_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1403_add_4_11 (.A0(LOSine[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15527), .COUT(n15528), .S0(MixerOutSin_11__N_236[9]), 
          .S1(MixerOutSin_11__N_236[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1403_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_1403_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_1403_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1403_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1403_add_4_9 (.A0(LOSine[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15526), .COUT(n15527), .S0(MixerOutSin_11__N_236[7]), 
          .S1(MixerOutSin_11__N_236[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1403_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_1403_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_1403_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1403_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1403_add_4_7 (.A0(LOSine[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15525), .COUT(n15526), .S0(MixerOutSin_11__N_236[5]), 
          .S1(MixerOutSin_11__N_236[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1403_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_1403_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_1403_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1403_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1403_add_4_5 (.A0(LOSine[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15524), .COUT(n15525), .S0(MixerOutSin_11__N_236[3]), 
          .S1(MixerOutSin_11__N_236[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1403_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_1403_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_1403_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1403_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1403_add_4_3 (.A0(LOSine[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15523), .COUT(n15524), .S0(MixerOutSin_11__N_236[1]), 
          .S1(MixerOutSin_11__N_236[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1403_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_1403_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_1403_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1403_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1403_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15523), .S1(MixerOutSin_11__N_236[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1403_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1403_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_1403_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1403_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_37 (.A0(d_tmp[70]), .B0(cout_adj_5001), .C0(n81_adj_5503), 
          .D0(n3_adj_4724), .A1(d_tmp[71]), .B1(cout_adj_5001), .C1(n78_adj_5502), 
          .D1(n2_adj_4725), .CIN(n15521), .S0(d6_71__N_1459[70]), .S1(d6_71__N_1459[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_35 (.A0(d_tmp[68]), .B0(cout_adj_5001), .C0(n87_adj_5505), 
          .D0(n5_adj_4722), .A1(d_tmp[69]), .B1(cout_adj_5001), .C1(n84_adj_5504), 
          .D1(n4_adj_4723), .CIN(n15520), .COUT(n15521), .S0(d6_71__N_1459[68]), 
          .S1(d6_71__N_1459[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_33 (.A0(d_tmp[66]), .B0(cout_adj_5001), .C0(n93_adj_5507), 
          .D0(n7_adj_4720), .A1(d_tmp[67]), .B1(cout_adj_5001), .C1(n90_adj_5506), 
          .D1(n6_adj_4721), .CIN(n15519), .COUT(n15520), .S0(d6_71__N_1459[66]), 
          .S1(d6_71__N_1459[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_31 (.A0(d_tmp[64]), .B0(cout_adj_5001), .C0(n99_adj_5509), 
          .D0(n9_adj_4718), .A1(d_tmp[65]), .B1(cout_adj_5001), .C1(n96_adj_5508), 
          .D1(n8_adj_4719), .CIN(n15518), .COUT(n15519), .S0(d6_71__N_1459[64]), 
          .S1(d6_71__N_1459[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_29 (.A0(d_tmp[62]), .B0(cout_adj_5001), .C0(n105_adj_5511), 
          .D0(n11_adj_4716), .A1(d_tmp[63]), .B1(cout_adj_5001), .C1(n102_adj_5510), 
          .D1(n10_adj_4717), .CIN(n15517), .COUT(n15518), .S0(d6_71__N_1459[62]), 
          .S1(d6_71__N_1459[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_27 (.A0(d_tmp[60]), .B0(cout_adj_5001), .C0(n111_adj_5513), 
          .D0(n13_adj_4714), .A1(d_tmp[61]), .B1(cout_adj_5001), .C1(n108_adj_5512), 
          .D1(n12_adj_4715), .CIN(n15516), .COUT(n15517), .S0(d6_71__N_1459[60]), 
          .S1(d6_71__N_1459[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_25 (.A0(d_tmp[58]), .B0(cout_adj_5001), .C0(n117_adj_5515), 
          .D0(n15_adj_4712), .A1(d_tmp[59]), .B1(cout_adj_5001), .C1(n114_adj_5514), 
          .D1(n14_adj_4713), .CIN(n15515), .COUT(n15516), .S0(d6_71__N_1459[58]), 
          .S1(d6_71__N_1459[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_23 (.A0(d_tmp[56]), .B0(cout_adj_5001), .C0(n123_adj_5517), 
          .D0(n17_adj_4710), .A1(d_tmp[57]), .B1(cout_adj_5001), .C1(n120_adj_5516), 
          .D1(n16_adj_4711), .CIN(n15514), .COUT(n15515), .S0(d6_71__N_1459[56]), 
          .S1(d6_71__N_1459[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_21 (.A0(d_tmp[54]), .B0(cout_adj_5001), .C0(n129_adj_5519), 
          .D0(n19_adj_4708), .A1(d_tmp[55]), .B1(cout_adj_5001), .C1(n126_adj_5518), 
          .D1(n18_adj_4709), .CIN(n15513), .COUT(n15514), .S0(d6_71__N_1459[54]), 
          .S1(d6_71__N_1459[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_19 (.A0(d_tmp[52]), .B0(cout_adj_5001), .C0(n135_adj_5521), 
          .D0(n21_adj_4706), .A1(d_tmp[53]), .B1(cout_adj_5001), .C1(n132_adj_5520), 
          .D1(n20_adj_4707), .CIN(n15512), .COUT(n15513), .S0(d6_71__N_1459[52]), 
          .S1(d6_71__N_1459[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_17 (.A0(d_tmp[50]), .B0(cout_adj_5001), .C0(n141_adj_5523), 
          .D0(n23_adj_4704), .A1(d_tmp[51]), .B1(cout_adj_5001), .C1(n138_adj_5522), 
          .D1(n22_adj_4705), .CIN(n15511), .COUT(n15512), .S0(d6_71__N_1459[50]), 
          .S1(d6_71__N_1459[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_15 (.A0(d_tmp[48]), .B0(cout_adj_5001), .C0(n147_adj_5525), 
          .D0(n25_adj_4702), .A1(d_tmp[49]), .B1(cout_adj_5001), .C1(n144_adj_5524), 
          .D1(n24_adj_4703), .CIN(n15510), .COUT(n15511), .S0(d6_71__N_1459[48]), 
          .S1(d6_71__N_1459[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_13 (.A0(d_tmp[46]), .B0(cout_adj_5001), .C0(n153_adj_5527), 
          .D0(n27_adj_4700), .A1(d_tmp[47]), .B1(cout_adj_5001), .C1(n150_adj_5526), 
          .D1(n26_adj_4701), .CIN(n15509), .COUT(n15510), .S0(d6_71__N_1459[46]), 
          .S1(d6_71__N_1459[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_11 (.A0(d_tmp[44]), .B0(cout_adj_5001), .C0(n159_adj_5529), 
          .D0(n29_adj_4698), .A1(d_tmp[45]), .B1(cout_adj_5001), .C1(n156_adj_5528), 
          .D1(n28_adj_4699), .CIN(n15508), .COUT(n15509), .S0(d6_71__N_1459[44]), 
          .S1(d6_71__N_1459[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_9 (.A0(d_tmp[42]), .B0(cout_adj_5001), .C0(n165_adj_5531), 
          .D0(n31_adj_4696), .A1(d_tmp[43]), .B1(cout_adj_5001), .C1(n162_adj_5530), 
          .D1(n30_adj_4697), .CIN(n15507), .COUT(n15508), .S0(d6_71__N_1459[42]), 
          .S1(d6_71__N_1459[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_7 (.A0(d_tmp[40]), .B0(cout_adj_5001), .C0(n171_adj_5533), 
          .D0(n33_adj_4694), .A1(d_tmp[41]), .B1(cout_adj_5001), .C1(n168_adj_5532), 
          .D1(n32_adj_4695), .CIN(n15506), .COUT(n15507), .S0(d6_71__N_1459[40]), 
          .S1(d6_71__N_1459[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_5 (.A0(d_tmp[38]), .B0(cout_adj_5001), .C0(n177_adj_5535), 
          .D0(n35_adj_4692), .A1(d_tmp[39]), .B1(cout_adj_5001), .C1(n174_adj_5534), 
          .D1(n34_adj_4693), .CIN(n15505), .COUT(n15506), .S0(d6_71__N_1459[38]), 
          .S1(d6_71__N_1459[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_3 (.A0(d_tmp[36]), .B0(cout_adj_5001), .C0(n183_adj_5537), 
          .D0(n37_adj_4690), .A1(d_tmp[37]), .B1(cout_adj_5001), .C1(n180_adj_5536), 
          .D1(n36_adj_4691), .CIN(n15504), .COUT(n15505), .S0(d6_71__N_1459[36]), 
          .S1(d6_71__N_1459[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1436_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1436_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5001), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15504));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1436_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1436_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1436_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_37 (.A0(d4_adj_5713[70]), .B0(cout_adj_5207), 
          .C0(n81_adj_5539), .D0(d5_adj_5714[70]), .A1(d4_adj_5713[71]), 
          .B1(cout_adj_5207), .C1(n78_adj_5538), .D1(d5_adj_5714[71]), 
          .CIN(n15499), .S0(d5_71__N_706_adj_5730[70]), .S1(d5_71__N_706_adj_5730[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_35 (.A0(d4_adj_5713[68]), .B0(cout_adj_5207), 
          .C0(n87_adj_5541), .D0(d5_adj_5714[68]), .A1(d4_adj_5713[69]), 
          .B1(cout_adj_5207), .C1(n84_adj_5540), .D1(d5_adj_5714[69]), 
          .CIN(n15498), .COUT(n15499), .S0(d5_71__N_706_adj_5730[68]), 
          .S1(d5_71__N_706_adj_5730[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_33 (.A0(d4_adj_5713[66]), .B0(cout_adj_5207), 
          .C0(n93_adj_5543), .D0(d5_adj_5714[66]), .A1(d4_adj_5713[67]), 
          .B1(cout_adj_5207), .C1(n90_adj_5542), .D1(d5_adj_5714[67]), 
          .CIN(n15497), .COUT(n15498), .S0(d5_71__N_706_adj_5730[66]), 
          .S1(d5_71__N_706_adj_5730[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_31 (.A0(d4_adj_5713[64]), .B0(cout_adj_5207), 
          .C0(n99_adj_5545), .D0(d5_adj_5714[64]), .A1(d4_adj_5713[65]), 
          .B1(cout_adj_5207), .C1(n96_adj_5544), .D1(d5_adj_5714[65]), 
          .CIN(n15496), .COUT(n15497), .S0(d5_71__N_706_adj_5730[64]), 
          .S1(d5_71__N_706_adj_5730[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_29 (.A0(d4_adj_5713[62]), .B0(cout_adj_5207), 
          .C0(n105_adj_5547), .D0(d5_adj_5714[62]), .A1(d4_adj_5713[63]), 
          .B1(cout_adj_5207), .C1(n102_adj_5546), .D1(d5_adj_5714[63]), 
          .CIN(n15495), .COUT(n15496), .S0(d5_71__N_706_adj_5730[62]), 
          .S1(d5_71__N_706_adj_5730[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_27 (.A0(d4_adj_5713[60]), .B0(cout_adj_5207), 
          .C0(n111_adj_5549), .D0(d5_adj_5714[60]), .A1(d4_adj_5713[61]), 
          .B1(cout_adj_5207), .C1(n108_adj_5548), .D1(d5_adj_5714[61]), 
          .CIN(n15494), .COUT(n15495), .S0(d5_71__N_706_adj_5730[60]), 
          .S1(d5_71__N_706_adj_5730[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_25 (.A0(d4_adj_5713[58]), .B0(cout_adj_5207), 
          .C0(n117_adj_5551), .D0(d5_adj_5714[58]), .A1(d4_adj_5713[59]), 
          .B1(cout_adj_5207), .C1(n114_adj_5550), .D1(d5_adj_5714[59]), 
          .CIN(n15493), .COUT(n15494), .S0(d5_71__N_706_adj_5730[58]), 
          .S1(d5_71__N_706_adj_5730[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_23 (.A0(d4_adj_5713[56]), .B0(cout_adj_5207), 
          .C0(n123_adj_5553), .D0(d5_adj_5714[56]), .A1(d4_adj_5713[57]), 
          .B1(cout_adj_5207), .C1(n120_adj_5552), .D1(d5_adj_5714[57]), 
          .CIN(n15492), .COUT(n15493), .S0(d5_71__N_706_adj_5730[56]), 
          .S1(d5_71__N_706_adj_5730[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_21 (.A0(d4_adj_5713[54]), .B0(cout_adj_5207), 
          .C0(n129_adj_5555), .D0(d5_adj_5714[54]), .A1(d4_adj_5713[55]), 
          .B1(cout_adj_5207), .C1(n126_adj_5554), .D1(d5_adj_5714[55]), 
          .CIN(n15491), .COUT(n15492), .S0(d5_71__N_706_adj_5730[54]), 
          .S1(d5_71__N_706_adj_5730[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_19 (.A0(d4_adj_5713[52]), .B0(cout_adj_5207), 
          .C0(n135_adj_5557), .D0(d5_adj_5714[52]), .A1(d4_adj_5713[53]), 
          .B1(cout_adj_5207), .C1(n132_adj_5556), .D1(d5_adj_5714[53]), 
          .CIN(n15490), .COUT(n15491), .S0(d5_71__N_706_adj_5730[52]), 
          .S1(d5_71__N_706_adj_5730[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_17 (.A0(d4_adj_5713[50]), .B0(cout_adj_5207), 
          .C0(n141_adj_5559), .D0(d5_adj_5714[50]), .A1(d4_adj_5713[51]), 
          .B1(cout_adj_5207), .C1(n138_adj_5558), .D1(d5_adj_5714[51]), 
          .CIN(n15489), .COUT(n15490), .S0(d5_71__N_706_adj_5730[50]), 
          .S1(d5_71__N_706_adj_5730[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_15 (.A0(d4_adj_5713[48]), .B0(cout_adj_5207), 
          .C0(n147_adj_5561), .D0(d5_adj_5714[48]), .A1(d4_adj_5713[49]), 
          .B1(cout_adj_5207), .C1(n144_adj_5560), .D1(d5_adj_5714[49]), 
          .CIN(n15488), .COUT(n15489), .S0(d5_71__N_706_adj_5730[48]), 
          .S1(d5_71__N_706_adj_5730[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_13 (.A0(d4_adj_5713[46]), .B0(cout_adj_5207), 
          .C0(n153_adj_5563), .D0(d5_adj_5714[46]), .A1(d4_adj_5713[47]), 
          .B1(cout_adj_5207), .C1(n150_adj_5562), .D1(d5_adj_5714[47]), 
          .CIN(n15487), .COUT(n15488), .S0(d5_71__N_706_adj_5730[46]), 
          .S1(d5_71__N_706_adj_5730[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_11 (.A0(d4_adj_5713[44]), .B0(cout_adj_5207), 
          .C0(n159_adj_5565), .D0(d5_adj_5714[44]), .A1(d4_adj_5713[45]), 
          .B1(cout_adj_5207), .C1(n156_adj_5564), .D1(d5_adj_5714[45]), 
          .CIN(n15486), .COUT(n15487), .S0(d5_71__N_706_adj_5730[44]), 
          .S1(d5_71__N_706_adj_5730[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_9 (.A0(d4_adj_5713[42]), .B0(cout_adj_5207), 
          .C0(n165_adj_5567), .D0(d5_adj_5714[42]), .A1(d4_adj_5713[43]), 
          .B1(cout_adj_5207), .C1(n162_adj_5566), .D1(d5_adj_5714[43]), 
          .CIN(n15485), .COUT(n15486), .S0(d5_71__N_706_adj_5730[42]), 
          .S1(d5_71__N_706_adj_5730[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_7 (.A0(d4_adj_5713[40]), .B0(cout_adj_5207), 
          .C0(n171_adj_5569), .D0(d5_adj_5714[40]), .A1(d4_adj_5713[41]), 
          .B1(cout_adj_5207), .C1(n168_adj_5568), .D1(d5_adj_5714[41]), 
          .CIN(n15484), .COUT(n15485), .S0(d5_71__N_706_adj_5730[40]), 
          .S1(d5_71__N_706_adj_5730[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_5 (.A0(d4_adj_5713[38]), .B0(cout_adj_5207), 
          .C0(n177_adj_5571), .D0(d5_adj_5714[38]), .A1(d4_adj_5713[39]), 
          .B1(cout_adj_5207), .C1(n174_adj_5570), .D1(d5_adj_5714[39]), 
          .CIN(n15483), .COUT(n15484), .S0(d5_71__N_706_adj_5730[38]), 
          .S1(d5_71__N_706_adj_5730[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_3 (.A0(d4_adj_5713[36]), .B0(cout_adj_5207), 
          .C0(n183_adj_5573), .D0(d5_adj_5714[36]), .A1(d4_adj_5713[37]), 
          .B1(cout_adj_5207), .C1(n180_adj_5572), .D1(d5_adj_5714[37]), 
          .CIN(n15482), .COUT(n15483), .S0(d5_71__N_706_adj_5730[36]), 
          .S1(d5_71__N_706_adj_5730[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1439_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1439_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5207), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15482));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1439_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1439_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_13 (.A0(LOCosine[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15478), .S0(MixerOutCos_11__N_250[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1406_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_1406_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_1406_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_11 (.A0(LOCosine[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15477), .COUT(n15478), .S0(MixerOutCos_11__N_250[9]), 
          .S1(MixerOutCos_11__N_250[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1406_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_1406_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_1406_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_9 (.A0(LOCosine[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15476), .COUT(n15477), .S0(MixerOutCos_11__N_250[7]), 
          .S1(MixerOutCos_11__N_250[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1406_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_1406_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_1406_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_7 (.A0(LOCosine[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15475), .COUT(n15476), .S0(MixerOutCos_11__N_250[5]), 
          .S1(MixerOutCos_11__N_250[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1406_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_1406_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_1406_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_5 (.A0(LOCosine[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15474), .COUT(n15475), .S0(MixerOutCos_11__N_250[3]), 
          .S1(MixerOutCos_11__N_250[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1406_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_1406_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_1406_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_3 (.A0(LOCosine[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15473), .COUT(n15474), .S0(MixerOutCos_11__N_250[1]), 
          .S1(MixerOutCos_11__N_250[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1406_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_1406_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_1406_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15473), .S1(MixerOutCos_11__N_250[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1406_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1406_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_1406_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_38 (.A0(d4[71]), .B0(d3[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15472), .S0(n78_adj_5249));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1535_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_36 (.A0(d4[69]), .B0(d3[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[70]), .B1(d3[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15471), .COUT(n15472), .S0(n84_adj_5251), .S1(n81_adj_5250));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_34 (.A0(d4[67]), .B0(d3[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[68]), .B1(d3[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15470), .COUT(n15471), .S0(n90_adj_5253), .S1(n87_adj_5252));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_32 (.A0(d4[65]), .B0(d3[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[66]), .B1(d3[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15469), .COUT(n15470), .S0(n96_adj_5255), .S1(n93_adj_5254));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_30 (.A0(d4[63]), .B0(d3[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[64]), .B1(d3[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15468), .COUT(n15469), .S0(n102_adj_5257), .S1(n99_adj_5256));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_28 (.A0(d4[61]), .B0(d3[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[62]), .B1(d3[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15467), .COUT(n15468), .S0(n108_adj_5259), .S1(n105_adj_5258));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_26 (.A0(d4[59]), .B0(d3[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[60]), .B1(d3[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15466), .COUT(n15467), .S0(n114_adj_5261), .S1(n111_adj_5260));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_24 (.A0(d4[57]), .B0(d3[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[58]), .B1(d3[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15465), .COUT(n15466), .S0(n120_adj_5263), .S1(n117_adj_5262));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_22 (.A0(d4[55]), .B0(d3[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[56]), .B1(d3[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15464), .COUT(n15465), .S0(n126_adj_5265), .S1(n123_adj_5264));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_20 (.A0(d4[53]), .B0(d3[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[54]), .B1(d3[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15463), .COUT(n15464), .S0(n132_adj_5267), .S1(n129_adj_5266));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_18 (.A0(d4[51]), .B0(d3[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[52]), .B1(d3[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15462), .COUT(n15463), .S0(n138_adj_5269), .S1(n135_adj_5268));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_16 (.A0(d4[49]), .B0(d3[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[50]), .B1(d3[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15461), .COUT(n15462), .S0(n144_adj_5271), .S1(n141_adj_5270));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_14 (.A0(d4[47]), .B0(d3[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[48]), .B1(d3[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15460), .COUT(n15461), .S0(n150_adj_5273), .S1(n147_adj_5272));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_12 (.A0(d4[45]), .B0(d3[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[46]), .B1(d3[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15459), .COUT(n15460), .S0(n156_adj_5275), .S1(n153_adj_5274));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_10 (.A0(d4[43]), .B0(d3[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[44]), .B1(d3[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15458), .COUT(n15459), .S0(n162_adj_5277), .S1(n159_adj_5276));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_8 (.A0(d4[41]), .B0(d3[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[42]), .B1(d3[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15457), .COUT(n15458), .S0(n168_adj_5279), .S1(n165_adj_5278));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_6 (.A0(d4[39]), .B0(d3[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[40]), .B1(d3[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15456), .COUT(n15457), .S0(n174_adj_5281), .S1(n171_adj_5280));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_6.INJECT1_1 = "NO";
    LUT4 i5034_1_lut_2_lut_3_lut (.A(ISquare[23]), .B(ISquare[22]), .C(ISquare[31]), 
         .Z(n23_adj_5022)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam i5034_1_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 i1_2_lut_rep_204_3_lut (.A(ISquare[23]), .B(ISquare[22]), .C(ISquare[31]), 
         .Z(n17826)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam i1_2_lut_rep_204_3_lut.init = 16'hfefe;
    LUT4 i2351_3_lut (.A(led_c_1), .B(n238), .C(n18053), .Z(n12254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2351_3_lut.init = 16'hcaca;
    CCU2C _add_1_1535_add_4_4 (.A0(d4[37]), .B0(d3[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[38]), .B1(d3[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15455), .COUT(n15456), .S0(n180_adj_5283), .S1(n177_adj_5282));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1535_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1535_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[36]), .B1(d3[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15455), .S1(n183_adj_5284));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1535_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1535_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1535_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1535_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_38 (.A0(d_d8[71]), .B0(d8[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15454), .S0(n78_adj_4575));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1577_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_36 (.A0(d_d8[69]), .B0(d8[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[70]), .B1(d8[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15453), .COUT(n15454), .S0(n84_adj_4573), .S1(n81_adj_4574));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_34 (.A0(d_d8[67]), .B0(d8[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[68]), .B1(d8[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15452), .COUT(n15453), .S0(n90_adj_4571), .S1(n87_adj_4572));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_32 (.A0(d_d8[65]), .B0(d8[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[66]), .B1(d8[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15451), .COUT(n15452), .S0(n96_adj_4569), .S1(n93_adj_4570));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_30 (.A0(d_d8[63]), .B0(d8[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[64]), .B1(d8[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15450), .COUT(n15451), .S0(n102_adj_4567), .S1(n99_adj_4568));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_28 (.A0(d_d8[61]), .B0(d8[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[62]), .B1(d8[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15449), .COUT(n15450), .S0(n108_adj_4565), .S1(n105_adj_4566));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_26 (.A0(d_d8[59]), .B0(d8[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[60]), .B1(d8[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15448), .COUT(n15449), .S0(n114_adj_4563), .S1(n111_adj_4564));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_24 (.A0(d_d8[57]), .B0(d8[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[58]), .B1(d8[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15447), .COUT(n15448), .S0(n120_adj_4561), .S1(n117_adj_4562));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_22 (.A0(d_d8[55]), .B0(d8[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[56]), .B1(d8[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15446), .COUT(n15447), .S0(n126), .S1(n123));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_20 (.A0(d_d8[53]), .B0(d8[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[54]), .B1(d8[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15445), .COUT(n15446), .S0(n132), .S1(n129));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_18 (.A0(d_d8[51]), .B0(d8[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[52]), .B1(d8[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15444), .COUT(n15445), .S0(n138), .S1(n135));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_16 (.A0(d_d8[49]), .B0(d8[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[50]), .B1(d8[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15443), .COUT(n15444), .S0(n144), .S1(n141));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_14 (.A0(d_d8[47]), .B0(d8[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[48]), .B1(d8[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15442), .COUT(n15443), .S0(n150), .S1(n147));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_12 (.A0(d_d8[45]), .B0(d8[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[46]), .B1(d8[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15441), .COUT(n15442), .S0(n156), .S1(n153));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_10 (.A0(d_d8[43]), .B0(d8[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[44]), .B1(d8[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15440), .COUT(n15441), .S0(n162), .S1(n159));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_8 (.A0(d_d8[41]), .B0(d8[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[42]), .B1(d8[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15439), .COUT(n15440), .S0(n168), .S1(n165));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_6 (.A0(d_d8[39]), .B0(d8[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[40]), .B1(d8[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15438), .COUT(n15439), .S0(n174), .S1(n171));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_4 (.A0(d_d8[37]), .B0(d8[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[38]), .B1(d8[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15437), .COUT(n15438), .S0(n180), .S1(n177));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1577_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1577_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[36]), .B1(d8[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15437), .S1(n183));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1577_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1577_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1577_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1577_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_38 (.A0(d5[71]), .B0(d4[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15436), .S0(n78_adj_5285));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1538_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_36 (.A0(d5[69]), .B0(d4[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[70]), .B1(d4[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15435), .COUT(n15436), .S0(n84_adj_5287), .S1(n81_adj_5286));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_34 (.A0(d5[67]), .B0(d4[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[68]), .B1(d4[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15434), .COUT(n15435), .S0(n90_adj_5289), .S1(n87_adj_5288));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_32 (.A0(d5[65]), .B0(d4[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[66]), .B1(d4[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15433), .COUT(n15434), .S0(n96_adj_5291), .S1(n93_adj_5290));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_30 (.A0(d5[63]), .B0(d4[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[64]), .B1(d4[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15432), .COUT(n15433), .S0(n102_adj_5293), .S1(n99_adj_5292));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_28 (.A0(d5[61]), .B0(d4[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[62]), .B1(d4[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15431), .COUT(n15432), .S0(n108_adj_5295), .S1(n105_adj_5294));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_26 (.A0(d5[59]), .B0(d4[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[60]), .B1(d4[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15430), .COUT(n15431), .S0(n114_adj_5297), .S1(n111_adj_5296));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_24 (.A0(d5[57]), .B0(d4[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[58]), .B1(d4[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15429), .COUT(n15430), .S0(n120_adj_5299), .S1(n117_adj_5298));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_22 (.A0(d5[55]), .B0(d4[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[56]), .B1(d4[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15428), .COUT(n15429), .S0(n126_adj_5301), .S1(n123_adj_5300));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_20 (.A0(d5[53]), .B0(d4[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[54]), .B1(d4[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15427), .COUT(n15428), .S0(n132_adj_5303), .S1(n129_adj_5302));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_18 (.A0(d5[51]), .B0(d4[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[52]), .B1(d4[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15426), .COUT(n15427), .S0(n138_adj_5305), .S1(n135_adj_5304));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_16 (.A0(d5[49]), .B0(d4[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[50]), .B1(d4[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15425), .COUT(n15426), .S0(n144_adj_5307), .S1(n141_adj_5306));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_14 (.A0(d5[47]), .B0(d4[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[48]), .B1(d4[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15424), .COUT(n15425), .S0(n150_adj_5309), .S1(n147_adj_5308));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_12 (.A0(d5[45]), .B0(d4[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[46]), .B1(d4[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15423), .COUT(n15424), .S0(n156_adj_5311), .S1(n153_adj_5310));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_12.INJECT1_1 = "NO";
    FD1P3AX phase_inc_carrGen_i0_i1 (.D(n1993), .SP(clk_80mhz_enable_1387), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i1.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i3 (.D(n12542), .SP(clk_80mhz_enable_1388), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i3.GSR = "ENABLED";
    LUT4 i5018_2_lut_3_lut (.A(ISquare[23]), .B(ISquare[22]), .C(ISquare[31]), 
         .Z(n14967)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam i5018_2_lut_3_lut.init = 16'h0e0e;
    FD1P3AX phase_inc_carrGen_i0_i5 (.D(n1989), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i5.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i7 (.D(n1987), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i7.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i11 (.D(n1983), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i11.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i15 (.D(n1979), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i15.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i19 (.D(n1975), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i19.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i21 (.D(n1973), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i21.GSR = "ENABLED";
    LUT4 i2074_3_lut_4_lut (.A(n17823), .B(n16869), .C(led_c_0), .D(n286_adj_5076), 
         .Z(n11968)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i2074_3_lut_4_lut.init = 16'hf780;
    LUT4 i19_4_lut_adj_70 (.A(n190_adj_5044), .B(n196), .C(n18053), .D(n17814), 
         .Z(n8_adj_4739)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i19_4_lut_adj_70.init = 16'hc0ca;
    FD1P3AX phase_inc_carrGen_i0_i24 (.D(n1970), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i24.GSR = "ENABLED";
    LUT4 i2082_3_lut_4_lut (.A(n17823), .B(n16869), .C(led_c_0), .D(n253_adj_5065), 
         .Z(n11976)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i2082_3_lut_4_lut.init = 16'hf780;
    FD1P3AX phase_inc_carrGen_i0_i26 (.D(n1968), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i26.GSR = "ENABLED";
    LUT4 mux_305_i43_4_lut (.A(n197), .B(n11995), .C(n17815), .D(n17809), 
         .Z(n1952)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i43_4_lut.init = 16'h0aca;
    FD1P3AX phase_inc_carrGen_i0_i30 (.D(n1964), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i30.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i32 (.D(n1962), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i32.GSR = "ENABLED";
    LUT4 i5008_1_lut_2_lut (.A(ISquare[23]), .B(ISquare[22]), .Z(n32_adj_5023)) /* synthesis lut_function=(!(A+(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam i5008_1_lut_2_lut.init = 16'h1111;
    FD1P3AX phase_inc_carrGen_i0_i34 (.D(n1960), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i34.GSR = "ENABLED";
    LUT4 i2101_3_lut (.A(n11994), .B(n193), .C(led_c_4), .Z(n11995)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2101_3_lut.init = 16'hcaca;
    LUT4 i2096_3_lut_4_lut (.A(n17823), .B(n16869), .C(led_c_0), .D(n202_adj_5048), 
         .Z(n11990)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i2096_3_lut_4_lut.init = 16'hf780;
    FD1P3AX phase_inc_carrGen_i0_i41 (.D(n1953), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i41.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i42 (.D(n1952), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[42]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i42.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i43 (.D(n1951), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i43.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i44 (.D(n1950), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[44]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i44.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i47 (.D(n1947), .SP(clk_80mhz_enable_1411), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i47.GSR = "ENABLED";
    LUT4 mux_305_i44_4_lut (.A(n194), .B(n2602), .C(n17815), .D(n17809), 
         .Z(n1951)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i44_4_lut.init = 16'h0aca;
    LUT4 led_c_0_bdd_4_lut (.A(led_c_0), .B(led_c_3), .C(led_c_2), .D(led_c_1), 
         .Z(n17778)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A !(B (C (D))+!B (D)))) */ ;
    defparam led_c_0_bdd_4_lut.init = 16'h7102;
    LUT4 i2104_3_lut_4_lut (.A(n17823), .B(n16869), .C(led_c_0), .D(n175_adj_5039), 
         .Z(n11998)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i2104_3_lut_4_lut.init = 16'hf780;
    FD1P3AX phase_inc_carrGen_i0_i52 (.D(n1942), .SP(o_Rx_DV), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen[52]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i52.GSR = "ENABLED";
    LUT4 mux_305_i45_4_lut (.A(n191), .B(n11997), .C(n17815), .D(n17809), 
         .Z(n1950)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i45_4_lut.init = 16'h0aca;
    LUT4 i3177_4_lut_4_lut (.A(led_c_4), .B(n17817), .C(n211), .D(n205_adj_5049), 
         .Z(n2609)) /* synthesis lut_function=(A (C)+!A !(B+!(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3177_4_lut_4_lut.init = 16'hb1a0;
    FD1P3AX phase_inc_carrGen_i0_i57 (.D(n1937), .SP(o_Rx_DV), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i57.GSR = "ENABLED";
    LUT4 i2103_3_lut (.A(n11996), .B(n187), .C(led_c_4), .Z(n11997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2103_3_lut.init = 16'hcaca;
    FD1P3AX phase_inc_carrGen_i0_i59 (.D(n1935), .SP(o_Rx_DV), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i59.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i60 (.D(n1934), .SP(o_Rx_DV), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen[60]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i60.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i61 (.D(n1933), .SP(o_Rx_DV), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i61.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i62 (.D(n1932), .SP(o_Rx_DV), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen[62]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i62.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i63 (.D(n1931), .SP(o_Rx_DV), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i63.GSR = "ENABLED";
    CCU2C _add_1_1472_add_4_30 (.A0(d_d8_adj_5720[27]), .B0(d8_adj_5719[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[28]), .B1(d8_adj_5719[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15916), .COUT(n15917), .S0(d9_71__N_1675_adj_5745[27]), 
          .S1(d9_71__N_1675_adj_5745[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_28 (.A0(d_d8_adj_5720[25]), .B0(d8_adj_5719[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[26]), .B1(d8_adj_5719[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15915), .COUT(n15916), .S0(d9_71__N_1675_adj_5745[25]), 
          .S1(d9_71__N_1675_adj_5745[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_26 (.A0(d_d8_adj_5720[23]), .B0(d8_adj_5719[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[24]), .B1(d8_adj_5719[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15914), .COUT(n15915), .S0(d9_71__N_1675_adj_5745[23]), 
          .S1(d9_71__N_1675_adj_5745[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_24 (.A0(d_d8_adj_5720[21]), .B0(d8_adj_5719[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[22]), .B1(d8_adj_5719[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15913), .COUT(n15914), .S0(d9_71__N_1675_adj_5745[21]), 
          .S1(d9_71__N_1675_adj_5745[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_22 (.A0(d_d8_adj_5720[19]), .B0(d8_adj_5719[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[20]), .B1(d8_adj_5719[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15912), .COUT(n15913), .S0(d9_71__N_1675_adj_5745[19]), 
          .S1(d9_71__N_1675_adj_5745[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_20 (.A0(d_d8_adj_5720[17]), .B0(d8_adj_5719[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[18]), .B1(d8_adj_5719[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15911), .COUT(n15912), .S0(d9_71__N_1675_adj_5745[17]), 
          .S1(d9_71__N_1675_adj_5745[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_18 (.A0(d_d8_adj_5720[15]), .B0(d8_adj_5719[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[16]), .B1(d8_adj_5719[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15910), .COUT(n15911), .S0(d9_71__N_1675_adj_5745[15]), 
          .S1(d9_71__N_1675_adj_5745[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_16 (.A0(d_d8_adj_5720[13]), .B0(d8_adj_5719[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[14]), .B1(d8_adj_5719[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15909), .COUT(n15910), .S0(d9_71__N_1675_adj_5745[13]), 
          .S1(d9_71__N_1675_adj_5745[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_14 (.A0(d_d8_adj_5720[11]), .B0(d8_adj_5719[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[12]), .B1(d8_adj_5719[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15908), .COUT(n15909), .S0(d9_71__N_1675_adj_5745[11]), 
          .S1(d9_71__N_1675_adj_5745[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_12 (.A0(d_d8_adj_5720[9]), .B0(d8_adj_5719[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[10]), .B1(d8_adj_5719[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15907), .COUT(n15908), .S0(d9_71__N_1675_adj_5745[9]), 
          .S1(d9_71__N_1675_adj_5745[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_10 (.A0(d_d8_adj_5720[7]), .B0(d8_adj_5719[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[8]), .B1(d8_adj_5719[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15906), .COUT(n15907), .S0(d9_71__N_1675_adj_5745[7]), 
          .S1(d9_71__N_1675_adj_5745[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_8 (.A0(d_d8_adj_5720[5]), .B0(d8_adj_5719[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[6]), .B1(d8_adj_5719[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15905), .COUT(n15906), .S0(d9_71__N_1675_adj_5745[5]), 
          .S1(d9_71__N_1675_adj_5745[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_6 (.A0(d_d8_adj_5720[3]), .B0(d8_adj_5719[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[4]), .B1(d8_adj_5719[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15904), .COUT(n15905), .S0(d9_71__N_1675_adj_5745[3]), 
          .S1(d9_71__N_1675_adj_5745[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_4 (.A0(d_d8_adj_5720[1]), .B0(d8_adj_5719[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[2]), .B1(d8_adj_5719[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15903), .COUT(n15904), .S0(d9_71__N_1675_adj_5745[1]), 
          .S1(d9_71__N_1675_adj_5745[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1472_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1472_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8_adj_5720[0]), .B1(d8_adj_5719[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15903), .S1(d9_71__N_1675_adj_5745[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1472_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1472_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1472_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1472_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_38 (.A0(d2[71]), .B0(d1[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15902), .S0(n78_adj_5118));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1529_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_36 (.A0(d2[69]), .B0(d1[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[70]), .B1(d1[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15901), .COUT(n15902), .S0(n84_adj_5120), .S1(n81_adj_5119));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_34 (.A0(d2[67]), .B0(d1[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[68]), .B1(d1[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15900), .COUT(n15901), .S0(n90_adj_5122), .S1(n87_adj_5121));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_32 (.A0(d2[65]), .B0(d1[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[66]), .B1(d1[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15899), .COUT(n15900), .S0(n96_adj_5124), .S1(n93_adj_5123));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_30 (.A0(d2[63]), .B0(d1[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[64]), .B1(d1[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15898), .COUT(n15899), .S0(n102_adj_5126), .S1(n99_adj_5125));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_28 (.A0(d2[61]), .B0(d1[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[62]), .B1(d1[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15897), .COUT(n15898), .S0(n108_adj_5128), .S1(n105_adj_5127));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_26 (.A0(d2[59]), .B0(d1[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[60]), .B1(d1[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15896), .COUT(n15897), .S0(n114_adj_5130), .S1(n111_adj_5129));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_24 (.A0(d2[57]), .B0(d1[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[58]), .B1(d1[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15895), .COUT(n15896), .S0(n120_adj_5132), .S1(n117_adj_5131));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_22 (.A0(d2[55]), .B0(d1[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[56]), .B1(d1[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15894), .COUT(n15895), .S0(n126_adj_5134), .S1(n123_adj_5133));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_20 (.A0(d2[53]), .B0(d1[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[54]), .B1(d1[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15893), .COUT(n15894), .S0(n132_adj_5136), .S1(n129_adj_5135));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_18 (.A0(d2[51]), .B0(d1[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[52]), .B1(d1[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15892), .COUT(n15893), .S0(n138_adj_5138), .S1(n135_adj_5137));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_16 (.A0(d2[49]), .B0(d1[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[50]), .B1(d1[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15891), .COUT(n15892), .S0(n144_adj_5140), .S1(n141_adj_5139));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_14 (.A0(d2[47]), .B0(d1[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[48]), .B1(d1[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15890), .COUT(n15891), .S0(n150_adj_5142), .S1(n147_adj_5141));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_12 (.A0(d2[45]), .B0(d1[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[46]), .B1(d1[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15889), .COUT(n15890), .S0(n156_adj_5144), .S1(n153_adj_5143));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_10 (.A0(d2[43]), .B0(d1[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[44]), .B1(d1[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15888), .COUT(n15889), .S0(n162_adj_5146), .S1(n159_adj_5145));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_8 (.A0(d2[41]), .B0(d1[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[42]), .B1(d1[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15887), .COUT(n15888), .S0(n168_adj_5148), .S1(n165_adj_5147));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_6 (.A0(d2[39]), .B0(d1[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[40]), .B1(d1[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15886), .COUT(n15887), .S0(n174_adj_5150), .S1(n171_adj_5149));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_4 (.A0(d2[37]), .B0(d1[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[38]), .B1(d1[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15885), .COUT(n15886), .S0(n180_adj_5152), .S1(n177_adj_5151));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1529_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1529_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[36]), .B1(d1[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15885), .S1(n183_adj_5153));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1529_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1529_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1529_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1529_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_20 (.A0(n916), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15884), .S0(d_out_d_11__N_2383[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1466_add_4_20.INIT0 = 16'h555f;
    defparam _add_1_1466_add_4_20.INIT1 = 16'h0000;
    defparam _add_1_1466_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_18 (.A0(ISquare[31]), .B0(n918), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(n917), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15883), .COUT(n15884));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1466_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1466_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1466_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_16 (.A0(n920), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(n919), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15882), .COUT(n15883));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1466_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1466_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1466_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_14 (.A0(d_out_d_11__N_1874[17]), .B0(n922), 
          .C0(GND_net), .D0(VCC_net), .A1(ISquare[31]), .B1(n17828), 
          .C1(n921), .D1(VCC_net), .CIN(n15881), .COUT(n15882));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1466_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1466_add_4_14.INIT1 = 16'he1e1;
    defparam _add_1_1466_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_12 (.A0(d_out_d_11__N_1878[17]), .B0(n924), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n923), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15880), .COUT(n15881));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1466_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1466_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1466_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_10 (.A0(d_out_d_11__N_1882[17]), .B0(n926), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n925), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15879), .COUT(n15880));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1466_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1466_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1466_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_8 (.A0(d_out_d_11__N_1886[17]), .B0(n928), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n927), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15878), .COUT(n15879));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1466_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1466_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1466_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_6 (.A0(d_out_d_11__N_1890[17]), .B0(n930), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n929), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15877), .COUT(n15878));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1466_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1466_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1466_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_4 (.A0(d_out_d_11__N_1892[17]), .B0(ISquare[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1892[17]), .B1(n931), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15876), .COUT(n15877));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1466_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1466_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1466_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1466_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15876));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1466_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1466_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1466_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1466_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_38 (.A0(d_d9_adj_5722[35]), .B0(d9_adj_5721[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15875), .S1(cout_adj_2808));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1469_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_36 (.A0(d_d9_adj_5722[33]), .B0(d9_adj_5721[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[34]), .B1(d9_adj_5721[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15874), .COUT(n15875));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_34 (.A0(d_d9_adj_5722[31]), .B0(d9_adj_5721[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[32]), .B1(d9_adj_5721[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15873), .COUT(n15874));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_32 (.A0(d_d9_adj_5722[29]), .B0(d9_adj_5721[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[30]), .B1(d9_adj_5721[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15872), .COUT(n15873));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_30 (.A0(d_d9_adj_5722[27]), .B0(d9_adj_5721[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[28]), .B1(d9_adj_5721[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15871), .COUT(n15872));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_28 (.A0(d_d9_adj_5722[25]), .B0(d9_adj_5721[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[26]), .B1(d9_adj_5721[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15870), .COUT(n15871));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_26 (.A0(d_d9_adj_5722[23]), .B0(d9_adj_5721[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[24]), .B1(d9_adj_5721[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15869), .COUT(n15870));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_24 (.A0(d_d9_adj_5722[21]), .B0(d9_adj_5721[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[22]), .B1(d9_adj_5721[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15868), .COUT(n15869));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_22 (.A0(d_d9_adj_5722[19]), .B0(d9_adj_5721[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[20]), .B1(d9_adj_5721[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15867), .COUT(n15868));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_20 (.A0(d_d9_adj_5722[17]), .B0(d9_adj_5721[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[18]), .B1(d9_adj_5721[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15866), .COUT(n15867));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_18 (.A0(d_d9_adj_5722[15]), .B0(d9_adj_5721[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[16]), .B1(d9_adj_5721[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15865), .COUT(n15866));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_16 (.A0(d_d9_adj_5722[13]), .B0(d9_adj_5721[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[14]), .B1(d9_adj_5721[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15864), .COUT(n15865));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_14 (.A0(d_d9_adj_5722[11]), .B0(d9_adj_5721[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[12]), .B1(d9_adj_5721[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15863), .COUT(n15864));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_12 (.A0(d_d9_adj_5722[9]), .B0(d9_adj_5721[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[10]), .B1(d9_adj_5721[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15862), .COUT(n15863));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_10 (.A0(d_d9_adj_5722[7]), .B0(d9_adj_5721[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[8]), .B1(d9_adj_5721[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15861), .COUT(n15862));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_8 (.A0(d_d9_adj_5722[5]), .B0(d9_adj_5721[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[6]), .B1(d9_adj_5721[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15860), .COUT(n15861));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_6 (.A0(d_d9_adj_5722[3]), .B0(d9_adj_5721[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[4]), .B1(d9_adj_5721[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15859), .COUT(n15860));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_4 (.A0(d_d9_adj_5722[1]), .B0(d9_adj_5721[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[2]), .B1(d9_adj_5721[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15858), .COUT(n15859));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1469_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1469_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9_adj_5722[0]), .B1(d9_adj_5721[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15858));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1469_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1469_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1469_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1469_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_28 (.A0(d_d_tmp_adj_5709[25]), .B0(d_tmp_adj_5708[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[26]), .B1(d_tmp_adj_5708[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16277), .COUT(n16278), .S0(d6_71__N_1459_adj_5742[25]), 
          .S1(d6_71__N_1459_adj_5742[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_28.INJECT1_1 = "NO";
    LUT4 mux_305_i48_4_lut (.A(n182), .B(n2598), .C(n17815), .D(n17809), 
         .Z(n1947)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i48_4_lut.init = 16'h0aca;
    CCU2C _add_1_1481_add_4_26 (.A0(d_d_tmp_adj_5709[23]), .B0(d_tmp_adj_5708[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[24]), .B1(d_tmp_adj_5708[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16276), .COUT(n16277), .S0(d6_71__N_1459_adj_5742[23]), 
          .S1(d6_71__N_1459_adj_5742[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_24 (.A0(d_d_tmp_adj_5709[21]), .B0(d_tmp_adj_5708[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[22]), .B1(d_tmp_adj_5708[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16275), .COUT(n16276), .S0(d6_71__N_1459_adj_5742[21]), 
          .S1(d6_71__N_1459_adj_5742[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_24.INJECT1_1 = "NO";
    LUT4 i19_4_lut_adj_71 (.A(n157_adj_5033), .B(n163), .C(led_c_4), .D(n17814), 
         .Z(n8_adj_4729)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i19_4_lut_adj_71.init = 16'hc0ca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n17823), .B(n16869), .C(n12538), .D(n18053), 
         .Z(n17069)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0007;
    CCU2C _add_1_1481_add_4_22 (.A0(d_d_tmp_adj_5709[19]), .B0(d_tmp_adj_5708[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[20]), .B1(d_tmp_adj_5708[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16274), .COUT(n16275), .S0(d6_71__N_1459_adj_5742[19]), 
          .S1(d6_71__N_1459_adj_5742[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_22.INJECT1_1 = "NO";
    LUT4 i19_4_lut_adj_72 (.A(n142_adj_5028), .B(n148), .C(n18053), .D(n17814), 
         .Z(n8_adj_4726)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i19_4_lut_adj_72.init = 16'hc0ca;
    LUT4 mux_305_i60_4_lut (.A(n146), .B(n2586), .C(n17815), .D(n17809), 
         .Z(n1935)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i60_4_lut.init = 16'h0aca;
    LUT4 mux_305_i61_4_lut (.A(n143), .B(n2585), .C(n17815), .D(n17809), 
         .Z(n1934)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i61_4_lut.init = 16'h0aca;
    CCU2C _add_1_1481_add_4_20 (.A0(d_d_tmp_adj_5709[17]), .B0(d_tmp_adj_5708[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[18]), .B1(d_tmp_adj_5708[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16273), .COUT(n16274), .S0(d6_71__N_1459_adj_5742[17]), 
          .S1(d6_71__N_1459_adj_5742[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_18 (.A0(d_d_tmp_adj_5709[15]), .B0(d_tmp_adj_5708[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[16]), .B1(d_tmp_adj_5708[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16272), .COUT(n16273), .S0(d6_71__N_1459_adj_5742[15]), 
          .S1(d6_71__N_1459_adj_5742[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_18.INJECT1_1 = "NO";
    LUT4 i2110_3_lut_4_lut (.A(n17823), .B(n16869), .C(led_c_0), .D(n154_adj_5032), 
         .Z(n12004)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i2110_3_lut_4_lut.init = 16'hf780;
    CCU2C _add_1_1481_add_4_16 (.A0(d_d_tmp_adj_5709[13]), .B0(d_tmp_adj_5708[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[14]), .B1(d_tmp_adj_5708[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16271), .COUT(n16272), .S0(d6_71__N_1459_adj_5742[13]), 
          .S1(d6_71__N_1459_adj_5742[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_14 (.A0(d_d_tmp_adj_5709[11]), .B0(d_tmp_adj_5708[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[12]), .B1(d_tmp_adj_5708[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16270), .COUT(n16271), .S0(d6_71__N_1459_adj_5742[11]), 
          .S1(d6_71__N_1459_adj_5742[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_12 (.A0(d_d_tmp_adj_5709[9]), .B0(d_tmp_adj_5708[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[10]), .B1(d_tmp_adj_5708[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16269), .COUT(n16270), .S0(d6_71__N_1459_adj_5742[9]), 
          .S1(d6_71__N_1459_adj_5742[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_12.INJECT1_1 = "NO";
    LUT4 i19_4_lut_adj_73 (.A(n130_adj_5024), .B(n136), .C(n18053), .D(n17814), 
         .Z(n8_adj_4730)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i19_4_lut_adj_73.init = 16'hc0ca;
    LUT4 i19_4_lut_adj_74 (.A(n127), .B(n133), .C(led_c_4), .D(n17814), 
         .Z(n8_adj_4727)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i19_4_lut_adj_74.init = 16'hc0ca;
    LUT4 i2084_3_lut_4_lut (.A(n17823), .B(n16869), .C(led_c_0), .D(n247_adj_5063), 
         .Z(n11978)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i2084_3_lut_4_lut.init = 16'hf780;
    LUT4 i19_4_lut_adj_75 (.A(n124), .B(n130), .C(n18053), .D(n17814), 
         .Z(n8_adj_4728)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i19_4_lut_adj_75.init = 16'hc0ca;
    CCU2C _add_1_1481_add_4_10 (.A0(d_d_tmp_adj_5709[7]), .B0(d_tmp_adj_5708[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[8]), .B1(d_tmp_adj_5708[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16268), .COUT(n16269), .S0(d6_71__N_1459_adj_5742[7]), 
          .S1(d6_71__N_1459_adj_5742[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_8 (.A0(d_d_tmp_adj_5709[5]), .B0(d_tmp_adj_5708[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[6]), .B1(d_tmp_adj_5708[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16267), .COUT(n16268), .S0(d6_71__N_1459_adj_5742[5]), 
          .S1(d6_71__N_1459_adj_5742[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_6 (.A0(d_d_tmp_adj_5709[3]), .B0(d_tmp_adj_5708[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[4]), .B1(d_tmp_adj_5708[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16266), .COUT(n16267), .S0(d6_71__N_1459_adj_5742[3]), 
          .S1(d6_71__N_1459_adj_5742[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1481_add_4_4 (.A0(d_d_tmp_adj_5709[1]), .B0(d_tmp_adj_5708[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[2]), .B1(d_tmp_adj_5708[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16265), .COUT(n16266), .S0(d6_71__N_1459_adj_5742[1]), 
          .S1(d6_71__N_1459_adj_5742[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1481_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_4.INJECT1_1 = "NO";
    LUT4 i6026_4_lut (.A(n17075), .B(n17022), .C(n17073), .D(n17778), 
         .Z(n12538)) /* synthesis lut_function=(!(A (B+(C (D))))) */ ;
    defparam i6026_4_lut.init = 16'h5777;
    CCU2C _add_1_1481_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp_adj_5709[0]), .B1(d_tmp_adj_5708[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16265), .S1(d6_71__N_1459_adj_5742[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1481_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1481_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1481_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1481_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_38 (.A0(d_d6_adj_5716[35]), .B0(d6_adj_5715[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16264), .S0(d7_71__N_1531_adj_5743[35]), 
          .S1(cout_adj_5464));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1478_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_36 (.A0(d_d6_adj_5716[33]), .B0(d6_adj_5715[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[34]), .B1(d6_adj_5715[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16263), .COUT(n16264), .S0(d7_71__N_1531_adj_5743[33]), 
          .S1(d7_71__N_1531_adj_5743[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_36.INJECT1_1 = "NO";
    LUT4 i2640_3_lut (.A(n305), .B(n2707), .C(n12538), .Z(n12545)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2640_3_lut.init = 16'hacac;
    CCU2C _add_1_1478_add_4_34 (.A0(d_d6_adj_5716[31]), .B0(d6_adj_5715[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[32]), .B1(d6_adj_5715[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16262), .COUT(n16263), .S0(d7_71__N_1531_adj_5743[31]), 
          .S1(d7_71__N_1531_adj_5743[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_32 (.A0(d_d6_adj_5716[29]), .B0(d6_adj_5715[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[30]), .B1(d6_adj_5715[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16261), .COUT(n16262), .S0(d7_71__N_1531_adj_5743[29]), 
          .S1(d7_71__N_1531_adj_5743[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_32.INJECT1_1 = "NO";
    LUT4 i3169_4_lut_4_lut (.A(n18053), .B(n17817), .C(n250), .D(n244_adj_5062), 
         .Z(n2622)) /* synthesis lut_function=(A (C)+!A !(B+!(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3169_4_lut_4_lut.init = 16'hb1a0;
    LUT4 i2654_4_lut (.A(n275), .B(n2629), .C(n12538), .D(n17813), .Z(n12559)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2654_4_lut.init = 16'hafac;
    LUT4 mux_339_i7_4_lut (.A(n3945), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i7_4_lut.init = 16'hcfca;
    LUT4 mux_843_i6_3_lut (.A(n295_adj_5079), .B(n301), .C(led_c_4), .Z(n3945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i6_3_lut.init = 16'hcaca;
    LUT4 i2638_4_lut (.A(n311), .B(n2641), .C(n12538), .D(n17813), .Z(n12543)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2638_4_lut.init = 16'hafac;
    LUT4 i3266_4_lut (.A(n317), .B(n17822), .C(n2711), .D(n12538), .Z(n12540)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i3266_4_lut.init = 16'h2230;
    CCU2C _add_1_1478_add_4_30 (.A0(d_d6_adj_5716[27]), .B0(d6_adj_5715[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[28]), .B1(d6_adj_5715[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16260), .COUT(n16261), .S0(d7_71__N_1531_adj_5743[27]), 
          .S1(d7_71__N_1531_adj_5743[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_30.INJECT1_1 = "NO";
    LUT4 mux_339_i3_4_lut (.A(n3949), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2711)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i3_4_lut.init = 16'hcfca;
    LUT4 i3136_2_lut (.A(n313), .B(led_c_4), .Z(n3949)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i3136_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_76 (.A(led_c_1), .B(n16867), .C(led_c_3), .D(n17832), 
         .Z(n17022)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_76.init = 16'h0400;
    CCU2C _add_1_1478_add_4_28 (.A0(d_d6_adj_5716[25]), .B0(d6_adj_5715[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[26]), .B1(d6_adj_5715[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16259), .COUT(n16260), .S0(d7_71__N_1531_adj_5743[25]), 
          .S1(d7_71__N_1531_adj_5743[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_28.INJECT1_1 = "NO";
    CCU2C add_3665_19 (.A0(d_out_d_11__N_1886[17]), .B0(n48_adj_5593), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), .B1(n45_adj_5592), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16492), .S0(n45_adj_5682), 
          .S1(d_out_d_11__N_1888[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3665_19.INIT0 = 16'h9995;
    defparam add_3665_19.INIT1 = 16'h9995;
    defparam add_3665_19.INJECT1_0 = "NO";
    defparam add_3665_19.INJECT1_1 = "NO";
    CCU2C add_3665_17 (.A0(d_out_d_11__N_1886[17]), .B0(n54_adj_5595), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), .B1(n51_adj_5594), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16491), .COUT(n16492), .S0(n51_adj_5684), 
          .S1(n48_adj_5683));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3665_17.INIT0 = 16'h9995;
    defparam add_3665_17.INIT1 = 16'h9995;
    defparam add_3665_17.INJECT1_0 = "NO";
    defparam add_3665_17.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_26 (.A0(d_d6_adj_5716[23]), .B0(d6_adj_5715[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[24]), .B1(d6_adj_5715[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16258), .COUT(n16259), .S0(d7_71__N_1531_adj_5743[23]), 
          .S1(d7_71__N_1531_adj_5743[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_26.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(led_c_4), .B(led_c_5), .Z(n17073)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    CCU2C _add_1_1478_add_4_24 (.A0(d_d6_adj_5716[21]), .B0(d6_adj_5715[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[22]), .B1(d6_adj_5715[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16257), .COUT(n16258), .S0(d7_71__N_1531_adj_5743[21]), 
          .S1(d7_71__N_1531_adj_5743[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_22 (.A0(d_d6_adj_5716[19]), .B0(d6_adj_5715[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[20]), .B1(d6_adj_5715[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16256), .COUT(n16257), .S0(d7_71__N_1531_adj_5743[19]), 
          .S1(d7_71__N_1531_adj_5743[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_20 (.A0(d_d6_adj_5716[17]), .B0(d6_adj_5715[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[18]), .B1(d6_adj_5715[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16255), .COUT(n16256), .S0(d7_71__N_1531_adj_5743[17]), 
          .S1(d7_71__N_1531_adj_5743[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_10 (.A0(d5[43]), .B0(d4[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[44]), .B1(d4[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15422), .COUT(n15423), .S0(n162_adj_5313), .S1(n159_adj_5312));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_8 (.A0(d5[41]), .B0(d4[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[42]), .B1(d4[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15421), .COUT(n15422), .S0(n168_adj_5315), .S1(n165_adj_5314));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_6 (.A0(d5[39]), .B0(d4[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[40]), .B1(d4[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15420), .COUT(n15421), .S0(n174_adj_5317), .S1(n171_adj_5316));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_4 (.A0(d5[37]), .B0(d4[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[38]), .B1(d4[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15419), .COUT(n15420), .S0(n180_adj_5319), .S1(n177_adj_5318));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1538_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1538_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[36]), .B1(d4[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15419), .S1(n183_adj_5320));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1538_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1538_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1538_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1538_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_37 (.A0(d3_adj_5712[70]), .B0(cout_adj_5206), 
          .C0(n81_adj_5410), .D0(d4_adj_5713[70]), .A1(d3_adj_5712[71]), 
          .B1(cout_adj_5206), .C1(n78_adj_5409), .D1(d4_adj_5713[71]), 
          .CIN(n15417), .S0(d4_71__N_634_adj_5729[70]), .S1(d4_71__N_634_adj_5729[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_35 (.A0(d3_adj_5712[68]), .B0(cout_adj_5206), 
          .C0(n87_adj_5412), .D0(d4_adj_5713[68]), .A1(d3_adj_5712[69]), 
          .B1(cout_adj_5206), .C1(n84_adj_5411), .D1(d4_adj_5713[69]), 
          .CIN(n15416), .COUT(n15417), .S0(d4_71__N_634_adj_5729[68]), 
          .S1(d4_71__N_634_adj_5729[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_33 (.A0(d3_adj_5712[66]), .B0(cout_adj_5206), 
          .C0(n93_adj_5414), .D0(d4_adj_5713[66]), .A1(d3_adj_5712[67]), 
          .B1(cout_adj_5206), .C1(n90_adj_5413), .D1(d4_adj_5713[67]), 
          .CIN(n15415), .COUT(n15416), .S0(d4_71__N_634_adj_5729[66]), 
          .S1(d4_71__N_634_adj_5729[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_31 (.A0(d3_adj_5712[64]), .B0(cout_adj_5206), 
          .C0(n99_adj_5416), .D0(d4_adj_5713[64]), .A1(d3_adj_5712[65]), 
          .B1(cout_adj_5206), .C1(n96_adj_5415), .D1(d4_adj_5713[65]), 
          .CIN(n15414), .COUT(n15415), .S0(d4_71__N_634_adj_5729[64]), 
          .S1(d4_71__N_634_adj_5729[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_29 (.A0(d3_adj_5712[62]), .B0(cout_adj_5206), 
          .C0(n105_adj_5418), .D0(d4_adj_5713[62]), .A1(d3_adj_5712[63]), 
          .B1(cout_adj_5206), .C1(n102_adj_5417), .D1(d4_adj_5713[63]), 
          .CIN(n15413), .COUT(n15414), .S0(d4_71__N_634_adj_5729[62]), 
          .S1(d4_71__N_634_adj_5729[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_27 (.A0(d3_adj_5712[60]), .B0(cout_adj_5206), 
          .C0(n111_adj_5420), .D0(d4_adj_5713[60]), .A1(d3_adj_5712[61]), 
          .B1(cout_adj_5206), .C1(n108_adj_5419), .D1(d4_adj_5713[61]), 
          .CIN(n15412), .COUT(n15413), .S0(d4_71__N_634_adj_5729[60]), 
          .S1(d4_71__N_634_adj_5729[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_25 (.A0(d3_adj_5712[58]), .B0(cout_adj_5206), 
          .C0(n117_adj_5422), .D0(d4_adj_5713[58]), .A1(d3_adj_5712[59]), 
          .B1(cout_adj_5206), .C1(n114_adj_5421), .D1(d4_adj_5713[59]), 
          .CIN(n15411), .COUT(n15412), .S0(d4_71__N_634_adj_5729[58]), 
          .S1(d4_71__N_634_adj_5729[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_23 (.A0(d3_adj_5712[56]), .B0(cout_adj_5206), 
          .C0(n123_adj_5424), .D0(d4_adj_5713[56]), .A1(d3_adj_5712[57]), 
          .B1(cout_adj_5206), .C1(n120_adj_5423), .D1(d4_adj_5713[57]), 
          .CIN(n15410), .COUT(n15411), .S0(d4_71__N_634_adj_5729[56]), 
          .S1(d4_71__N_634_adj_5729[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_21 (.A0(d3_adj_5712[54]), .B0(cout_adj_5206), 
          .C0(n129_adj_5426), .D0(d4_adj_5713[54]), .A1(d3_adj_5712[55]), 
          .B1(cout_adj_5206), .C1(n126_adj_5425), .D1(d4_adj_5713[55]), 
          .CIN(n15409), .COUT(n15410), .S0(d4_71__N_634_adj_5729[54]), 
          .S1(d4_71__N_634_adj_5729[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_19 (.A0(d3_adj_5712[52]), .B0(cout_adj_5206), 
          .C0(n135_adj_5428), .D0(d4_adj_5713[52]), .A1(d3_adj_5712[53]), 
          .B1(cout_adj_5206), .C1(n132_adj_5427), .D1(d4_adj_5713[53]), 
          .CIN(n15408), .COUT(n15409), .S0(d4_71__N_634_adj_5729[52]), 
          .S1(d4_71__N_634_adj_5729[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_17 (.A0(d3_adj_5712[50]), .B0(cout_adj_5206), 
          .C0(n141_adj_5430), .D0(d4_adj_5713[50]), .A1(d3_adj_5712[51]), 
          .B1(cout_adj_5206), .C1(n138_adj_5429), .D1(d4_adj_5713[51]), 
          .CIN(n15407), .COUT(n15408), .S0(d4_71__N_634_adj_5729[50]), 
          .S1(d4_71__N_634_adj_5729[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_15 (.A0(d3_adj_5712[48]), .B0(cout_adj_5206), 
          .C0(n147_adj_5432), .D0(d4_adj_5713[48]), .A1(d3_adj_5712[49]), 
          .B1(cout_adj_5206), .C1(n144_adj_5431), .D1(d4_adj_5713[49]), 
          .CIN(n15406), .COUT(n15407), .S0(d4_71__N_634_adj_5729[48]), 
          .S1(d4_71__N_634_adj_5729[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_13 (.A0(d3_adj_5712[46]), .B0(cout_adj_5206), 
          .C0(n153_adj_5434), .D0(d4_adj_5713[46]), .A1(d3_adj_5712[47]), 
          .B1(cout_adj_5206), .C1(n150_adj_5433), .D1(d4_adj_5713[47]), 
          .CIN(n15405), .COUT(n15406), .S0(d4_71__N_634_adj_5729[46]), 
          .S1(d4_71__N_634_adj_5729[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_11 (.A0(d3_adj_5712[44]), .B0(cout_adj_5206), 
          .C0(n159_adj_5436), .D0(d4_adj_5713[44]), .A1(d3_adj_5712[45]), 
          .B1(cout_adj_5206), .C1(n156_adj_5435), .D1(d4_adj_5713[45]), 
          .CIN(n15404), .COUT(n15405), .S0(d4_71__N_634_adj_5729[44]), 
          .S1(d4_71__N_634_adj_5729[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_9 (.A0(d3_adj_5712[42]), .B0(cout_adj_5206), 
          .C0(n165_adj_5438), .D0(d4_adj_5713[42]), .A1(d3_adj_5712[43]), 
          .B1(cout_adj_5206), .C1(n162_adj_5437), .D1(d4_adj_5713[43]), 
          .CIN(n15403), .COUT(n15404), .S0(d4_71__N_634_adj_5729[42]), 
          .S1(d4_71__N_634_adj_5729[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_7 (.A0(d3_adj_5712[40]), .B0(cout_adj_5206), 
          .C0(n171_adj_5440), .D0(d4_adj_5713[40]), .A1(d3_adj_5712[41]), 
          .B1(cout_adj_5206), .C1(n168_adj_5439), .D1(d4_adj_5713[41]), 
          .CIN(n15402), .COUT(n15403), .S0(d4_71__N_634_adj_5729[40]), 
          .S1(d4_71__N_634_adj_5729[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_5 (.A0(d3_adj_5712[38]), .B0(cout_adj_5206), 
          .C0(n177_adj_5442), .D0(d4_adj_5713[38]), .A1(d3_adj_5712[39]), 
          .B1(cout_adj_5206), .C1(n174_adj_5441), .D1(d4_adj_5713[39]), 
          .CIN(n15401), .COUT(n15402), .S0(d4_71__N_634_adj_5729[38]), 
          .S1(d4_71__N_634_adj_5729[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_3 (.A0(d3_adj_5712[36]), .B0(cout_adj_5206), 
          .C0(n183_adj_5444), .D0(d4_adj_5713[36]), .A1(d3_adj_5712[37]), 
          .B1(cout_adj_5206), .C1(n180_adj_5443), .D1(d4_adj_5713[37]), 
          .CIN(n15400), .COUT(n15401), .S0(d4_71__N_634_adj_5729[36]), 
          .S1(d4_71__N_634_adj_5729[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1442_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1442_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5206), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15400));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1442_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1442_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1442_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_37 (.A0(d2_adj_5711[70]), .B0(cout_adj_4836), 
          .C0(n81_adj_5322), .D0(d3_adj_5712[70]), .A1(d2_adj_5711[71]), 
          .B1(cout_adj_4836), .C1(n78_adj_5321), .D1(d3_adj_5712[71]), 
          .CIN(n15393), .S0(d3_71__N_562_adj_5728[70]), .S1(d3_71__N_562_adj_5728[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_35 (.A0(d2_adj_5711[68]), .B0(cout_adj_4836), 
          .C0(n87_adj_5324), .D0(d3_adj_5712[68]), .A1(d2_adj_5711[69]), 
          .B1(cout_adj_4836), .C1(n84_adj_5323), .D1(d3_adj_5712[69]), 
          .CIN(n15392), .COUT(n15393), .S0(d3_71__N_562_adj_5728[68]), 
          .S1(d3_71__N_562_adj_5728[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_33 (.A0(d2_adj_5711[66]), .B0(cout_adj_4836), 
          .C0(n93_adj_5326), .D0(d3_adj_5712[66]), .A1(d2_adj_5711[67]), 
          .B1(cout_adj_4836), .C1(n90_adj_5325), .D1(d3_adj_5712[67]), 
          .CIN(n15391), .COUT(n15392), .S0(d3_71__N_562_adj_5728[66]), 
          .S1(d3_71__N_562_adj_5728[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_31 (.A0(d2_adj_5711[64]), .B0(cout_adj_4836), 
          .C0(n99_adj_5328), .D0(d3_adj_5712[64]), .A1(d2_adj_5711[65]), 
          .B1(cout_adj_4836), .C1(n96_adj_5327), .D1(d3_adj_5712[65]), 
          .CIN(n15390), .COUT(n15391), .S0(d3_71__N_562_adj_5728[64]), 
          .S1(d3_71__N_562_adj_5728[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_29 (.A0(d2_adj_5711[62]), .B0(cout_adj_4836), 
          .C0(n105_adj_5330), .D0(d3_adj_5712[62]), .A1(d2_adj_5711[63]), 
          .B1(cout_adj_4836), .C1(n102_adj_5329), .D1(d3_adj_5712[63]), 
          .CIN(n15389), .COUT(n15390), .S0(d3_71__N_562_adj_5728[62]), 
          .S1(d3_71__N_562_adj_5728[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_27 (.A0(d2_adj_5711[60]), .B0(cout_adj_4836), 
          .C0(n111_adj_5332), .D0(d3_adj_5712[60]), .A1(d2_adj_5711[61]), 
          .B1(cout_adj_4836), .C1(n108_adj_5331), .D1(d3_adj_5712[61]), 
          .CIN(n15388), .COUT(n15389), .S0(d3_71__N_562_adj_5728[60]), 
          .S1(d3_71__N_562_adj_5728[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_25 (.A0(d2_adj_5711[58]), .B0(cout_adj_4836), 
          .C0(n117_adj_5334), .D0(d3_adj_5712[58]), .A1(d2_adj_5711[59]), 
          .B1(cout_adj_4836), .C1(n114_adj_5333), .D1(d3_adj_5712[59]), 
          .CIN(n15387), .COUT(n15388), .S0(d3_71__N_562_adj_5728[58]), 
          .S1(d3_71__N_562_adj_5728[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_23 (.A0(d2_adj_5711[56]), .B0(cout_adj_4836), 
          .C0(n123_adj_5336), .D0(d3_adj_5712[56]), .A1(d2_adj_5711[57]), 
          .B1(cout_adj_4836), .C1(n120_adj_5335), .D1(d3_adj_5712[57]), 
          .CIN(n15386), .COUT(n15387), .S0(d3_71__N_562_adj_5728[56]), 
          .S1(d3_71__N_562_adj_5728[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_21 (.A0(d2_adj_5711[54]), .B0(cout_adj_4836), 
          .C0(n129_adj_5338), .D0(d3_adj_5712[54]), .A1(d2_adj_5711[55]), 
          .B1(cout_adj_4836), .C1(n126_adj_5337), .D1(d3_adj_5712[55]), 
          .CIN(n15385), .COUT(n15386), .S0(d3_71__N_562_adj_5728[54]), 
          .S1(d3_71__N_562_adj_5728[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_19 (.A0(d2_adj_5711[52]), .B0(cout_adj_4836), 
          .C0(n135_adj_5340), .D0(d3_adj_5712[52]), .A1(d2_adj_5711[53]), 
          .B1(cout_adj_4836), .C1(n132_adj_5339), .D1(d3_adj_5712[53]), 
          .CIN(n15384), .COUT(n15385), .S0(d3_71__N_562_adj_5728[52]), 
          .S1(d3_71__N_562_adj_5728[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_17 (.A0(d2_adj_5711[50]), .B0(cout_adj_4836), 
          .C0(n141_adj_5342), .D0(d3_adj_5712[50]), .A1(d2_adj_5711[51]), 
          .B1(cout_adj_4836), .C1(n138_adj_5341), .D1(d3_adj_5712[51]), 
          .CIN(n15383), .COUT(n15384), .S0(d3_71__N_562_adj_5728[50]), 
          .S1(d3_71__N_562_adj_5728[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_15 (.A0(d2_adj_5711[48]), .B0(cout_adj_4836), 
          .C0(n147_adj_5344), .D0(d3_adj_5712[48]), .A1(d2_adj_5711[49]), 
          .B1(cout_adj_4836), .C1(n144_adj_5343), .D1(d3_adj_5712[49]), 
          .CIN(n15382), .COUT(n15383), .S0(d3_71__N_562_adj_5728[48]), 
          .S1(d3_71__N_562_adj_5728[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_13 (.A0(d2_adj_5711[46]), .B0(cout_adj_4836), 
          .C0(n153_adj_5346), .D0(d3_adj_5712[46]), .A1(d2_adj_5711[47]), 
          .B1(cout_adj_4836), .C1(n150_adj_5345), .D1(d3_adj_5712[47]), 
          .CIN(n15381), .COUT(n15382), .S0(d3_71__N_562_adj_5728[46]), 
          .S1(d3_71__N_562_adj_5728[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_11 (.A0(d2_adj_5711[44]), .B0(cout_adj_4836), 
          .C0(n159_adj_5348), .D0(d3_adj_5712[44]), .A1(d2_adj_5711[45]), 
          .B1(cout_adj_4836), .C1(n156_adj_5347), .D1(d3_adj_5712[45]), 
          .CIN(n15380), .COUT(n15381), .S0(d3_71__N_562_adj_5728[44]), 
          .S1(d3_71__N_562_adj_5728[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_9 (.A0(d2_adj_5711[42]), .B0(cout_adj_4836), 
          .C0(n165_adj_5350), .D0(d3_adj_5712[42]), .A1(d2_adj_5711[43]), 
          .B1(cout_adj_4836), .C1(n162_adj_5349), .D1(d3_adj_5712[43]), 
          .CIN(n15379), .COUT(n15380), .S0(d3_71__N_562_adj_5728[42]), 
          .S1(d3_71__N_562_adj_5728[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_7 (.A0(d2_adj_5711[40]), .B0(cout_adj_4836), 
          .C0(n171_adj_5352), .D0(d3_adj_5712[40]), .A1(d2_adj_5711[41]), 
          .B1(cout_adj_4836), .C1(n168_adj_5351), .D1(d3_adj_5712[41]), 
          .CIN(n15378), .COUT(n15379), .S0(d3_71__N_562_adj_5728[40]), 
          .S1(d3_71__N_562_adj_5728[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_5 (.A0(d2_adj_5711[38]), .B0(cout_adj_4836), 
          .C0(n177_adj_5354), .D0(d3_adj_5712[38]), .A1(d2_adj_5711[39]), 
          .B1(cout_adj_4836), .C1(n174_adj_5353), .D1(d3_adj_5712[39]), 
          .CIN(n15377), .COUT(n15378), .S0(d3_71__N_562_adj_5728[38]), 
          .S1(d3_71__N_562_adj_5728[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_3 (.A0(d2_adj_5711[36]), .B0(cout_adj_4836), 
          .C0(n183_adj_5356), .D0(d3_adj_5712[36]), .A1(d2_adj_5711[37]), 
          .B1(cout_adj_4836), .C1(n180_adj_5355), .D1(d3_adj_5712[37]), 
          .CIN(n15376), .COUT(n15377), .S0(d3_71__N_562_adj_5728[36]), 
          .S1(d3_71__N_562_adj_5728[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1445_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1445_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1445_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_4836), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15376));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1445_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1445_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1445_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1445_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_38 (.A0(d3_adj_5712[71]), .B0(d2_adj_5711[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15372), .S0(n78_adj_5321));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1547_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_36 (.A0(d3_adj_5712[69]), .B0(d2_adj_5711[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[70]), .B1(d2_adj_5711[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15371), .COUT(n15372), .S0(n84_adj_5323), 
          .S1(n81_adj_5322));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_34 (.A0(d3_adj_5712[67]), .B0(d2_adj_5711[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[68]), .B1(d2_adj_5711[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15370), .COUT(n15371), .S0(n90_adj_5325), 
          .S1(n87_adj_5324));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_32 (.A0(d3_adj_5712[65]), .B0(d2_adj_5711[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[66]), .B1(d2_adj_5711[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15369), .COUT(n15370), .S0(n96_adj_5327), 
          .S1(n93_adj_5326));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_30 (.A0(d3_adj_5712[63]), .B0(d2_adj_5711[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[64]), .B1(d2_adj_5711[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15368), .COUT(n15369), .S0(n102_adj_5329), 
          .S1(n99_adj_5328));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_28 (.A0(d3_adj_5712[61]), .B0(d2_adj_5711[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[62]), .B1(d2_adj_5711[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15367), .COUT(n15368), .S0(n108_adj_5331), 
          .S1(n105_adj_5330));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_26 (.A0(d3_adj_5712[59]), .B0(d2_adj_5711[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[60]), .B1(d2_adj_5711[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15366), .COUT(n15367), .S0(n114_adj_5333), 
          .S1(n111_adj_5332));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_24 (.A0(d3_adj_5712[57]), .B0(d2_adj_5711[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[58]), .B1(d2_adj_5711[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15365), .COUT(n15366), .S0(n120_adj_5335), 
          .S1(n117_adj_5334));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_22 (.A0(d3_adj_5712[55]), .B0(d2_adj_5711[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[56]), .B1(d2_adj_5711[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15364), .COUT(n15365), .S0(n126_adj_5337), 
          .S1(n123_adj_5336));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_20 (.A0(d3_adj_5712[53]), .B0(d2_adj_5711[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[54]), .B1(d2_adj_5711[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15363), .COUT(n15364), .S0(n132_adj_5339), 
          .S1(n129_adj_5338));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_18 (.A0(d3_adj_5712[51]), .B0(d2_adj_5711[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[52]), .B1(d2_adj_5711[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15362), .COUT(n15363), .S0(n138_adj_5341), 
          .S1(n135_adj_5340));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_16 (.A0(d3_adj_5712[49]), .B0(d2_adj_5711[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[50]), .B1(d2_adj_5711[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15361), .COUT(n15362), .S0(n144_adj_5343), 
          .S1(n141_adj_5342));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_14 (.A0(d3_adj_5712[47]), .B0(d2_adj_5711[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[48]), .B1(d2_adj_5711[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15360), .COUT(n15361), .S0(n150_adj_5345), 
          .S1(n147_adj_5344));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_12 (.A0(d3_adj_5712[45]), .B0(d2_adj_5711[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[46]), .B1(d2_adj_5711[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15359), .COUT(n15360), .S0(n156_adj_5347), 
          .S1(n153_adj_5346));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_10 (.A0(d3_adj_5712[43]), .B0(d2_adj_5711[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[44]), .B1(d2_adj_5711[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15358), .COUT(n15359), .S0(n162_adj_5349), 
          .S1(n159_adj_5348));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_8 (.A0(d3_adj_5712[41]), .B0(d2_adj_5711[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[42]), .B1(d2_adj_5711[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15357), .COUT(n15358), .S0(n168_adj_5351), 
          .S1(n165_adj_5350));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_6 (.A0(d3_adj_5712[39]), .B0(d2_adj_5711[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[40]), .B1(d2_adj_5711[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15356), .COUT(n15357), .S0(n174_adj_5353), 
          .S1(n171_adj_5352));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_4 (.A0(d3_adj_5712[37]), .B0(d2_adj_5711[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5712[38]), .B1(d2_adj_5711[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15355), .COUT(n15356), .S0(n180_adj_5355), 
          .S1(n177_adj_5354));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1547_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1547_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d3_adj_5712[36]), .B1(d2_adj_5711[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15355), .S1(n183_adj_5356));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1547_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1547_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1547_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1547_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_37 (.A0(d1_adj_5710[70]), .B0(cout_adj_4835), 
          .C0(n81_adj_5609), .D0(d2_adj_5711[70]), .A1(d1_adj_5710[71]), 
          .B1(cout_adj_4835), .C1(n78_adj_5608), .D1(d2_adj_5711[71]), 
          .CIN(n15353), .S0(d2_71__N_490_adj_5727[70]), .S1(d2_71__N_490_adj_5727[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_35 (.A0(d1_adj_5710[68]), .B0(cout_adj_4835), 
          .C0(n87_adj_5611), .D0(d2_adj_5711[68]), .A1(d1_adj_5710[69]), 
          .B1(cout_adj_4835), .C1(n84_adj_5610), .D1(d2_adj_5711[69]), 
          .CIN(n15352), .COUT(n15353), .S0(d2_71__N_490_adj_5727[68]), 
          .S1(d2_71__N_490_adj_5727[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_33 (.A0(d1_adj_5710[66]), .B0(cout_adj_4835), 
          .C0(n93_adj_5613), .D0(d2_adj_5711[66]), .A1(d1_adj_5710[67]), 
          .B1(cout_adj_4835), .C1(n90_adj_5612), .D1(d2_adj_5711[67]), 
          .CIN(n15351), .COUT(n15352), .S0(d2_71__N_490_adj_5727[66]), 
          .S1(d2_71__N_490_adj_5727[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_31 (.A0(d1_adj_5710[64]), .B0(cout_adj_4835), 
          .C0(n99_adj_5615), .D0(d2_adj_5711[64]), .A1(d1_adj_5710[65]), 
          .B1(cout_adj_4835), .C1(n96_adj_5614), .D1(d2_adj_5711[65]), 
          .CIN(n15350), .COUT(n15351), .S0(d2_71__N_490_adj_5727[64]), 
          .S1(d2_71__N_490_adj_5727[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_29 (.A0(d1_adj_5710[62]), .B0(cout_adj_4835), 
          .C0(n105_adj_5617), .D0(d2_adj_5711[62]), .A1(d1_adj_5710[63]), 
          .B1(cout_adj_4835), .C1(n102_adj_5616), .D1(d2_adj_5711[63]), 
          .CIN(n15349), .COUT(n15350), .S0(d2_71__N_490_adj_5727[62]), 
          .S1(d2_71__N_490_adj_5727[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_27 (.A0(d1_adj_5710[60]), .B0(cout_adj_4835), 
          .C0(n111_adj_5619), .D0(d2_adj_5711[60]), .A1(d1_adj_5710[61]), 
          .B1(cout_adj_4835), .C1(n108_adj_5618), .D1(d2_adj_5711[61]), 
          .CIN(n15348), .COUT(n15349), .S0(d2_71__N_490_adj_5727[60]), 
          .S1(d2_71__N_490_adj_5727[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_25 (.A0(d1_adj_5710[58]), .B0(cout_adj_4835), 
          .C0(n117_adj_5621), .D0(d2_adj_5711[58]), .A1(d1_adj_5710[59]), 
          .B1(cout_adj_4835), .C1(n114_adj_5620), .D1(d2_adj_5711[59]), 
          .CIN(n15347), .COUT(n15348), .S0(d2_71__N_490_adj_5727[58]), 
          .S1(d2_71__N_490_adj_5727[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_23 (.A0(d1_adj_5710[56]), .B0(cout_adj_4835), 
          .C0(n123_adj_5623), .D0(d2_adj_5711[56]), .A1(d1_adj_5710[57]), 
          .B1(cout_adj_4835), .C1(n120_adj_5622), .D1(d2_adj_5711[57]), 
          .CIN(n15346), .COUT(n15347), .S0(d2_71__N_490_adj_5727[56]), 
          .S1(d2_71__N_490_adj_5727[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_21 (.A0(d1_adj_5710[54]), .B0(cout_adj_4835), 
          .C0(n129_adj_5625), .D0(d2_adj_5711[54]), .A1(d1_adj_5710[55]), 
          .B1(cout_adj_4835), .C1(n126_adj_5624), .D1(d2_adj_5711[55]), 
          .CIN(n15345), .COUT(n15346), .S0(d2_71__N_490_adj_5727[54]), 
          .S1(d2_71__N_490_adj_5727[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_19 (.A0(d1_adj_5710[52]), .B0(cout_adj_4835), 
          .C0(n135_adj_5627), .D0(d2_adj_5711[52]), .A1(d1_adj_5710[53]), 
          .B1(cout_adj_4835), .C1(n132_adj_5626), .D1(d2_adj_5711[53]), 
          .CIN(n15344), .COUT(n15345), .S0(d2_71__N_490_adj_5727[52]), 
          .S1(d2_71__N_490_adj_5727[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_17 (.A0(d1_adj_5710[50]), .B0(cout_adj_4835), 
          .C0(n141_adj_5629), .D0(d2_adj_5711[50]), .A1(d1_adj_5710[51]), 
          .B1(cout_adj_4835), .C1(n138_adj_5628), .D1(d2_adj_5711[51]), 
          .CIN(n15343), .COUT(n15344), .S0(d2_71__N_490_adj_5727[50]), 
          .S1(d2_71__N_490_adj_5727[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_15 (.A0(d1_adj_5710[48]), .B0(cout_adj_4835), 
          .C0(n147_adj_5631), .D0(d2_adj_5711[48]), .A1(d1_adj_5710[49]), 
          .B1(cout_adj_4835), .C1(n144_adj_5630), .D1(d2_adj_5711[49]), 
          .CIN(n15342), .COUT(n15343), .S0(d2_71__N_490_adj_5727[48]), 
          .S1(d2_71__N_490_adj_5727[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_13 (.A0(d1_adj_5710[46]), .B0(cout_adj_4835), 
          .C0(n153_adj_5633), .D0(d2_adj_5711[46]), .A1(d1_adj_5710[47]), 
          .B1(cout_adj_4835), .C1(n150_adj_5632), .D1(d2_adj_5711[47]), 
          .CIN(n15341), .COUT(n15342), .S0(d2_71__N_490_adj_5727[46]), 
          .S1(d2_71__N_490_adj_5727[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_11 (.A0(d1_adj_5710[44]), .B0(cout_adj_4835), 
          .C0(n159_adj_5635), .D0(d2_adj_5711[44]), .A1(d1_adj_5710[45]), 
          .B1(cout_adj_4835), .C1(n156_adj_5634), .D1(d2_adj_5711[45]), 
          .CIN(n15340), .COUT(n15341), .S0(d2_71__N_490_adj_5727[44]), 
          .S1(d2_71__N_490_adj_5727[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_9 (.A0(d1_adj_5710[42]), .B0(cout_adj_4835), 
          .C0(n165_adj_5637), .D0(d2_adj_5711[42]), .A1(d1_adj_5710[43]), 
          .B1(cout_adj_4835), .C1(n162_adj_5636), .D1(d2_adj_5711[43]), 
          .CIN(n15339), .COUT(n15340), .S0(d2_71__N_490_adj_5727[42]), 
          .S1(d2_71__N_490_adj_5727[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_7 (.A0(d1_adj_5710[40]), .B0(cout_adj_4835), 
          .C0(n171_adj_5639), .D0(d2_adj_5711[40]), .A1(d1_adj_5710[41]), 
          .B1(cout_adj_4835), .C1(n168_adj_5638), .D1(d2_adj_5711[41]), 
          .CIN(n15338), .COUT(n15339), .S0(d2_71__N_490_adj_5727[40]), 
          .S1(d2_71__N_490_adj_5727[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_5 (.A0(d1_adj_5710[38]), .B0(cout_adj_4835), 
          .C0(n177_adj_5641), .D0(d2_adj_5711[38]), .A1(d1_adj_5710[39]), 
          .B1(cout_adj_4835), .C1(n174_adj_5640), .D1(d2_adj_5711[39]), 
          .CIN(n15337), .COUT(n15338), .S0(d2_71__N_490_adj_5727[38]), 
          .S1(d2_71__N_490_adj_5727[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_3 (.A0(d1_adj_5710[36]), .B0(cout_adj_4835), 
          .C0(n183_adj_5643), .D0(d2_adj_5711[36]), .A1(d1_adj_5710[37]), 
          .B1(cout_adj_4835), .C1(n180_adj_5642), .D1(d2_adj_5711[37]), 
          .CIN(n15336), .COUT(n15337), .S0(d2_71__N_490_adj_5727[36]), 
          .S1(d2_71__N_490_adj_5727[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1448_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1448_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1448_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_4835), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15336));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1448_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1448_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1448_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1448_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_37 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n81_adj_5358), .D0(d1_adj_5710[70]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n78_adj_5357), .D1(d1_adj_5710[71]), 
          .CIN(n15331), .S0(d1_71__N_418_adj_5726[70]), .S1(d1_71__N_418_adj_5726[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_35 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n87_adj_5360), .D0(d1_adj_5710[68]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n84_adj_5359), .D1(d1_adj_5710[69]), 
          .CIN(n15330), .COUT(n15331), .S0(d1_71__N_418_adj_5726[68]), 
          .S1(d1_71__N_418_adj_5726[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_33 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n93_adj_5362), .D0(d1_adj_5710[66]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n90_adj_5361), .D1(d1_adj_5710[67]), 
          .CIN(n15329), .COUT(n15330), .S0(d1_71__N_418_adj_5726[66]), 
          .S1(d1_71__N_418_adj_5726[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_31 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n99_adj_5364), .D0(d1_adj_5710[64]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n96_adj_5363), .D1(d1_adj_5710[65]), 
          .CIN(n15328), .COUT(n15329), .S0(d1_71__N_418_adj_5726[64]), 
          .S1(d1_71__N_418_adj_5726[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_29 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n105_adj_5366), .D0(d1_adj_5710[62]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n102_adj_5365), .D1(d1_adj_5710[63]), 
          .CIN(n15327), .COUT(n15328), .S0(d1_71__N_418_adj_5726[62]), 
          .S1(d1_71__N_418_adj_5726[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_27 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n111_adj_5368), .D0(d1_adj_5710[60]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n108_adj_5367), .D1(d1_adj_5710[61]), 
          .CIN(n15326), .COUT(n15327), .S0(d1_71__N_418_adj_5726[60]), 
          .S1(d1_71__N_418_adj_5726[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_25 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n117_adj_5370), .D0(d1_adj_5710[58]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n114_adj_5369), .D1(d1_adj_5710[59]), 
          .CIN(n15325), .COUT(n15326), .S0(d1_71__N_418_adj_5726[58]), 
          .S1(d1_71__N_418_adj_5726[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_23 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n123_adj_5372), .D0(d1_adj_5710[56]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n120_adj_5371), .D1(d1_adj_5710[57]), 
          .CIN(n15324), .COUT(n15325), .S0(d1_71__N_418_adj_5726[56]), 
          .S1(d1_71__N_418_adj_5726[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_21 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n129_adj_5374), .D0(d1_adj_5710[54]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n126_adj_5373), .D1(d1_adj_5710[55]), 
          .CIN(n15323), .COUT(n15324), .S0(d1_71__N_418_adj_5726[54]), 
          .S1(d1_71__N_418_adj_5726[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_19 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n135_adj_5376), .D0(d1_adj_5710[52]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n132_adj_5375), .D1(d1_adj_5710[53]), 
          .CIN(n15322), .COUT(n15323), .S0(d1_71__N_418_adj_5726[52]), 
          .S1(d1_71__N_418_adj_5726[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_17 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n141_adj_5378), .D0(d1_adj_5710[50]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n138_adj_5377), .D1(d1_adj_5710[51]), 
          .CIN(n15321), .COUT(n15322), .S0(d1_71__N_418_adj_5726[50]), 
          .S1(d1_71__N_418_adj_5726[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_15 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n147_adj_5380), .D0(d1_adj_5710[48]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n144_adj_5379), .D1(d1_adj_5710[49]), 
          .CIN(n15320), .COUT(n15321), .S0(d1_71__N_418_adj_5726[48]), 
          .S1(d1_71__N_418_adj_5726[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_13 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n153_adj_5382), .D0(d1_adj_5710[46]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n150_adj_5381), .D1(d1_adj_5710[47]), 
          .CIN(n15319), .COUT(n15320), .S0(d1_71__N_418_adj_5726[46]), 
          .S1(d1_71__N_418_adj_5726[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_11 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n159_adj_5384), .D0(d1_adj_5710[44]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n156_adj_5383), .D1(d1_adj_5710[45]), 
          .CIN(n15318), .COUT(n15319), .S0(d1_71__N_418_adj_5726[44]), 
          .S1(d1_71__N_418_adj_5726[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_9 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n165_adj_5386), .D0(d1_adj_5710[42]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n162_adj_5385), .D1(d1_adj_5710[43]), 
          .CIN(n15317), .COUT(n15318), .S0(d1_71__N_418_adj_5726[42]), 
          .S1(d1_71__N_418_adj_5726[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_7 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n171_adj_5388), .D0(d1_adj_5710[40]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n168_adj_5387), .D1(d1_adj_5710[41]), 
          .CIN(n15316), .COUT(n15317), .S0(d1_71__N_418_adj_5726[40]), 
          .S1(d1_71__N_418_adj_5726[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_5 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n177_adj_5390), .D0(d1_adj_5710[38]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n174_adj_5389), .D1(d1_adj_5710[39]), 
          .CIN(n15315), .COUT(n15316), .S0(d1_71__N_418_adj_5726[38]), 
          .S1(d1_71__N_418_adj_5726[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_3 (.A0(MixerOutCos[11]), .B0(cout_adj_2809), 
          .C0(n183_adj_5392), .D0(d1_adj_5710[36]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_2809), .C1(n180_adj_5391), .D1(d1_adj_5710[37]), 
          .CIN(n15314), .COUT(n15315), .S0(d1_71__N_418_adj_5726[36]), 
          .S1(d1_71__N_418_adj_5726[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1451_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1451_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1451_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_2809), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15314));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1451_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1451_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1451_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1451_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_38 (.A0(d1_adj_5710[71]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15310), .S0(n78_adj_5357));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1541_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_36 (.A0(d1_adj_5710[69]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[70]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15309), .COUT(n15310), .S0(n84_adj_5359), 
          .S1(n81_adj_5358));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_34 (.A0(d1_adj_5710[67]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[68]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15308), .COUT(n15309), .S0(n90_adj_5361), 
          .S1(n87_adj_5360));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_32 (.A0(d1_adj_5710[65]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[66]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15307), .COUT(n15308), .S0(n96_adj_5363), 
          .S1(n93_adj_5362));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_30 (.A0(d1_adj_5710[63]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[64]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15306), .COUT(n15307), .S0(n102_adj_5365), 
          .S1(n99_adj_5364));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_28 (.A0(d1_adj_5710[61]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[62]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15305), .COUT(n15306), .S0(n108_adj_5367), 
          .S1(n105_adj_5366));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_26 (.A0(d1_adj_5710[59]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[60]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15304), .COUT(n15305), .S0(n114_adj_5369), 
          .S1(n111_adj_5368));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_24 (.A0(d1_adj_5710[57]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[58]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15303), .COUT(n15304), .S0(n120_adj_5371), 
          .S1(n117_adj_5370));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_22 (.A0(d1_adj_5710[55]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[56]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15302), .COUT(n15303), .S0(n126_adj_5373), 
          .S1(n123_adj_5372));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_20 (.A0(d1_adj_5710[53]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[54]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15301), .COUT(n15302), .S0(n132_adj_5375), 
          .S1(n129_adj_5374));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_18 (.A0(d1_adj_5710[51]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[52]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15300), .COUT(n15301), .S0(n138_adj_5377), 
          .S1(n135_adj_5376));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_16 (.A0(d1_adj_5710[49]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[50]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15299), .COUT(n15300), .S0(n144_adj_5379), 
          .S1(n141_adj_5378));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_14 (.A0(d1_adj_5710[47]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[48]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15298), .COUT(n15299), .S0(n150_adj_5381), 
          .S1(n147_adj_5380));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_12 (.A0(d1_adj_5710[45]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[46]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15297), .COUT(n15298), .S0(n156_adj_5383), 
          .S1(n153_adj_5382));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_10 (.A0(d1_adj_5710[43]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[44]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15296), .COUT(n15297), .S0(n162_adj_5385), 
          .S1(n159_adj_5384));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_8 (.A0(d1_adj_5710[41]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[42]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15295), .COUT(n15296), .S0(n168_adj_5387), 
          .S1(n165_adj_5386));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_6 (.A0(d1_adj_5710[39]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[40]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15294), .COUT(n15295), .S0(n174_adj_5389), 
          .S1(n171_adj_5388));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_4 (.A0(d1_adj_5710[37]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[38]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15293), .COUT(n15294), .S0(n180_adj_5391), 
          .S1(n177_adj_5390));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1541_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1541_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d1_adj_5710[36]), .B1(MixerOutCos[11]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15293), .S1(n183_adj_5392));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1541_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1541_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1541_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1541_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_37 (.A0(d1[70]), .B0(cout_adj_4558), .C0(n81_adj_5119), 
          .D0(d2[70]), .A1(d1[71]), .B1(cout_adj_4558), .C1(n78_adj_5118), 
          .D1(d2[71]), .CIN(n15291), .S0(d2_71__N_490[70]), .S1(d2_71__N_490[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_35 (.A0(d1[68]), .B0(cout_adj_4558), .C0(n87_adj_5121), 
          .D0(d2[68]), .A1(d1[69]), .B1(cout_adj_4558), .C1(n84_adj_5120), 
          .D1(d2[69]), .CIN(n15290), .COUT(n15291), .S0(d2_71__N_490[68]), 
          .S1(d2_71__N_490[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_33 (.A0(d1[66]), .B0(cout_adj_4558), .C0(n93_adj_5123), 
          .D0(d2[66]), .A1(d1[67]), .B1(cout_adj_4558), .C1(n90_adj_5122), 
          .D1(d2[67]), .CIN(n15289), .COUT(n15290), .S0(d2_71__N_490[66]), 
          .S1(d2_71__N_490[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_31 (.A0(d1[64]), .B0(cout_adj_4558), .C0(n99_adj_5125), 
          .D0(d2[64]), .A1(d1[65]), .B1(cout_adj_4558), .C1(n96_adj_5124), 
          .D1(d2[65]), .CIN(n15288), .COUT(n15289), .S0(d2_71__N_490[64]), 
          .S1(d2_71__N_490[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_29 (.A0(d1[62]), .B0(cout_adj_4558), .C0(n105_adj_5127), 
          .D0(d2[62]), .A1(d1[63]), .B1(cout_adj_4558), .C1(n102_adj_5126), 
          .D1(d2[63]), .CIN(n15287), .COUT(n15288), .S0(d2_71__N_490[62]), 
          .S1(d2_71__N_490[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_27 (.A0(d1[60]), .B0(cout_adj_4558), .C0(n111_adj_5129), 
          .D0(d2[60]), .A1(d1[61]), .B1(cout_adj_4558), .C1(n108_adj_5128), 
          .D1(d2[61]), .CIN(n15286), .COUT(n15287), .S0(d2_71__N_490[60]), 
          .S1(d2_71__N_490[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_25 (.A0(d1[58]), .B0(cout_adj_4558), .C0(n117_adj_5131), 
          .D0(d2[58]), .A1(d1[59]), .B1(cout_adj_4558), .C1(n114_adj_5130), 
          .D1(d2[59]), .CIN(n15285), .COUT(n15286), .S0(d2_71__N_490[58]), 
          .S1(d2_71__N_490[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_23 (.A0(d1[56]), .B0(cout_adj_4558), .C0(n123_adj_5133), 
          .D0(d2[56]), .A1(d1[57]), .B1(cout_adj_4558), .C1(n120_adj_5132), 
          .D1(d2[57]), .CIN(n15284), .COUT(n15285), .S0(d2_71__N_490[56]), 
          .S1(d2_71__N_490[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_21 (.A0(d1[54]), .B0(cout_adj_4558), .C0(n129_adj_5135), 
          .D0(d2[54]), .A1(d1[55]), .B1(cout_adj_4558), .C1(n126_adj_5134), 
          .D1(d2[55]), .CIN(n15283), .COUT(n15284), .S0(d2_71__N_490[54]), 
          .S1(d2_71__N_490[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_19 (.A0(d1[52]), .B0(cout_adj_4558), .C0(n135_adj_5137), 
          .D0(d2[52]), .A1(d1[53]), .B1(cout_adj_4558), .C1(n132_adj_5136), 
          .D1(d2[53]), .CIN(n15282), .COUT(n15283), .S0(d2_71__N_490[52]), 
          .S1(d2_71__N_490[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_17 (.A0(d1[50]), .B0(cout_adj_4558), .C0(n141_adj_5139), 
          .D0(d2[50]), .A1(d1[51]), .B1(cout_adj_4558), .C1(n138_adj_5138), 
          .D1(d2[51]), .CIN(n15281), .COUT(n15282), .S0(d2_71__N_490[50]), 
          .S1(d2_71__N_490[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_15 (.A0(d1[48]), .B0(cout_adj_4558), .C0(n147_adj_5141), 
          .D0(d2[48]), .A1(d1[49]), .B1(cout_adj_4558), .C1(n144_adj_5140), 
          .D1(d2[49]), .CIN(n15280), .COUT(n15281), .S0(d2_71__N_490[48]), 
          .S1(d2_71__N_490[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_13 (.A0(d1[46]), .B0(cout_adj_4558), .C0(n153_adj_5143), 
          .D0(d2[46]), .A1(d1[47]), .B1(cout_adj_4558), .C1(n150_adj_5142), 
          .D1(d2[47]), .CIN(n15279), .COUT(n15280), .S0(d2_71__N_490[46]), 
          .S1(d2_71__N_490[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_11 (.A0(d1[44]), .B0(cout_adj_4558), .C0(n159_adj_5145), 
          .D0(d2[44]), .A1(d1[45]), .B1(cout_adj_4558), .C1(n156_adj_5144), 
          .D1(d2[45]), .CIN(n15278), .COUT(n15279), .S0(d2_71__N_490[44]), 
          .S1(d2_71__N_490[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_9 (.A0(d1[42]), .B0(cout_adj_4558), .C0(n165_adj_5147), 
          .D0(d2[42]), .A1(d1[43]), .B1(cout_adj_4558), .C1(n162_adj_5146), 
          .D1(d2[43]), .CIN(n15277), .COUT(n15278), .S0(d2_71__N_490[42]), 
          .S1(d2_71__N_490[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_7 (.A0(d1[40]), .B0(cout_adj_4558), .C0(n171_adj_5149), 
          .D0(d2[40]), .A1(d1[41]), .B1(cout_adj_4558), .C1(n168_adj_5148), 
          .D1(d2[41]), .CIN(n15276), .COUT(n15277), .S0(d2_71__N_490[40]), 
          .S1(d2_71__N_490[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_5 (.A0(d1[38]), .B0(cout_adj_4558), .C0(n177_adj_5151), 
          .D0(d2[38]), .A1(d1[39]), .B1(cout_adj_4558), .C1(n174_adj_5150), 
          .D1(d2[39]), .CIN(n15275), .COUT(n15276), .S0(d2_71__N_490[38]), 
          .S1(d2_71__N_490[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_3 (.A0(d1[36]), .B0(cout_adj_4558), .C0(n183_adj_5153), 
          .D0(d2[36]), .A1(d1[37]), .B1(cout_adj_4558), .C1(n180_adj_5152), 
          .D1(d2[37]), .CIN(n15274), .COUT(n15275), .S0(d2_71__N_490[36]), 
          .S1(d2_71__N_490[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1463_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1463_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1463_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_4558), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15274));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1463_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1463_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1463_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1463_add_4_1.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_64 (.A0(phase_inc_carrGen1[62]), .B0(phase_accum[62]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[63]), .B1(phase_accum[63]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15269), .S0(n135_adj_5003), 
          .S1(n132_adj_5002));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_64.INIT0 = 16'h666a;
    defparam phase_accum_add_4_64.INIT1 = 16'h666a;
    defparam phase_accum_add_4_64.INJECT1_0 = "NO";
    defparam phase_accum_add_4_64.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_62 (.A0(phase_inc_carrGen1[60]), .B0(phase_accum[60]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[61]), .B1(phase_accum[61]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15268), .COUT(n15269), .S0(n141_adj_5005), 
          .S1(n138_adj_5004));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_62.INIT0 = 16'h666a;
    defparam phase_accum_add_4_62.INIT1 = 16'h666a;
    defparam phase_accum_add_4_62.INJECT1_0 = "NO";
    defparam phase_accum_add_4_62.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_60 (.A0(phase_inc_carrGen1[58]), .B0(phase_accum[58]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[59]), .B1(phase_accum[59]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15267), .COUT(n15268), .S0(n147_adj_5007), 
          .S1(n144_adj_5006));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_60.INIT0 = 16'h666a;
    defparam phase_accum_add_4_60.INIT1 = 16'h666a;
    defparam phase_accum_add_4_60.INJECT1_0 = "NO";
    defparam phase_accum_add_4_60.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_58 (.A0(phase_inc_carrGen1[56]), .B0(phase_accum[56]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[57]), .B1(phase_accum[57]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15266), .COUT(n15267), .S0(n153_adj_5009), 
          .S1(n150_adj_5008));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_58.INIT0 = 16'h666a;
    defparam phase_accum_add_4_58.INIT1 = 16'h666a;
    defparam phase_accum_add_4_58.INJECT1_0 = "NO";
    defparam phase_accum_add_4_58.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_56 (.A0(phase_inc_carrGen1[54]), .B0(phase_accum_adj_5702[54]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[55]), .B1(phase_accum_adj_5702[55]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15265), .COUT(n15266), .S0(n159_adj_5011), 
          .S1(n156_adj_5010));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_56.INIT0 = 16'h666a;
    defparam phase_accum_add_4_56.INIT1 = 16'h666a;
    defparam phase_accum_add_4_56.INJECT1_0 = "NO";
    defparam phase_accum_add_4_56.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_54 (.A0(phase_inc_carrGen1[52]), .B0(phase_accum_adj_5702[52]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[53]), .B1(phase_accum_adj_5702[53]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15264), .COUT(n15265), .S0(n165_adj_5013), 
          .S1(n162_adj_5012));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_54.INIT0 = 16'h666a;
    defparam phase_accum_add_4_54.INIT1 = 16'h666a;
    defparam phase_accum_add_4_54.INJECT1_0 = "NO";
    defparam phase_accum_add_4_54.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_52 (.A0(phase_inc_carrGen1[50]), .B0(phase_accum_adj_5702[50]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[51]), .B1(phase_accum_adj_5702[51]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15263), .COUT(n15264), .S0(n171_adj_5015), 
          .S1(n168_adj_5014));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_52.INIT0 = 16'h666a;
    defparam phase_accum_add_4_52.INIT1 = 16'h666a;
    defparam phase_accum_add_4_52.INJECT1_0 = "NO";
    defparam phase_accum_add_4_52.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_50 (.A0(phase_inc_carrGen1[48]), .B0(phase_accum_adj_5702[48]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[49]), .B1(phase_accum_adj_5702[49]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15262), .COUT(n15263), .S0(n177_adj_5017), 
          .S1(n174_adj_5016));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_50.INIT0 = 16'h666a;
    defparam phase_accum_add_4_50.INIT1 = 16'h666a;
    defparam phase_accum_add_4_50.INJECT1_0 = "NO";
    defparam phase_accum_add_4_50.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_48 (.A0(phase_inc_carrGen1[46]), .B0(phase_accum_adj_5702[46]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[47]), .B1(phase_accum_adj_5702[47]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15261), .COUT(n15262), .S0(n183_adj_5019), 
          .S1(n180_adj_5018));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_48.INIT0 = 16'h666a;
    defparam phase_accum_add_4_48.INIT1 = 16'h666a;
    defparam phase_accum_add_4_48.INJECT1_0 = "NO";
    defparam phase_accum_add_4_48.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_46 (.A0(phase_inc_carrGen1[44]), .B0(phase_accum_adj_5702[44]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[45]), .B1(phase_accum_adj_5702[45]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15260), .COUT(n15261), .S0(n189), 
          .S1(n186));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_46.INIT0 = 16'h666a;
    defparam phase_accum_add_4_46.INIT1 = 16'h666a;
    defparam phase_accum_add_4_46.INJECT1_0 = "NO";
    defparam phase_accum_add_4_46.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_44 (.A0(phase_inc_carrGen1[42]), .B0(phase_accum_adj_5702[42]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[43]), .B1(phase_accum_adj_5702[43]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15259), .COUT(n15260), .S0(n195), 
          .S1(n192));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_44.INIT0 = 16'h666a;
    defparam phase_accum_add_4_44.INIT1 = 16'h666a;
    defparam phase_accum_add_4_44.INJECT1_0 = "NO";
    defparam phase_accum_add_4_44.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_42 (.A0(phase_inc_carrGen1[40]), .B0(phase_accum_adj_5702[40]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[41]), .B1(phase_accum_adj_5702[41]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15258), .COUT(n15259), .S0(n201), 
          .S1(n198));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_42.INIT0 = 16'h666a;
    defparam phase_accum_add_4_42.INIT1 = 16'h666a;
    defparam phase_accum_add_4_42.INJECT1_0 = "NO";
    defparam phase_accum_add_4_42.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_40 (.A0(phase_inc_carrGen1[38]), .B0(phase_accum_adj_5702[38]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[39]), .B1(phase_accum_adj_5702[39]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15257), .COUT(n15258), .S0(n207), 
          .S1(n204));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_40.INIT0 = 16'h666a;
    defparam phase_accum_add_4_40.INIT1 = 16'h666a;
    defparam phase_accum_add_4_40.INJECT1_0 = "NO";
    defparam phase_accum_add_4_40.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_38 (.A0(phase_inc_carrGen1[36]), .B0(phase_accum_adj_5702[36]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[37]), .B1(phase_accum_adj_5702[37]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15256), .COUT(n15257), .S0(n213_adj_5020), 
          .S1(n210));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_38.INIT0 = 16'h666a;
    defparam phase_accum_add_4_38.INIT1 = 16'h666a;
    defparam phase_accum_add_4_38.INJECT1_0 = "NO";
    defparam phase_accum_add_4_38.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_36 (.A0(phase_inc_carrGen1[34]), .B0(phase_accum_adj_5702[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[35]), .B1(phase_accum_adj_5702[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15255), .COUT(n15256), .S0(n219), 
          .S1(n216));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_36.INIT0 = 16'h666a;
    defparam phase_accum_add_4_36.INIT1 = 16'h666a;
    defparam phase_accum_add_4_36.INJECT1_0 = "NO";
    defparam phase_accum_add_4_36.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_34 (.A0(phase_inc_carrGen1[32]), .B0(phase_accum_adj_5702[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[33]), .B1(phase_accum_adj_5702[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15254), .COUT(n15255), .S0(n225), 
          .S1(n222));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_34.INIT0 = 16'h666a;
    defparam phase_accum_add_4_34.INIT1 = 16'h666a;
    defparam phase_accum_add_4_34.INJECT1_0 = "NO";
    defparam phase_accum_add_4_34.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_32 (.A0(phase_inc_carrGen1[30]), .B0(phase_accum_adj_5702[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[31]), .B1(phase_accum_adj_5702[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15253), .COUT(n15254), .S0(n231), 
          .S1(n228));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_32.INIT0 = 16'h666a;
    defparam phase_accum_add_4_32.INIT1 = 16'h666a;
    defparam phase_accum_add_4_32.INJECT1_0 = "NO";
    defparam phase_accum_add_4_32.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_30 (.A0(phase_inc_carrGen1[28]), .B0(phase_accum_adj_5702[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[29]), .B1(phase_accum_adj_5702[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15252), .COUT(n15253), .S0(n237), 
          .S1(n234));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_30.INIT0 = 16'h666a;
    defparam phase_accum_add_4_30.INIT1 = 16'h666a;
    defparam phase_accum_add_4_30.INJECT1_0 = "NO";
    defparam phase_accum_add_4_30.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_28 (.A0(phase_inc_carrGen1[26]), .B0(phase_accum_adj_5702[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[27]), .B1(phase_accum_adj_5702[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15251), .COUT(n15252), .S0(n243), 
          .S1(n240));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_28.INIT0 = 16'h666a;
    defparam phase_accum_add_4_28.INIT1 = 16'h666a;
    defparam phase_accum_add_4_28.INJECT1_0 = "NO";
    defparam phase_accum_add_4_28.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_26 (.A0(phase_inc_carrGen1[24]), .B0(phase_accum_adj_5702[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[25]), .B1(phase_accum_adj_5702[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15250), .COUT(n15251), .S0(n249), 
          .S1(n246));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_26.INIT0 = 16'h666a;
    defparam phase_accum_add_4_26.INIT1 = 16'h666a;
    defparam phase_accum_add_4_26.INJECT1_0 = "NO";
    defparam phase_accum_add_4_26.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_24 (.A0(phase_inc_carrGen1[22]), .B0(phase_accum_adj_5702[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[23]), .B1(phase_accum_adj_5702[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15249), .COUT(n15250), .S0(n255), 
          .S1(n252));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_24.INIT0 = 16'h666a;
    defparam phase_accum_add_4_24.INIT1 = 16'h666a;
    defparam phase_accum_add_4_24.INJECT1_0 = "NO";
    defparam phase_accum_add_4_24.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_22 (.A0(phase_inc_carrGen1[20]), .B0(phase_accum_adj_5702[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[21]), .B1(phase_accum_adj_5702[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15248), .COUT(n15249), .S0(n261), 
          .S1(n258));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_22.INIT0 = 16'h666a;
    defparam phase_accum_add_4_22.INIT1 = 16'h666a;
    defparam phase_accum_add_4_22.INJECT1_0 = "NO";
    defparam phase_accum_add_4_22.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_20 (.A0(phase_inc_carrGen1[18]), .B0(phase_accum_adj_5702[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[19]), .B1(phase_accum_adj_5702[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15247), .COUT(n15248), .S0(n267), 
          .S1(n264));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_20.INIT0 = 16'h666a;
    defparam phase_accum_add_4_20.INIT1 = 16'h666a;
    defparam phase_accum_add_4_20.INJECT1_0 = "NO";
    defparam phase_accum_add_4_20.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_18 (.A0(phase_inc_carrGen1[16]), .B0(phase_accum_adj_5702[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[17]), .B1(phase_accum_adj_5702[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15246), .COUT(n15247), .S0(n273), 
          .S1(n270));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_18.INIT0 = 16'h666a;
    defparam phase_accum_add_4_18.INIT1 = 16'h666a;
    defparam phase_accum_add_4_18.INJECT1_0 = "NO";
    defparam phase_accum_add_4_18.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_16 (.A0(phase_inc_carrGen1[14]), .B0(phase_accum_adj_5702[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[15]), .B1(phase_accum_adj_5702[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15245), .COUT(n15246), .S0(n279), 
          .S1(n276));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_16.INIT0 = 16'h666a;
    defparam phase_accum_add_4_16.INIT1 = 16'h666a;
    defparam phase_accum_add_4_16.INJECT1_0 = "NO";
    defparam phase_accum_add_4_16.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_14 (.A0(phase_inc_carrGen1[12]), .B0(phase_accum_adj_5702[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[13]), .B1(phase_accum_adj_5702[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15244), .COUT(n15245), .S0(n285), 
          .S1(n282));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_14.INIT0 = 16'h666a;
    defparam phase_accum_add_4_14.INIT1 = 16'h666a;
    defparam phase_accum_add_4_14.INJECT1_0 = "NO";
    defparam phase_accum_add_4_14.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_12 (.A0(phase_inc_carrGen1[10]), .B0(phase_accum_adj_5702[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[11]), .B1(phase_accum_adj_5702[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15243), .COUT(n15244), .S0(n291), 
          .S1(n288));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_12.INIT0 = 16'h666a;
    defparam phase_accum_add_4_12.INIT1 = 16'h666a;
    defparam phase_accum_add_4_12.INJECT1_0 = "NO";
    defparam phase_accum_add_4_12.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_10 (.A0(phase_inc_carrGen1[8]), .B0(phase_accum_adj_5702[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[9]), .B1(phase_accum_adj_5702[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15242), .COUT(n15243), .S0(n297), 
          .S1(n294));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_10.INIT0 = 16'h666a;
    defparam phase_accum_add_4_10.INIT1 = 16'h666a;
    defparam phase_accum_add_4_10.INJECT1_0 = "NO";
    defparam phase_accum_add_4_10.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_8 (.A0(phase_inc_carrGen1[6]), .B0(phase_accum_adj_5702[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[7]), .B1(phase_accum_adj_5702[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15241), .COUT(n15242), .S0(n303), 
          .S1(n300));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_8.INIT0 = 16'h666a;
    defparam phase_accum_add_4_8.INIT1 = 16'h666a;
    defparam phase_accum_add_4_8.INJECT1_0 = "NO";
    defparam phase_accum_add_4_8.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_6 (.A0(phase_inc_carrGen1[4]), .B0(phase_accum_adj_5702[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[5]), .B1(phase_accum_adj_5702[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15240), .COUT(n15241), .S0(n309), 
          .S1(n306));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_6.INIT0 = 16'h666a;
    defparam phase_accum_add_4_6.INIT1 = 16'h666a;
    defparam phase_accum_add_4_6.INJECT1_0 = "NO";
    defparam phase_accum_add_4_6.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_4 (.A0(phase_inc_carrGen1[2]), .B0(phase_accum_adj_5702[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[3]), .B1(phase_accum_adj_5702[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15239), .COUT(n15240), .S0(n315), 
          .S1(n312));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_4.INIT0 = 16'h666a;
    defparam phase_accum_add_4_4.INIT1 = 16'h666a;
    defparam phase_accum_add_4_4.INJECT1_0 = "NO";
    defparam phase_accum_add_4_4.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_2 (.A0(phase_inc_carrGen1[0]), .B0(phase_accum_adj_5702[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[1]), .B1(phase_accum_adj_5702[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15239), .S1(n318));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_2.INIT0 = 16'h0008;
    defparam phase_accum_add_4_2.INIT1 = 16'h666a;
    defparam phase_accum_add_4_2.INJECT1_0 = "NO";
    defparam phase_accum_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15237), .S0(cout_adj_5021));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1604_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1604_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_36 (.A0(d1[34]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[35]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15236), .COUT(n15237), .S0(d1_71__N_418[34]), 
          .S1(d1_71__N_418[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_34 (.A0(d1[32]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[33]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15235), .COUT(n15236), .S0(d1_71__N_418[32]), 
          .S1(d1_71__N_418[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_32 (.A0(d1[30]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[31]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15234), .COUT(n15235), .S0(d1_71__N_418[30]), 
          .S1(d1_71__N_418[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_30 (.A0(d1[28]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[29]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15233), .COUT(n15234), .S0(d1_71__N_418[28]), 
          .S1(d1_71__N_418[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_28 (.A0(d1[26]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[27]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15232), .COUT(n15233), .S0(d1_71__N_418[26]), 
          .S1(d1_71__N_418[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_26 (.A0(d1[24]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[25]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15231), .COUT(n15232), .S0(d1_71__N_418[24]), 
          .S1(d1_71__N_418[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_24 (.A0(d1[22]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[23]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15230), .COUT(n15231), .S0(d1_71__N_418[22]), 
          .S1(d1_71__N_418[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_22 (.A0(d1[20]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[21]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15229), .COUT(n15230), .S0(d1_71__N_418[20]), 
          .S1(d1_71__N_418[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_20 (.A0(d1[18]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[19]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15228), .COUT(n15229), .S0(d1_71__N_418[18]), 
          .S1(d1_71__N_418[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_18 (.A0(d1[16]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[17]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15227), .COUT(n15228), .S0(d1_71__N_418[16]), 
          .S1(d1_71__N_418[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_16 (.A0(d1[14]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[15]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15226), .COUT(n15227), .S0(d1_71__N_418[14]), 
          .S1(d1_71__N_418[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_14 (.A0(d1[12]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[13]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15225), .COUT(n15226), .S0(d1_71__N_418[12]), 
          .S1(d1_71__N_418[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_12 (.A0(d1[10]), .B0(MixerOutSin[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[11]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15224), .COUT(n15225), .S0(d1_71__N_418[10]), 
          .S1(d1_71__N_418[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_10 (.A0(d1[8]), .B0(MixerOutSin[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[9]), .B1(MixerOutSin[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15223), .COUT(n15224), .S0(d1_71__N_418[8]), 
          .S1(d1_71__N_418[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_8 (.A0(d1[6]), .B0(MixerOutSin[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[7]), .B1(MixerOutSin[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15222), .COUT(n15223), .S0(d1_71__N_418[6]), 
          .S1(d1_71__N_418[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_6 (.A0(d1[4]), .B0(MixerOutSin[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[5]), .B1(MixerOutSin[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15221), .COUT(n15222), .S0(d1_71__N_418[4]), 
          .S1(d1_71__N_418[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_4 (.A0(d1[2]), .B0(MixerOutSin[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[3]), .B1(MixerOutSin[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15220), .COUT(n15221), .S0(d1_71__N_418[2]), 
          .S1(d1_71__N_418[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1604_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1604_add_4_2 (.A0(d1[0]), .B0(MixerOutSin[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[1]), .B1(MixerOutSin[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15220), .S1(d1_71__N_418[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1604_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1604_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1604_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1604_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_63 (.A0(phase_inc_carrGen[62]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[63]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15217), .S0(n133), .S1(n130));
    defparam _add_1_1607_add_4_63.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_63.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_63.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_63.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_61 (.A0(phase_inc_carrGen[60]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[61]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15216), .COUT(n15217), .S0(n139), 
          .S1(n136));
    defparam _add_1_1607_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_61.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_61.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_59 (.A0(phase_inc_carrGen[58]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[59]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15215), .COUT(n15216), .S0(n145), 
          .S1(n142));
    defparam _add_1_1607_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_57 (.A0(phase_inc_carrGen[56]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[57]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15214), .COUT(n15215), .S0(n151), 
          .S1(n148));
    defparam _add_1_1607_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_55 (.A0(phase_inc_carrGen[54]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[55]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15213), .COUT(n15214), .S0(n157), 
          .S1(n154));
    defparam _add_1_1607_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_53 (.A0(phase_inc_carrGen[52]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[53]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15212), .COUT(n15213), .S0(n163), 
          .S1(n160));
    defparam _add_1_1607_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_51 (.A0(phase_inc_carrGen[50]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[51]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15211), .COUT(n15212), .S0(n169), 
          .S1(n166));
    defparam _add_1_1607_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_49 (.A0(phase_inc_carrGen[48]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[49]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15210), .COUT(n15211), .S0(n175), 
          .S1(n172));
    defparam _add_1_1607_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_47 (.A0(phase_inc_carrGen[46]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[47]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15209), .COUT(n15210), .S0(n181), 
          .S1(n178));
    defparam _add_1_1607_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_1607_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_45 (.A0(phase_inc_carrGen[44]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[45]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15208), .COUT(n15209), .S0(n187), 
          .S1(n184));
    defparam _add_1_1607_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_45.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_43 (.A0(phase_inc_carrGen[42]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[43]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15207), .COUT(n15208), .S0(n193), 
          .S1(n190));
    defparam _add_1_1607_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_43.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_41 (.A0(phase_inc_carrGen[40]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[41]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15206), .COUT(n15207), .S0(n199), 
          .S1(n196));
    defparam _add_1_1607_add_4_41.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_39 (.A0(phase_inc_carrGen[38]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[39]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15205), .COUT(n15206), .S0(n205), 
          .S1(n202));
    defparam _add_1_1607_add_4_39.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_37 (.A0(phase_inc_carrGen[36]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[37]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15204), .COUT(n15205), .S0(n211), 
          .S1(n208));
    defparam _add_1_1607_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_35 (.A0(phase_inc_carrGen[34]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[35]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15203), .COUT(n15204), .S0(n217), 
          .S1(n214));
    defparam _add_1_1607_add_4_35.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_33 (.A0(phase_inc_carrGen[32]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[33]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15202), .COUT(n15203), .S0(n223), 
          .S1(n220));
    defparam _add_1_1607_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_31 (.A0(phase_inc_carrGen[30]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[31]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15201), .COUT(n15202), .S0(n229), 
          .S1(n226));
    defparam _add_1_1607_add_4_31.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_29 (.A0(phase_inc_carrGen[28]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[29]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15200), .COUT(n15201), .S0(n235), 
          .S1(n232));
    defparam _add_1_1607_add_4_29.INIT0 = 16'haaa0;
    defparam _add_1_1607_add_4_29.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_27 (.A0(phase_inc_carrGen[26]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[27]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15199), .COUT(n15200), .S0(n241), 
          .S1(n238));
    defparam _add_1_1607_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_25 (.A0(phase_inc_carrGen[24]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[25]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15198), .COUT(n15199), .S0(n247), 
          .S1(n244));
    defparam _add_1_1607_add_4_25.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_25.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_23 (.A0(phase_inc_carrGen[22]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[23]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15197), .COUT(n15198), .S0(n253), 
          .S1(n250));
    defparam _add_1_1607_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_21 (.A0(phase_inc_carrGen[20]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[21]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15196), .COUT(n15197), .S0(n259), 
          .S1(n256));
    defparam _add_1_1607_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_19 (.A0(phase_inc_carrGen[18]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[19]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15195), .COUT(n15196), .S0(n265), 
          .S1(n262));
    defparam _add_1_1607_add_4_19.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_17 (.A0(phase_inc_carrGen[16]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[17]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15194), .COUT(n15195), .S0(n271), 
          .S1(n268));
    defparam _add_1_1607_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1607_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_15 (.A0(phase_inc_carrGen[14]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[15]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15193), .COUT(n15194), .S0(n277), 
          .S1(n274));
    defparam _add_1_1607_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_13 (.A0(phase_inc_carrGen[12]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[13]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15192), .COUT(n15193), .S0(n283), 
          .S1(n280));
    defparam _add_1_1607_add_4_13.INIT0 = 16'h555f;
    defparam _add_1_1607_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_11 (.A0(phase_inc_carrGen[10]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[11]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15191), .COUT(n15192), .S0(n289), 
          .S1(n286));
    defparam _add_1_1607_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1607_add_4_11.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_9 (.A0(phase_inc_carrGen[8]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[9]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15190), .COUT(n15191), .S0(n295), 
          .S1(n292));
    defparam _add_1_1607_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1607_add_4_9.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_7 (.A0(phase_inc_carrGen[6]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[7]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15189), .COUT(n15190), .S0(n301), 
          .S1(n298));
    defparam _add_1_1607_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1607_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_5 (.A0(phase_inc_carrGen[4]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[5]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15188), .COUT(n15189), .S0(n307), 
          .S1(n304));
    defparam _add_1_1607_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1607_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_3 (.A0(phase_inc_carrGen[2]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[3]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15187), .COUT(n15188), .S0(n313), 
          .S1(n310));
    defparam _add_1_1607_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1607_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1607_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1607_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15187), .S1(n316));
    defparam _add_1_1607_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1607_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1607_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1607_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_61 (.A0(phase_inc_carrGen[63]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15186), .S0(n124));
    defparam _add_1_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_add_4_61.INIT1 = 16'h0000;
    defparam _add_1_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_add_4_61.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_59 (.A0(phase_inc_carrGen[61]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[62]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15185), .COUT(n15186), .S0(n130_adj_5024), 
          .S1(n127));
    defparam _add_1_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_57 (.A0(phase_inc_carrGen[59]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[60]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15184), .COUT(n15185), .S0(n136_adj_5026), 
          .S1(n133_adj_5025));
    defparam _add_1_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_55 (.A0(phase_inc_carrGen[57]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[58]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15183), .COUT(n15184), .S0(n142_adj_5028), 
          .S1(n139_adj_5027));
    defparam _add_1_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_53 (.A0(phase_inc_carrGen[55]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[56]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15182), .COUT(n15183), .S0(n148_adj_5030), 
          .S1(n145_adj_5029));
    defparam _add_1_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_51 (.A0(phase_inc_carrGen[53]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[54]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15181), .COUT(n15182), .S0(n154_adj_5032), 
          .S1(n151_adj_5031));
    defparam _add_1_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_49 (.A0(phase_inc_carrGen[51]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[52]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15180), .COUT(n15181), .S0(n160_adj_5034), 
          .S1(n157_adj_5033));
    defparam _add_1_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_47 (.A0(phase_inc_carrGen[49]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[50]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15179), .COUT(n15180), .S0(n166_adj_5036), 
          .S1(n163_adj_5035));
    defparam _add_1_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_45 (.A0(phase_inc_carrGen[47]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[48]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15178), .COUT(n15179), .S0(n172_adj_5038), 
          .S1(n169_adj_5037));
    defparam _add_1_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_add_4_45.INIT1 = 16'haaa0;
    defparam _add_1_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_43 (.A0(phase_inc_carrGen[45]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[46]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15177), .COUT(n15178), .S0(n178_adj_5040), 
          .S1(n175_adj_5039));
    defparam _add_1_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_add_4_43.INIT1 = 16'h555f;
    defparam _add_1_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_41 (.A0(phase_inc_carrGen[43]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[44]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15176), .COUT(n15177), .S0(n184_adj_5042), 
          .S1(n181_adj_5041));
    defparam _add_1_add_4_41.INIT0 = 16'haaa0;
    defparam _add_1_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_39 (.A0(phase_inc_carrGen[41]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[42]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15175), .COUT(n15176), .S0(n190_adj_5044), 
          .S1(n187_adj_5043));
    defparam _add_1_add_4_39.INIT0 = 16'haaa0;
    defparam _add_1_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_37 (.A0(phase_inc_carrGen[39]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[40]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15174), .COUT(n15175), .S0(n196_adj_5046), 
          .S1(n193_adj_5045));
    defparam _add_1_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_35 (.A0(phase_inc_carrGen[37]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[38]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15173), .COUT(n15174), .S0(n202_adj_5048), 
          .S1(n199_adj_5047));
    defparam _add_1_add_4_35.INIT0 = 16'haaa0;
    defparam _add_1_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_33 (.A0(phase_inc_carrGen[35]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[36]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15172), .COUT(n15173), .S0(n208_adj_5050), 
          .S1(n205_adj_5049));
    defparam _add_1_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_31 (.A0(phase_inc_carrGen[33]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[34]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15171), .COUT(n15172), .S0(n214_adj_5052), 
          .S1(n211_adj_5051));
    defparam _add_1_add_4_31.INIT0 = 16'haaa0;
    defparam _add_1_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_29 (.A0(phase_inc_carrGen[31]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[32]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15170), .COUT(n15171), .S0(n220_adj_5054), 
          .S1(n217_adj_5053));
    defparam _add_1_add_4_29.INIT0 = 16'h555f;
    defparam _add_1_add_4_29.INIT1 = 16'haaa0;
    defparam _add_1_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_27 (.A0(phase_inc_carrGen[29]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[30]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15169), .COUT(n15170), .S0(n226_adj_5056), 
          .S1(n223_adj_5055));
    defparam _add_1_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_25 (.A0(phase_inc_carrGen[27]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[28]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15168), .COUT(n15169), .S0(n232_adj_5058), 
          .S1(n229_adj_5057));
    defparam _add_1_add_4_25.INIT0 = 16'haaa0;
    defparam _add_1_add_4_25.INIT1 = 16'haaa0;
    defparam _add_1_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_23 (.A0(phase_inc_carrGen[25]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[26]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15167), .COUT(n15168), .S0(n238_adj_5060), 
          .S1(n235_adj_5059));
    defparam _add_1_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_21 (.A0(phase_inc_carrGen[23]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[24]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15166), .COUT(n15167), .S0(n244_adj_5062), 
          .S1(n241_adj_5061));
    defparam _add_1_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_19 (.A0(phase_inc_carrGen[21]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[22]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15165), .COUT(n15166), .S0(n250_adj_5064), 
          .S1(n247_adj_5063));
    defparam _add_1_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_17 (.A0(phase_inc_carrGen[19]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[20]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15164), .COUT(n15165), .S0(n256_adj_5066), 
          .S1(n253_adj_5065));
    defparam _add_1_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_add_4_17.INIT1 = 16'h555f;
    defparam _add_1_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_15 (.A0(phase_inc_carrGen[17]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[18]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15163), .COUT(n15164), .S0(n262_adj_5068), 
          .S1(n259_adj_5067));
    defparam _add_1_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_add_4_15.INIT1 = 16'h555f;
    defparam _add_1_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_13 (.A0(phase_inc_carrGen[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[16]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15162), .COUT(n15163), .S0(n268_adj_5070), 
          .S1(n265_adj_5069));
    defparam _add_1_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_add_4_13.INIT1 = 16'h555f;
    defparam _add_1_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_11 (.A0(phase_inc_carrGen[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15161), .COUT(n15162), .S0(n274_adj_5072), 
          .S1(n271_adj_5071));
    defparam _add_1_add_4_11.INIT0 = 16'h555f;
    defparam _add_1_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_9 (.A0(phase_inc_carrGen[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15160), .COUT(n15161), .S0(n280_adj_5074), 
          .S1(n277_adj_5073));
    defparam _add_1_add_4_9.INIT0 = 16'h555f;
    defparam _add_1_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_7 (.A0(phase_inc_carrGen[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15159), .COUT(n15160), .S0(n286_adj_5076), 
          .S1(n283_adj_5075));
    defparam _add_1_add_4_7.INIT0 = 16'h555f;
    defparam _add_1_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_5 (.A0(phase_inc_carrGen[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15158), .COUT(n15159), .S0(n292_adj_5078), 
          .S1(n289_adj_5077));
    defparam _add_1_add_4_5.INIT0 = 16'h555f;
    defparam _add_1_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_3 (.A0(phase_inc_carrGen[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_carrGen[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15157), .COUT(n15158), .S0(n298_adj_5080), 
          .S1(n295_adj_5079));
    defparam _add_1_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(phase_inc_carrGen[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15157), .S1(n301_adj_5081));
    defparam _add_1_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_38 (.A0(d1[71]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15156), .S0(n78_adj_5082));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1526_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_36 (.A0(d1[69]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[70]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15155), .COUT(n15156), .S0(n84_adj_5084), 
          .S1(n81_adj_5083));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_34 (.A0(d1[67]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[68]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15154), .COUT(n15155), .S0(n90_adj_5086), 
          .S1(n87_adj_5085));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_32 (.A0(d1[65]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[66]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15153), .COUT(n15154), .S0(n96_adj_5088), 
          .S1(n93_adj_5087));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_30 (.A0(d1[63]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[64]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15152), .COUT(n15153), .S0(n102_adj_5090), 
          .S1(n99_adj_5089));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_28 (.A0(d1[61]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[62]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15151), .COUT(n15152), .S0(n108_adj_5092), 
          .S1(n105_adj_5091));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_26 (.A0(d1[59]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[60]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15150), .COUT(n15151), .S0(n114_adj_5094), 
          .S1(n111_adj_5093));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_24 (.A0(d1[57]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[58]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15149), .COUT(n15150), .S0(n120_adj_5096), 
          .S1(n117_adj_5095));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_22 (.A0(d1[55]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[56]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15148), .COUT(n15149), .S0(n126_adj_5098), 
          .S1(n123_adj_5097));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_20 (.A0(d1[53]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[54]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15147), .COUT(n15148), .S0(n132_adj_5100), 
          .S1(n129_adj_5099));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_18 (.A0(d1[51]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[52]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15146), .COUT(n15147), .S0(n138_adj_5102), 
          .S1(n135_adj_5101));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_16 (.A0(d1[49]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[50]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15145), .COUT(n15146), .S0(n144_adj_5104), 
          .S1(n141_adj_5103));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_14 (.A0(d1[47]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[48]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15144), .COUT(n15145), .S0(n150_adj_5106), 
          .S1(n147_adj_5105));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_12 (.A0(d1[45]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[46]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15143), .COUT(n15144), .S0(n156_adj_5108), 
          .S1(n153_adj_5107));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_10 (.A0(d1[43]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[44]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15142), .COUT(n15143), .S0(n162_adj_5110), 
          .S1(n159_adj_5109));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_8 (.A0(d1[41]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[42]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15141), .COUT(n15142), .S0(n168_adj_5112), 
          .S1(n165_adj_5111));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_6 (.A0(d1[39]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[40]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15140), .COUT(n15141), .S0(n174_adj_5114), 
          .S1(n171_adj_5113));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_4 (.A0(d1[37]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[38]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15139), .COUT(n15140), .S0(n180_adj_5116), 
          .S1(n177_adj_5115));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1526_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1526_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[36]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15139), .S1(n183_adj_5117));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1526_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1526_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1526_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1526_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_38 (.A0(d_d9[71]), .B0(d9[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15138), .S0(n78_adj_4560));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1580_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_36 (.A0(d_d9[69]), .B0(d9[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[70]), .B1(d9[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15137), .COUT(n15138), .S0(n84), .S1(n81_adj_4559));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_34 (.A0(d_d9[67]), .B0(d9[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[68]), .B1(d9[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15136), .COUT(n15137), .S0(n90), .S1(n87));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_32 (.A0(d_d9[65]), .B0(d9[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[66]), .B1(d9[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15135), .COUT(n15136), .S0(n96), .S1(n93));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_30 (.A0(d_d9[63]), .B0(d9[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[64]), .B1(d9[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15134), .COUT(n15135), .S0(n102), .S1(n99));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_28 (.A0(d_d9[61]), .B0(d9[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[62]), .B1(d9[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15133), .COUT(n15134), .S0(n108), .S1(n105));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_26 (.A0(d_d9[59]), .B0(d9[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[60]), .B1(d9[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15132), .COUT(n15133), .S0(n114), .S1(n111));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_24 (.A0(d_d9[57]), .B0(d9[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[58]), .B1(d9[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15131), .COUT(n15132), .S0(n120), .S1(n117));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_22 (.A0(d_d9[55]), .B0(d9[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[56]), .B1(d9[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15130), .COUT(n15131));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_20 (.A0(d_d9[53]), .B0(d9[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[54]), .B1(d9[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15129), .COUT(n15130));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_18 (.A0(d_d9[51]), .B0(d9[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[52]), .B1(d9[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15128), .COUT(n15129));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_16 (.A0(d_d9[49]), .B0(d9[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[50]), .B1(d9[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15127), .COUT(n15128));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_14 (.A0(d_d9[47]), .B0(d9[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[48]), .B1(d9[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15126), .COUT(n15127));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_12 (.A0(d_d9[45]), .B0(d9[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[46]), .B1(d9[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15125), .COUT(n15126));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_10 (.A0(d_d9[43]), .B0(d9[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[44]), .B1(d9[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15124), .COUT(n15125));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_8 (.A0(d_d9[41]), .B0(d9[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[42]), .B1(d9[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15123), .COUT(n15124));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_6 (.A0(d_d9[39]), .B0(d9[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[40]), .B1(d9[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15122), .COUT(n15123));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_4 (.A0(d_d9[37]), .B0(d9[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[38]), .B1(d9[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15121), .COUT(n15122));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1580_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1580_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[36]), .B1(d9[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15121));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1580_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1580_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1580_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1580_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15120), .S0(cout_adj_4267));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1368_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1368_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_36 (.A0(d4[34]), .B0(d3[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[35]), .B1(d3[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15119), .COUT(n15120), .S0(d4_71__N_634[34]), .S1(d4_71__N_634[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_34 (.A0(d4[32]), .B0(d3[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[33]), .B1(d3[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15118), .COUT(n15119), .S0(d4_71__N_634[32]), .S1(d4_71__N_634[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_32 (.A0(d4[30]), .B0(d3[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[31]), .B1(d3[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15117), .COUT(n15118), .S0(d4_71__N_634[30]), .S1(d4_71__N_634[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_30 (.A0(d4[28]), .B0(d3[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[29]), .B1(d3[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15116), .COUT(n15117), .S0(d4_71__N_634[28]), .S1(d4_71__N_634[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_28 (.A0(d4[26]), .B0(d3[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[27]), .B1(d3[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15115), .COUT(n15116), .S0(d4_71__N_634[26]), .S1(d4_71__N_634[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_26 (.A0(d4[24]), .B0(d3[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[25]), .B1(d3[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15114), .COUT(n15115), .S0(d4_71__N_634[24]), .S1(d4_71__N_634[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_24 (.A0(d4[22]), .B0(d3[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[23]), .B1(d3[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15113), .COUT(n15114), .S0(d4_71__N_634[22]), .S1(d4_71__N_634[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_22 (.A0(d4[20]), .B0(d3[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[21]), .B1(d3[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15112), .COUT(n15113), .S0(d4_71__N_634[20]), .S1(d4_71__N_634[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_20 (.A0(d4[18]), .B0(d3[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[19]), .B1(d3[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15111), .COUT(n15112), .S0(d4_71__N_634[18]), .S1(d4_71__N_634[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_18 (.A0(d4[16]), .B0(d3[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[17]), .B1(d3[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15110), .COUT(n15111), .S0(d4_71__N_634[16]), .S1(d4_71__N_634[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_16 (.A0(d4[14]), .B0(d3[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[15]), .B1(d3[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15109), .COUT(n15110), .S0(d4_71__N_634[14]), .S1(d4_71__N_634[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_14 (.A0(d4[12]), .B0(d3[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[13]), .B1(d3[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15108), .COUT(n15109), .S0(d4_71__N_634[12]), .S1(d4_71__N_634[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_12 (.A0(d4[10]), .B0(d3[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[11]), .B1(d3[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15107), .COUT(n15108), .S0(d4_71__N_634[10]), .S1(d4_71__N_634[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_10 (.A0(d4[8]), .B0(d3[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[9]), .B1(d3[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15106), .COUT(n15107), .S0(d4_71__N_634[8]), .S1(d4_71__N_634[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_8 (.A0(d4[6]), .B0(d3[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[7]), .B1(d3[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15105), 
          .COUT(n15106), .S0(d4_71__N_634[6]), .S1(d4_71__N_634[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_6 (.A0(d4[4]), .B0(d3[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[5]), .B1(d3[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15104), 
          .COUT(n15105), .S0(d4_71__N_634[4]), .S1(d4_71__N_634[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_4 (.A0(d4[2]), .B0(d3[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[3]), .B1(d3[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15103), 
          .COUT(n15104), .S0(d4_71__N_634[2]), .S1(d4_71__N_634[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1368_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1368_add_4_2 (.A0(d4[0]), .B0(d3[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[1]), .B1(d3[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15103), 
          .S1(d4_71__N_634[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1368_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1368_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1368_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1368_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_38 (.A0(d_d_tmp_adj_5709[71]), .B0(d_tmp_adj_5708[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15101), .S0(n78_adj_4842));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1583_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_36 (.A0(d_d_tmp_adj_5709[69]), .B0(d_tmp_adj_5708[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[70]), .B1(d_tmp_adj_5708[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15100), .COUT(n15101), .S0(n84_adj_4844), 
          .S1(n81_adj_4843));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_34 (.A0(d_d_tmp_adj_5709[67]), .B0(d_tmp_adj_5708[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[68]), .B1(d_tmp_adj_5708[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15099), .COUT(n15100), .S0(n90_adj_4846), 
          .S1(n87_adj_4845));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_32 (.A0(d_d_tmp_adj_5709[65]), .B0(d_tmp_adj_5708[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[66]), .B1(d_tmp_adj_5708[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15098), .COUT(n15099), .S0(n96_adj_4848), 
          .S1(n93_adj_4847));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_30 (.A0(d_d_tmp_adj_5709[63]), .B0(d_tmp_adj_5708[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[64]), .B1(d_tmp_adj_5708[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15097), .COUT(n15098), .S0(n102_adj_4850), 
          .S1(n99_adj_4849));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_28 (.A0(d_d_tmp_adj_5709[61]), .B0(d_tmp_adj_5708[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[62]), .B1(d_tmp_adj_5708[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15096), .COUT(n15097), .S0(n108_adj_4852), 
          .S1(n105_adj_4851));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_26 (.A0(d_d_tmp_adj_5709[59]), .B0(d_tmp_adj_5708[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[60]), .B1(d_tmp_adj_5708[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15095), .COUT(n15096), .S0(n114_adj_4854), 
          .S1(n111_adj_4853));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_24 (.A0(d_d_tmp_adj_5709[57]), .B0(d_tmp_adj_5708[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[58]), .B1(d_tmp_adj_5708[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15094), .COUT(n15095), .S0(n120_adj_4856), 
          .S1(n117_adj_4855));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_22 (.A0(d_d_tmp_adj_5709[55]), .B0(d_tmp_adj_5708[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[56]), .B1(d_tmp_adj_5708[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15093), .COUT(n15094), .S0(n126_adj_4858), 
          .S1(n123_adj_4857));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_20 (.A0(d_d_tmp_adj_5709[53]), .B0(d_tmp_adj_5708[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[54]), .B1(d_tmp_adj_5708[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15092), .COUT(n15093), .S0(n132_adj_4860), 
          .S1(n129_adj_4859));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_18 (.A0(d_d_tmp_adj_5709[51]), .B0(d_tmp_adj_5708[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[52]), .B1(d_tmp_adj_5708[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15091), .COUT(n15092), .S0(n138_adj_4862), 
          .S1(n135_adj_4861));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_16 (.A0(d_d_tmp_adj_5709[49]), .B0(d_tmp_adj_5708[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[50]), .B1(d_tmp_adj_5708[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15090), .COUT(n15091), .S0(n144_adj_4864), 
          .S1(n141_adj_4863));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_14 (.A0(d_d_tmp_adj_5709[47]), .B0(d_tmp_adj_5708[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[48]), .B1(d_tmp_adj_5708[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15089), .COUT(n15090), .S0(n150_adj_4866), 
          .S1(n147_adj_4865));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_12 (.A0(d_d_tmp_adj_5709[45]), .B0(d_tmp_adj_5708[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[46]), .B1(d_tmp_adj_5708[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15088), .COUT(n15089), .S0(n156_adj_4868), 
          .S1(n153_adj_4867));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_10 (.A0(d_d_tmp_adj_5709[43]), .B0(d_tmp_adj_5708[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[44]), .B1(d_tmp_adj_5708[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15087), .COUT(n15088), .S0(n162_adj_4870), 
          .S1(n159_adj_4869));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_8 (.A0(d_d_tmp_adj_5709[41]), .B0(d_tmp_adj_5708[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[42]), .B1(d_tmp_adj_5708[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15086), .COUT(n15087), .S0(n168_adj_4872), 
          .S1(n165_adj_4871));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_6 (.A0(d_d_tmp_adj_5709[39]), .B0(d_tmp_adj_5708[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[40]), .B1(d_tmp_adj_5708[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15085), .COUT(n15086), .S0(n174_adj_4874), 
          .S1(n171_adj_4873));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_4 (.A0(d_d_tmp_adj_5709[37]), .B0(d_tmp_adj_5708[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5709[38]), .B1(d_tmp_adj_5708[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15084), .COUT(n15085), .S0(n180_adj_4876), 
          .S1(n177_adj_4875));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1583_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1583_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp_adj_5709[36]), .B1(d_tmp_adj_5708[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15084), .S1(n183_adj_4877));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1583_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1583_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1583_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1583_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15083), .S0(cout_adj_2810));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1371_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1371_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_36 (.A0(d5[34]), .B0(d4[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[35]), .B1(d4[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15082), .COUT(n15083), .S0(d5_71__N_706[34]), .S1(d5_71__N_706[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_34 (.A0(d5[32]), .B0(d4[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[33]), .B1(d4[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15081), .COUT(n15082), .S0(d5_71__N_706[32]), .S1(d5_71__N_706[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_32 (.A0(d5[30]), .B0(d4[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[31]), .B1(d4[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15080), .COUT(n15081), .S0(d5_71__N_706[30]), .S1(d5_71__N_706[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_30 (.A0(d5[28]), .B0(d4[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[29]), .B1(d4[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15079), .COUT(n15080), .S0(d5_71__N_706[28]), .S1(d5_71__N_706[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_28 (.A0(d5[26]), .B0(d4[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[27]), .B1(d4[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15078), .COUT(n15079), .S0(d5_71__N_706[26]), .S1(d5_71__N_706[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_26 (.A0(d5[24]), .B0(d4[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[25]), .B1(d4[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15077), .COUT(n15078), .S0(d5_71__N_706[24]), .S1(d5_71__N_706[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_24 (.A0(d5[22]), .B0(d4[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[23]), .B1(d4[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15076), .COUT(n15077), .S0(d5_71__N_706[22]), .S1(d5_71__N_706[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_22 (.A0(d5[20]), .B0(d4[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[21]), .B1(d4[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15075), .COUT(n15076), .S0(d5_71__N_706[20]), .S1(d5_71__N_706[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_20 (.A0(d5[18]), .B0(d4[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[19]), .B1(d4[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15074), .COUT(n15075), .S0(d5_71__N_706[18]), .S1(d5_71__N_706[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_18 (.A0(d5[16]), .B0(d4[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[17]), .B1(d4[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15073), .COUT(n15074), .S0(d5_71__N_706[16]), .S1(d5_71__N_706[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_16 (.A0(d5[14]), .B0(d4[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[15]), .B1(d4[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15072), .COUT(n15073), .S0(d5_71__N_706[14]), .S1(d5_71__N_706[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_14 (.A0(d5[12]), .B0(d4[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[13]), .B1(d4[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15071), .COUT(n15072), .S0(d5_71__N_706[12]), .S1(d5_71__N_706[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_12 (.A0(d5[10]), .B0(d4[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[11]), .B1(d4[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15070), .COUT(n15071), .S0(d5_71__N_706[10]), .S1(d5_71__N_706[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_10 (.A0(d5[8]), .B0(d4[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[9]), .B1(d4[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15069), .COUT(n15070), .S0(d5_71__N_706[8]), .S1(d5_71__N_706[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_8 (.A0(d5[6]), .B0(d4[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[7]), .B1(d4[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15068), 
          .COUT(n15069), .S0(d5_71__N_706[6]), .S1(d5_71__N_706[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_6 (.A0(d5[4]), .B0(d4[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[5]), .B1(d4[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15067), 
          .COUT(n15068), .S0(d5_71__N_706[4]), .S1(d5_71__N_706[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_4 (.A0(d5[2]), .B0(d4[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[3]), .B1(d4[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15066), 
          .COUT(n15067), .S0(d5_71__N_706[2]), .S1(d5_71__N_706[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1371_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1371_add_4_2 (.A0(d5[0]), .B0(d4[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[1]), .B1(d4[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15066), 
          .S1(d5_71__N_706[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1371_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1371_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1371_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1371_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_38 (.A0(d_d8[35]), .B0(d8[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15064), .S0(d9_71__N_1675[35]), .S1(cout_adj_5461));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1487_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_36 (.A0(d_d8[33]), .B0(d8[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[34]), .B1(d8[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15063), .COUT(n15064), .S0(d9_71__N_1675[33]), .S1(d9_71__N_1675[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_34 (.A0(d_d8[31]), .B0(d8[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[32]), .B1(d8[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15062), .COUT(n15063), .S0(d9_71__N_1675[31]), .S1(d9_71__N_1675[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_32 (.A0(d_d8[29]), .B0(d8[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[30]), .B1(d8[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15061), .COUT(n15062), .S0(d9_71__N_1675[29]), .S1(d9_71__N_1675[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_30 (.A0(d_d8[27]), .B0(d8[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[28]), .B1(d8[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15060), .COUT(n15061), .S0(d9_71__N_1675[27]), .S1(d9_71__N_1675[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_28 (.A0(d_d8[25]), .B0(d8[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[26]), .B1(d8[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15059), .COUT(n15060), .S0(d9_71__N_1675[25]), .S1(d9_71__N_1675[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_26 (.A0(d_d8[23]), .B0(d8[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[24]), .B1(d8[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15058), .COUT(n15059), .S0(d9_71__N_1675[23]), .S1(d9_71__N_1675[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_24 (.A0(d_d8[21]), .B0(d8[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[22]), .B1(d8[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15057), .COUT(n15058), .S0(d9_71__N_1675[21]), .S1(d9_71__N_1675[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_22 (.A0(d_d8[19]), .B0(d8[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[20]), .B1(d8[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15056), .COUT(n15057), .S0(d9_71__N_1675[19]), .S1(d9_71__N_1675[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_20 (.A0(d_d8[17]), .B0(d8[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[18]), .B1(d8[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15055), .COUT(n15056), .S0(d9_71__N_1675[17]), .S1(d9_71__N_1675[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_18 (.A0(d_d8[15]), .B0(d8[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[16]), .B1(d8[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15054), .COUT(n15055), .S0(d9_71__N_1675[15]), .S1(d9_71__N_1675[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_16 (.A0(d_d8[13]), .B0(d8[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[14]), .B1(d8[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15053), .COUT(n15054), .S0(d9_71__N_1675[13]), .S1(d9_71__N_1675[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_14 (.A0(d_d8[11]), .B0(d8[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[12]), .B1(d8[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15052), .COUT(n15053), .S0(d9_71__N_1675[11]), .S1(d9_71__N_1675[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_12 (.A0(d_d8[9]), .B0(d8[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[10]), .B1(d8[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15051), .COUT(n15052), .S0(d9_71__N_1675[9]), .S1(d9_71__N_1675[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_10 (.A0(d_d8[7]), .B0(d8[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[8]), .B1(d8[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15050), .COUT(n15051), .S0(d9_71__N_1675[7]), .S1(d9_71__N_1675[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_8 (.A0(d_d8[5]), .B0(d8[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[6]), .B1(d8[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15049), .COUT(n15050), .S0(d9_71__N_1675[5]), .S1(d9_71__N_1675[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_6 (.A0(d_d8[3]), .B0(d8[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[4]), .B1(d8[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15048), .COUT(n15049), .S0(d9_71__N_1675[3]), .S1(d9_71__N_1675[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_4 (.A0(d_d8[1]), .B0(d8[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[2]), .B1(d8[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15047), .COUT(n15048), .S0(d9_71__N_1675[1]), .S1(d9_71__N_1675[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1487_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1487_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[0]), .B1(d8[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15047), .S1(d9_71__N_1675[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1487_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1487_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1487_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1487_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_38 (.A0(d_d6_adj_5716[71]), .B0(d6_adj_5715[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15046), .S0(n78_adj_4878));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1586_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_36 (.A0(d_d6_adj_5716[69]), .B0(d6_adj_5715[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[70]), .B1(d6_adj_5715[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15045), .COUT(n15046), .S0(n84_adj_4880), 
          .S1(n81_adj_4879));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_34 (.A0(d_d6_adj_5716[67]), .B0(d6_adj_5715[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[68]), .B1(d6_adj_5715[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15044), .COUT(n15045), .S0(n90_adj_4882), 
          .S1(n87_adj_4881));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_32 (.A0(d_d6_adj_5716[65]), .B0(d6_adj_5715[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[66]), .B1(d6_adj_5715[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15043), .COUT(n15044), .S0(n96_adj_4884), 
          .S1(n93_adj_4883));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_30 (.A0(d_d6_adj_5716[63]), .B0(d6_adj_5715[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[64]), .B1(d6_adj_5715[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15042), .COUT(n15043), .S0(n102_adj_4886), 
          .S1(n99_adj_4885));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_28 (.A0(d_d6_adj_5716[61]), .B0(d6_adj_5715[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[62]), .B1(d6_adj_5715[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15041), .COUT(n15042), .S0(n108_adj_4888), 
          .S1(n105_adj_4887));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_26 (.A0(d_d6_adj_5716[59]), .B0(d6_adj_5715[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[60]), .B1(d6_adj_5715[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15040), .COUT(n15041), .S0(n114_adj_4890), 
          .S1(n111_adj_4889));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_24 (.A0(d_d6_adj_5716[57]), .B0(d6_adj_5715[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[58]), .B1(d6_adj_5715[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15039), .COUT(n15040), .S0(n120_adj_4892), 
          .S1(n117_adj_4891));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_22 (.A0(d_d6_adj_5716[55]), .B0(d6_adj_5715[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[56]), .B1(d6_adj_5715[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15038), .COUT(n15039), .S0(n126_adj_4894), 
          .S1(n123_adj_4893));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_20 (.A0(d_d6_adj_5716[53]), .B0(d6_adj_5715[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[54]), .B1(d6_adj_5715[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15037), .COUT(n15038), .S0(n132_adj_4896), 
          .S1(n129_adj_4895));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_18 (.A0(d_d6_adj_5716[51]), .B0(d6_adj_5715[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[52]), .B1(d6_adj_5715[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15036), .COUT(n15037), .S0(n138_adj_4898), 
          .S1(n135_adj_4897));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_16 (.A0(d_d6_adj_5716[49]), .B0(d6_adj_5715[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[50]), .B1(d6_adj_5715[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15035), .COUT(n15036), .S0(n144_adj_4900), 
          .S1(n141_adj_4899));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_14 (.A0(d_d6_adj_5716[47]), .B0(d6_adj_5715[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[48]), .B1(d6_adj_5715[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15034), .COUT(n15035), .S0(n150_adj_4902), 
          .S1(n147_adj_4901));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_12 (.A0(d_d6_adj_5716[45]), .B0(d6_adj_5715[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[46]), .B1(d6_adj_5715[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15033), .COUT(n15034), .S0(n156_adj_4904), 
          .S1(n153_adj_4903));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_10 (.A0(d_d6_adj_5716[43]), .B0(d6_adj_5715[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[44]), .B1(d6_adj_5715[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15032), .COUT(n15033), .S0(n162_adj_4906), 
          .S1(n159_adj_4905));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_8 (.A0(d_d6_adj_5716[41]), .B0(d6_adj_5715[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[42]), .B1(d6_adj_5715[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15031), .COUT(n15032), .S0(n168_adj_4908), 
          .S1(n165_adj_4907));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_6 (.A0(d_d6_adj_5716[39]), .B0(d6_adj_5715[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[40]), .B1(d6_adj_5715[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15030), .COUT(n15031), .S0(n174_adj_4910), 
          .S1(n171_adj_4909));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_4 (.A0(d_d6_adj_5716[37]), .B0(d6_adj_5715[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[38]), .B1(d6_adj_5715[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15029), .COUT(n15030), .S0(n180_adj_4912), 
          .S1(n177_adj_4911));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1586_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1586_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6_adj_5716[36]), .B1(d6_adj_5715[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15029), .S1(n183_adj_4913));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1586_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1586_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1586_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1586_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_38 (.A0(d_d7_adj_5718[71]), .B0(d7_adj_5717[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15028), .S0(n78_adj_4914));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1589_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_36 (.A0(d_d7_adj_5718[69]), .B0(d7_adj_5717[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[70]), .B1(d7_adj_5717[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15027), .COUT(n15028), .S0(n84_adj_4916), 
          .S1(n81_adj_4915));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_34 (.A0(d_d7_adj_5718[67]), .B0(d7_adj_5717[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[68]), .B1(d7_adj_5717[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15026), .COUT(n15027), .S0(n90_adj_4918), 
          .S1(n87_adj_4917));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_32 (.A0(d_d7_adj_5718[65]), .B0(d7_adj_5717[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[66]), .B1(d7_adj_5717[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15025), .COUT(n15026), .S0(n96_adj_4920), 
          .S1(n93_adj_4919));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_30 (.A0(d_d7_adj_5718[63]), .B0(d7_adj_5717[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[64]), .B1(d7_adj_5717[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15024), .COUT(n15025), .S0(n102_adj_4922), 
          .S1(n99_adj_4921));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_28 (.A0(d_d7_adj_5718[61]), .B0(d7_adj_5717[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[62]), .B1(d7_adj_5717[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15023), .COUT(n15024), .S0(n108_adj_4924), 
          .S1(n105_adj_4923));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_26 (.A0(d_d7_adj_5718[59]), .B0(d7_adj_5717[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[60]), .B1(d7_adj_5717[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15022), .COUT(n15023), .S0(n114_adj_4926), 
          .S1(n111_adj_4925));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_24 (.A0(d_d7_adj_5718[57]), .B0(d7_adj_5717[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[58]), .B1(d7_adj_5717[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15021), .COUT(n15022), .S0(n120_adj_4928), 
          .S1(n117_adj_4927));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_22 (.A0(d_d7_adj_5718[55]), .B0(d7_adj_5717[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[56]), .B1(d7_adj_5717[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15020), .COUT(n15021), .S0(n126_adj_4930), 
          .S1(n123_adj_4929));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_20 (.A0(d_d7_adj_5718[53]), .B0(d7_adj_5717[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[54]), .B1(d7_adj_5717[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15019), .COUT(n15020), .S0(n132_adj_4932), 
          .S1(n129_adj_4931));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_18 (.A0(d_d7_adj_5718[51]), .B0(d7_adj_5717[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[52]), .B1(d7_adj_5717[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15018), .COUT(n15019), .S0(n138_adj_4934), 
          .S1(n135_adj_4933));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_16 (.A0(d_d7_adj_5718[49]), .B0(d7_adj_5717[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[50]), .B1(d7_adj_5717[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15017), .COUT(n15018), .S0(n144_adj_4936), 
          .S1(n141_adj_4935));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_14 (.A0(d_d7_adj_5718[47]), .B0(d7_adj_5717[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[48]), .B1(d7_adj_5717[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15016), .COUT(n15017), .S0(n150_adj_4938), 
          .S1(n147_adj_4937));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_12 (.A0(d_d7_adj_5718[45]), .B0(d7_adj_5717[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[46]), .B1(d7_adj_5717[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15015), .COUT(n15016), .S0(n156_adj_4940), 
          .S1(n153_adj_4939));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_10 (.A0(d_d7_adj_5718[43]), .B0(d7_adj_5717[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[44]), .B1(d7_adj_5717[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15014), .COUT(n15015), .S0(n162_adj_4942), 
          .S1(n159_adj_4941));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_8 (.A0(d_d7_adj_5718[41]), .B0(d7_adj_5717[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[42]), .B1(d7_adj_5717[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15013), .COUT(n15014), .S0(n168_adj_4944), 
          .S1(n165_adj_4943));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_6 (.A0(d_d7_adj_5718[39]), .B0(d7_adj_5717[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[40]), .B1(d7_adj_5717[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15012), .COUT(n15013), .S0(n174_adj_4946), 
          .S1(n171_adj_4945));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_4 (.A0(d_d7_adj_5718[37]), .B0(d7_adj_5717[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[38]), .B1(d7_adj_5717[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15011), .COUT(n15012), .S0(n180_adj_4948), 
          .S1(n177_adj_4947));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1589_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1589_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7_adj_5718[36]), .B1(d7_adj_5717[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15011), .S1(n183_adj_4949));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1589_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1589_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1589_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1589_add_4_2.INJECT1_1 = "NO";
    FD1S3AX ISquare_e3__i2 (.D(n123_adj_5247), .CK(CIC1_out_clkSin), .Q(ISquare[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i2.GSR = "ENABLED";
    CCU2C _add_1_1374_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15010), .S0(cout_adj_2809));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1374_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1374_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_36 (.A0(d1_adj_5710[34]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[35]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15009), .COUT(n15010), .S0(d1_71__N_418_adj_5726[34]), 
          .S1(d1_71__N_418_adj_5726[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_34 (.A0(d1_adj_5710[32]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[33]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15008), .COUT(n15009), .S0(d1_71__N_418_adj_5726[32]), 
          .S1(d1_71__N_418_adj_5726[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_32 (.A0(d1_adj_5710[30]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[31]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15007), .COUT(n15008), .S0(d1_71__N_418_adj_5726[30]), 
          .S1(d1_71__N_418_adj_5726[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_30 (.A0(d1_adj_5710[28]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[29]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15006), .COUT(n15007), .S0(d1_71__N_418_adj_5726[28]), 
          .S1(d1_71__N_418_adj_5726[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_28 (.A0(d1_adj_5710[26]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[27]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15005), .COUT(n15006), .S0(d1_71__N_418_adj_5726[26]), 
          .S1(d1_71__N_418_adj_5726[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_26 (.A0(d1_adj_5710[24]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[25]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15004), .COUT(n15005), .S0(d1_71__N_418_adj_5726[24]), 
          .S1(d1_71__N_418_adj_5726[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_24 (.A0(d1_adj_5710[22]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[23]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15003), .COUT(n15004), .S0(d1_71__N_418_adj_5726[22]), 
          .S1(d1_71__N_418_adj_5726[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_22 (.A0(d1_adj_5710[20]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[21]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15002), .COUT(n15003), .S0(d1_71__N_418_adj_5726[20]), 
          .S1(d1_71__N_418_adj_5726[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_20 (.A0(d1_adj_5710[18]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[19]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15001), .COUT(n15002), .S0(d1_71__N_418_adj_5726[18]), 
          .S1(d1_71__N_418_adj_5726[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_12 (.A0(d1_adj_5710[10]), .B0(MixerOutCos[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[11]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14997), .COUT(n14998), .S0(d1_71__N_418_adj_5726[10]), 
          .S1(d1_71__N_418_adj_5726[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_12.INJECT1_1 = "NO";
    LUT4 i2799_2_lut (.A(n18096), .B(led_c_7), .Z(n12710)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i2799_2_lut.init = 16'h8888;
    CCU2C _add_1_1374_add_4_18 (.A0(d1_adj_5710[16]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[17]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15000), .COUT(n15001), .S0(d1_71__N_418_adj_5726[16]), 
          .S1(d1_71__N_418_adj_5726[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_8 (.A0(d1_adj_5710[6]), .B0(MixerOutCos[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[7]), .B1(MixerOutCos[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14995), .COUT(n14996), .S0(d1_71__N_418_adj_5726[6]), 
          .S1(d1_71__N_418_adj_5726[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_16 (.A0(d1_adj_5710[14]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[15]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14999), .COUT(n15000), .S0(d1_71__N_418_adj_5726[14]), 
          .S1(d1_71__N_418_adj_5726[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_6 (.A0(d1_adj_5710[4]), .B0(MixerOutCos[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[5]), .B1(MixerOutCos[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14994), .COUT(n14995), .S0(d1_71__N_418_adj_5726[4]), 
          .S1(d1_71__N_418_adj_5726[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1374_add_4_4 (.A0(d1_adj_5710[2]), .B0(MixerOutCos[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[3]), .B1(MixerOutCos[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14993), .COUT(n14994), .S0(d1_71__N_418_adj_5726[2]), 
          .S1(d1_71__N_418_adj_5726[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_4.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut (.A(n17809), .B(n17815), .C(n18096), .D(n17812), 
         .Z(clk_80mhz_enable_23)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf0b0;
    CCU2C _add_1_1374_add_4_10 (.A0(d1_adj_5710[8]), .B0(MixerOutCos[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[9]), .B1(MixerOutCos[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14996), .COUT(n14997), .S0(d1_71__N_418_adj_5726[8]), 
          .S1(d1_71__N_418_adj_5726[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_10.INJECT1_1 = "NO";
    LUT4 i1_3_lut (.A(led_c_3), .B(led_c_2), .C(led_c_6), .Z(n16829)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut.init = 16'hfefe;
    CCU2C _add_1_1374_add_4_14 (.A0(d1_adj_5710[12]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[13]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14998), .COUT(n14999), .S0(d1_71__N_418_adj_5726[12]), 
          .S1(d1_71__N_418_adj_5726[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1374_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_14.INJECT1_1 = "NO";
    CCU2C add_3665_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1886[17]), .C0(n60_adj_5597), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1886[17]), 
          .C1(n57_adj_5596), .D1(VCC_net), .CIN(n16490), .COUT(n16491), 
          .S0(n57_adj_5686), .S1(n54_adj_5685));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3665_15.INIT0 = 16'h6969;
    defparam add_3665_15.INIT1 = 16'h6969;
    defparam add_3665_15.INJECT1_0 = "NO";
    defparam add_3665_15.INJECT1_1 = "NO";
    CCU2C add_3665_13 (.A0(d_out_d_11__N_1886[17]), .B0(n66_adj_5599), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1886[17]), 
          .C1(n63_adj_5598), .D1(VCC_net), .CIN(n16489), .COUT(n16490), 
          .S0(n63_adj_5688), .S1(n60_adj_5687));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3665_13.INIT0 = 16'h9995;
    defparam add_3665_13.INIT1 = 16'h6969;
    defparam add_3665_13.INJECT1_0 = "NO";
    defparam add_3665_13.INJECT1_1 = "NO";
    CCU2C add_3665_11 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(n72_adj_5601), .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), 
          .B1(n17826), .C1(n69_adj_5600), .D1(VCC_net), .CIN(n16488), 
          .COUT(n16489), .S0(n69_adj_5690), .S1(n66_adj_5689));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3665_11.INIT0 = 16'h9696;
    defparam add_3665_11.INIT1 = 16'h6969;
    defparam add_3665_11.INJECT1_0 = "NO";
    defparam add_3665_11.INJECT1_1 = "NO";
    CCU2C add_3665_9 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(n78_adj_5603), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(n75_adj_5602), .D1(VCC_net), 
          .CIN(n16487), .COUT(n16488), .S0(n75_adj_5692), .S1(n72_adj_5691));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3665_9.INIT0 = 16'h9696;
    defparam add_3665_9.INIT1 = 16'h9696;
    defparam add_3665_9.INJECT1_0 = "NO";
    defparam add_3665_9.INJECT1_1 = "NO";
    CCU2C add_3665_7 (.A0(d_out_d_11__N_1882[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(n84_adj_5605), .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(n81_adj_5604), .D1(VCC_net), 
          .CIN(n16486), .COUT(n16487), .S0(n81_adj_5694), .S1(n78_adj_5693));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3665_7.INIT0 = 16'h9696;
    defparam add_3665_7.INIT1 = 16'h9696;
    defparam add_3665_7.INJECT1_0 = "NO";
    defparam add_3665_7.INJECT1_1 = "NO";
    CCU2C add_3665_5 (.A0(n90_adj_5607), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1884[17]), .B1(d_out_d_11__N_1886[17]), .C1(n87_adj_5606), 
          .D1(VCC_net), .CIN(n16485), .COUT(n16486), .S0(n87_adj_5696), 
          .S1(n84_adj_5695));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3665_5.INIT0 = 16'haaa0;
    defparam add_3665_5.INIT1 = 16'h9696;
    defparam add_3665_5.INJECT1_0 = "NO";
    defparam add_3665_5.INJECT1_1 = "NO";
    CCU2C add_3665_3 (.A0(d_out_d_11__N_1886[17]), .B0(ISquare[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16484), .COUT(n16485), .S1(n90_adj_5697));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3665_3.INIT0 = 16'h666a;
    defparam add_3665_3.INIT1 = 16'h555f;
    defparam add_3665_3.INJECT1_0 = "NO";
    defparam add_3665_3.INJECT1_1 = "NO";
    CCU2C add_3665_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1886[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16484));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3665_1.INIT0 = 16'h0000;
    defparam add_3665_1.INIT1 = 16'haaaf;
    defparam add_3665_1.INJECT1_0 = "NO";
    defparam add_3665_1.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_37 (.A0(d_d9[71]), .B0(d9[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15857), .S0(n76));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_37.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_37.INIT1 = 16'h0000;
    defparam _add_1_1424_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_37.INJECT1_1 = "NO";
    CCU2C add_3666_15 (.A0(d_out_d_11__N_1875), .B0(d_out_d_11__N_1876[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1875), .B1(d_out_d_11__N_1876[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16478), .S0(n37_adj_5681), 
          .S1(d_out_d_11__N_1878[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3666_15.INIT0 = 16'h666a;
    defparam add_3666_15.INIT1 = 16'h666a;
    defparam add_3666_15.INJECT1_0 = "NO";
    defparam add_3666_15.INJECT1_1 = "NO";
    CCU2C add_3666_13 (.A0(d_out_d_11__N_1876[17]), .B0(n36_adj_2795), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n33_adj_2796), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16477), .COUT(n16478), .S0(n43), 
          .S1(n40));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3666_13.INIT0 = 16'h9995;
    defparam add_3666_13.INIT1 = 16'h9995;
    defparam add_3666_13.INJECT1_0 = "NO";
    defparam add_3666_13.INJECT1_1 = "NO";
    CCU2C add_3666_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1876[17]), .C0(n42), 
          .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n39), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16476), .COUT(n16477), .S0(n49), .S1(n46));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3666_11.INIT0 = 16'h6969;
    defparam add_3666_11.INIT1 = 16'h9995;
    defparam add_3666_11.INJECT1_0 = "NO";
    defparam add_3666_11.INJECT1_1 = "NO";
    CCU2C add_3666_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1876[17]), .C0(n48), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1876[17]), 
          .C1(n45), .D1(VCC_net), .CIN(n16475), .COUT(n16476), .S0(n55), 
          .S1(n52));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3666_9.INIT0 = 16'h6969;
    defparam add_3666_9.INIT1 = 16'h6969;
    defparam add_3666_9.INJECT1_0 = "NO";
    defparam add_3666_9.INJECT1_1 = "NO";
    FD1S3AX ISquare_e3__i3 (.D(n120_adj_5246), .CK(CIC1_out_clkSin), .Q(ISquare[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i3.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i4 (.D(n117_adj_5245), .CK(CIC1_out_clkSin), .Q(ISquare[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i4.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i5 (.D(n114_adj_5244), .CK(CIC1_out_clkSin), .Q(ISquare[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i5.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i6 (.D(n111_adj_5243), .CK(CIC1_out_clkSin), .Q(ISquare[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i6.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i7 (.D(n108_adj_5242), .CK(CIC1_out_clkSin), .Q(ISquare[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i7.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i8 (.D(n105_adj_5241), .CK(CIC1_out_clkSin), .Q(ISquare[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i8.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i9 (.D(n102_adj_5240), .CK(CIC1_out_clkSin), .Q(ISquare[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i9.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i10 (.D(n99_adj_5239), .CK(CIC1_out_clkSin), .Q(ISquare[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i10.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i11 (.D(n96_adj_5238), .CK(CIC1_out_clkSin), .Q(ISquare[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i11.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i12 (.D(n93_adj_5237), .CK(CIC1_out_clkSin), .Q(ISquare[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i12.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i13 (.D(n90_adj_5236), .CK(CIC1_out_clkSin), .Q(ISquare[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i13.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i14 (.D(n87_adj_5235), .CK(CIC1_out_clkSin), .Q(ISquare[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i14.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i15 (.D(n84_adj_5234), .CK(CIC1_out_clkSin), .Q(ISquare[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i15.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i16 (.D(n81_adj_5233), .CK(CIC1_out_clkSin), .Q(ISquare[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i16.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i17 (.D(n78_adj_5232), .CK(CIC1_out_clkSin), .Q(ISquare[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i17.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i18 (.D(n75_adj_5231), .CK(CIC1_out_clkSin), .Q(ISquare[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i18.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i19 (.D(n72_adj_5230), .CK(CIC1_out_clkSin), .Q(ISquare[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i19.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i20 (.D(n69_adj_5229), .CK(CIC1_out_clkSin), .Q(ISquare[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i20.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i21 (.D(n66_adj_5228), .CK(CIC1_out_clkSin), .Q(ISquare[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i21.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i22 (.D(n63_adj_5227), .CK(CIC1_out_clkSin), .Q(ISquare[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i22.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i23 (.D(n60_adj_5226), .CK(CIC1_out_clkSin), .Q(ISquare[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i23.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i24 (.D(n57_adj_5225), .CK(CIC1_out_clkSin), .Q(ISquare[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i24.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i25 (.D(n54_adj_5224), .CK(CIC1_out_clkSin), .Q(ISquare[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i25.GSR = "ENABLED";
    CCU2C add_3666_7 (.A0(d_out_d_11__N_1876[17]), .B0(n17826), .C0(n54), 
          .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n51), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16474), .COUT(n16475), .S0(n61), .S1(n58));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3666_7.INIT0 = 16'h6969;
    defparam add_3666_7.INIT1 = 16'h9995;
    defparam add_3666_7.INJECT1_0 = "NO";
    defparam add_3666_7.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_adj_77 (.A(n17809), .B(n17815), .C(n18096), .D(n17810), 
         .Z(clk_80mhz_enable_1387)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;
    defparam i1_3_lut_4_lut_adj_77.init = 16'hf0b0;
    CCU2C add_3666_5 (.A0(n60), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(d_out_d_11__N_1876[17]), .C1(n57), 
          .D1(VCC_net), .CIN(n16473), .COUT(n16474), .S0(n67), .S1(n64));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3666_5.INIT0 = 16'haaa0;
    defparam add_3666_5.INIT1 = 16'h9696;
    defparam add_3666_5.INJECT1_0 = "NO";
    defparam add_3666_5.INJECT1_1 = "NO";
    CCU2C add_3666_3 (.A0(d_out_d_11__N_1876[17]), .B0(ISquare[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16472), .COUT(n16473), .S1(n70));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3666_3.INIT0 = 16'h666a;
    defparam add_3666_3.INIT1 = 16'h555f;
    defparam add_3666_3.INJECT1_0 = "NO";
    defparam add_3666_3.INJECT1_1 = "NO";
    CCU2C add_3666_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1876[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16472));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3666_1.INIT0 = 16'h0000;
    defparam add_3666_1.INIT1 = 16'haaaf;
    defparam add_3666_1.INJECT1_0 = "NO";
    defparam add_3666_1.INJECT1_1 = "NO";
    GSR GSR_INST (.GSR(VCC_net));
    CCU2C add_3655_19 (.A0(d_out_d_11__N_1882[17]), .B0(n48_adj_5191), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n45_adj_5190), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16466), .S0(n45_adj_5393), 
          .S1(d_out_d_11__N_1884[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3655_19.INIT0 = 16'h9995;
    defparam add_3655_19.INIT1 = 16'h9995;
    defparam add_3655_19.INJECT1_0 = "NO";
    defparam add_3655_19.INJECT1_1 = "NO";
    CCU2C add_3655_17 (.A0(d_out_d_11__N_1882[17]), .B0(n54_adj_5193), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n51_adj_5192), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16465), .COUT(n16466), .S0(n51_adj_5395), 
          .S1(n48_adj_5394));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3655_17.INIT0 = 16'h9995;
    defparam add_3655_17.INIT1 = 16'h9995;
    defparam add_3655_17.INJECT1_0 = "NO";
    defparam add_3655_17.INJECT1_1 = "NO";
    CCU2C add_3655_15 (.A0(d_out_d_11__N_1882[17]), .B0(n60_adj_5195), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n57_adj_5194), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16464), .COUT(n16465), .S0(n57_adj_5397), 
          .S1(n54_adj_5396));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3655_15.INIT0 = 16'h9995;
    defparam add_3655_15.INIT1 = 16'h9995;
    defparam add_3655_15.INJECT1_0 = "NO";
    defparam add_3655_15.INJECT1_1 = "NO";
    FD1P3IX phase_inc_carrGen_i0_i8 (.D(n12547), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i8.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i6 (.D(n12545), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i6.GSR = "ENABLED";
    FD1P3IX phase_inc_carrGen_i0_i4 (.D(n12543), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i4.GSR = "ENABLED";
    CCU2C add_3655_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1882[17]), .C0(n66_adj_5197), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1882[17]), 
          .C1(n63_adj_5196), .D1(VCC_net), .CIN(n16463), .COUT(n16464), 
          .S0(n63_adj_5399), .S1(n60_adj_5398));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3655_13.INIT0 = 16'h6969;
    defparam add_3655_13.INIT1 = 16'h6969;
    defparam add_3655_13.INJECT1_0 = "NO";
    defparam add_3655_13.INJECT1_1 = "NO";
    FD1P3AX phase_inc_carrGen_i0_i2 (.D(n12540), .SP(clk_80mhz_enable_1408), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i2.GSR = "ENABLED";
    CCU2C add_3655_11 (.A0(d_out_d_11__N_1882[17]), .B0(n72_adj_5199), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1882[17]), 
          .C1(n69_adj_5198), .D1(VCC_net), .CIN(n16462), .COUT(n16463), 
          .S0(n69_adj_5401), .S1(n66_adj_5400));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3655_11.INIT0 = 16'h9995;
    defparam add_3655_11.INIT1 = 16'h6969;
    defparam add_3655_11.INJECT1_0 = "NO";
    defparam add_3655_11.INJECT1_1 = "NO";
    CCU2C add_3655_9 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1882[17]), 
          .C0(n78_adj_5201), .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), 
          .B1(n17826), .C1(n75_adj_5200), .D1(VCC_net), .CIN(n16461), 
          .COUT(n16462), .S0(n75_adj_5403), .S1(n72_adj_5402));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3655_9.INIT0 = 16'h9696;
    defparam add_3655_9.INIT1 = 16'h6969;
    defparam add_3655_9.INJECT1_0 = "NO";
    defparam add_3655_9.INJECT1_1 = "NO";
    CCU2C add_3655_7 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1882[17]), 
          .C0(n84_adj_5203), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1882[17]), .C1(n81_adj_5202), .D1(VCC_net), 
          .CIN(n16460), .COUT(n16461), .S0(n81_adj_5405), .S1(n78_adj_5404));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3655_7.INIT0 = 16'h9696;
    defparam add_3655_7.INIT1 = 16'h9696;
    defparam add_3655_7.INJECT1_0 = "NO";
    defparam add_3655_7.INJECT1_1 = "NO";
    CCU2C add_3655_5 (.A0(n90_adj_5205), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1880[17]), .B1(d_out_d_11__N_1882[17]), .C1(n87_adj_5204), 
          .D1(VCC_net), .CIN(n16459), .COUT(n16460), .S0(n87_adj_5407), 
          .S1(n84_adj_5406));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3655_5.INIT0 = 16'haaa0;
    defparam add_3655_5.INIT1 = 16'h9696;
    defparam add_3655_5.INJECT1_0 = "NO";
    defparam add_3655_5.INJECT1_1 = "NO";
    CCU2C add_3655_3 (.A0(d_out_d_11__N_1882[17]), .B0(ISquare[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16458), .COUT(n16459), .S1(n90_adj_5408));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3655_3.INIT0 = 16'h666a;
    defparam add_3655_3.INIT1 = 16'h555f;
    defparam add_3655_3.INJECT1_0 = "NO";
    defparam add_3655_3.INJECT1_1 = "NO";
    CCU2C add_3655_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1882[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16458));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3655_1.INIT0 = 16'h0000;
    defparam add_3655_1.INIT1 = 16'haaaf;
    defparam add_3655_1.INJECT1_0 = "NO";
    defparam add_3655_1.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_35 (.A0(d_d9[69]), .B0(d9[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[70]), .B1(d9[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15856), .COUT(n15857), .S0(n82), .S1(n79));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_35.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_35.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_35.INJECT1_1 = "NO";
    FD1P3IX CICGain__i1 (.D(n17032), .SP(clk_80mhz_enable_1411), .CD(n12710), 
            .CK(clk_80mhz), .Q(CICGain[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam CICGain__i1.GSR = "ENABLED";
    CCU2C add_3667_19 (.A0(d_out_d_11__N_1884[17]), .B0(n48_adj_5394), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n45_adj_5393), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16452), .S0(n45_adj_5592), 
          .S1(d_out_d_11__N_1886[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3667_19.INIT0 = 16'h9995;
    defparam add_3667_19.INIT1 = 16'h9995;
    defparam add_3667_19.INJECT1_0 = "NO";
    defparam add_3667_19.INJECT1_1 = "NO";
    CCU2C add_3667_17 (.A0(d_out_d_11__N_1884[17]), .B0(n54_adj_5396), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n51_adj_5395), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16451), .COUT(n16452), .S0(n51_adj_5594), 
          .S1(n48_adj_5593));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3667_17.INIT0 = 16'h9995;
    defparam add_3667_17.INIT1 = 16'h9995;
    defparam add_3667_17.INJECT1_0 = "NO";
    defparam add_3667_17.INJECT1_1 = "NO";
    CCU2C add_3667_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1884[17]), .C0(n60_adj_5398), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n57_adj_5397), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16450), .COUT(n16451), .S0(n57_adj_5596), 
          .S1(n54_adj_5595));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3667_15.INIT0 = 16'h6969;
    defparam add_3667_15.INIT1 = 16'h9995;
    defparam add_3667_15.INJECT1_0 = "NO";
    defparam add_3667_15.INJECT1_1 = "NO";
    CCU2C add_3667_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1884[17]), .C0(n66_adj_5400), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1884[17]), 
          .C1(n63_adj_5399), .D1(VCC_net), .CIN(n16449), .COUT(n16450), 
          .S0(n63_adj_5598), .S1(n60_adj_5597));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3667_13.INIT0 = 16'h6969;
    defparam add_3667_13.INIT1 = 16'h6969;
    defparam add_3667_13.INJECT1_0 = "NO";
    defparam add_3667_13.INJECT1_1 = "NO";
    CCU2C add_3667_11 (.A0(d_out_d_11__N_1884[17]), .B0(n17826), .C0(n72_adj_5402), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n69_adj_5401), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16448), .COUT(n16449), .S0(n69_adj_5600), 
          .S1(n66_adj_5599));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3667_11.INIT0 = 16'h6969;
    defparam add_3667_11.INIT1 = 16'h9995;
    defparam add_3667_11.INJECT1_0 = "NO";
    defparam add_3667_11.INJECT1_1 = "NO";
    CCU2C add_3667_9 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(n78_adj_5404), .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1884[17]), .C1(n75_adj_5403), .D1(VCC_net), 
          .CIN(n16447), .COUT(n16448), .S0(n75_adj_5602), .S1(n72_adj_5601));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3667_9.INIT0 = 16'h9696;
    defparam add_3667_9.INIT1 = 16'h9696;
    defparam add_3667_9.INJECT1_0 = "NO";
    defparam add_3667_9.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_33 (.A0(d_d9[67]), .B0(d9[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[68]), .B1(d9[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15855), .COUT(n15856), .S0(n88), .S1(n85));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_33.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_33.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_31 (.A0(d_d9[65]), .B0(d9[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[66]), .B1(d9[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15854), .COUT(n15855), .S0(n94), .S1(n91));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_31.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_31.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_29 (.A0(d_d9[63]), .B0(d9[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[64]), .B1(d9[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15853), .COUT(n15854), .S0(n100), .S1(n97));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_29.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_29.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_27 (.A0(d_d9[61]), .B0(d9[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[62]), .B1(d9[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15852), .COUT(n15853), .S0(n106), .S1(n103));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_27.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_27.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_25 (.A0(d_d9[59]), .B0(d9[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[60]), .B1(d9[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15851), .COUT(n15852), .S0(n112), .S1(n109));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_25.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_25.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_23 (.A0(d_d9[57]), .B0(d9[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[58]), .B1(d9[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15850), .COUT(n15851), .S0(n118), .S1(n115));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_23.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_23.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_21 (.A0(d_d9[55]), .B0(d9[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[56]), .B1(d9[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15849), .COUT(n15850));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_21.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_21.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_19 (.A0(d_d9[53]), .B0(d9[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[54]), .B1(d9[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15848), .COUT(n15849));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_19.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_19.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_17 (.A0(d_d9[51]), .B0(d9[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[52]), .B1(d9[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15847), .COUT(n15848));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_17.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_17.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_15 (.A0(d_d9[49]), .B0(d9[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[50]), .B1(d9[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15846), .COUT(n15847));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_15.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_15.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_13 (.A0(d_d9[47]), .B0(d9[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[48]), .B1(d9[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15845), .COUT(n15846));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_13.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_13.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_11 (.A0(d_d9[45]), .B0(d9[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[46]), .B1(d9[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15844), .COUT(n15845));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_9 (.A0(d_d9[43]), .B0(d9[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[44]), .B1(d9[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15843), .COUT(n15844));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_7 (.A0(d_d9[41]), .B0(d9[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[42]), .B1(d9[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15842), .COUT(n15843));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_5 (.A0(d_d9[39]), .B0(d9[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[40]), .B1(d9[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15841), .COUT(n15842));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_3 (.A0(d_d9[37]), .B0(d9[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[38]), .B1(d9[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15840), .COUT(n15841));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_1424_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[36]), .B1(d9[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15840));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1424_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1424_add_4_1.INIT1 = 16'h9995;
    defparam _add_1_1424_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_38 (.A0(d3[71]), .B0(d2[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15839), .S0(n78_adj_5154));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1532_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_36 (.A0(d3[69]), .B0(d2[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[70]), .B1(d2[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15838), .COUT(n15839), .S0(n84_adj_5156), .S1(n81_adj_5155));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_34 (.A0(d3[67]), .B0(d2[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[68]), .B1(d2[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15837), .COUT(n15838), .S0(n90_adj_5158), .S1(n87_adj_5157));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_32 (.A0(d3[65]), .B0(d2[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[66]), .B1(d2[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15836), .COUT(n15837), .S0(n96_adj_5160), .S1(n93_adj_5159));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_30 (.A0(d3[63]), .B0(d2[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[64]), .B1(d2[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15835), .COUT(n15836), .S0(n102_adj_5162), .S1(n99_adj_5161));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_28 (.A0(d3[61]), .B0(d2[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[62]), .B1(d2[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15834), .COUT(n15835), .S0(n108_adj_5164), .S1(n105_adj_5163));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_26 (.A0(d3[59]), .B0(d2[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[60]), .B1(d2[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15833), .COUT(n15834), .S0(n114_adj_5166), .S1(n111_adj_5165));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_24 (.A0(d3[57]), .B0(d2[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[58]), .B1(d2[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15832), .COUT(n15833), .S0(n120_adj_5168), .S1(n117_adj_5167));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_22 (.A0(d3[55]), .B0(d2[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[56]), .B1(d2[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15831), .COUT(n15832), .S0(n126_adj_5170), .S1(n123_adj_5169));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_20 (.A0(d3[53]), .B0(d2[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[54]), .B1(d2[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15830), .COUT(n15831), .S0(n132_adj_5172), .S1(n129_adj_5171));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_18 (.A0(d3[51]), .B0(d2[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[52]), .B1(d2[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15829), .COUT(n15830), .S0(n138_adj_5174), .S1(n135_adj_5173));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_16 (.A0(d3[49]), .B0(d2[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[50]), .B1(d2[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15828), .COUT(n15829), .S0(n144_adj_5176), .S1(n141_adj_5175));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_14 (.A0(d3[47]), .B0(d2[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[48]), .B1(d2[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15827), .COUT(n15828), .S0(n150_adj_5178), .S1(n147_adj_5177));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_12 (.A0(d3[45]), .B0(d2[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[46]), .B1(d2[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15826), .COUT(n15827), .S0(n156_adj_5180), .S1(n153_adj_5179));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_10 (.A0(d3[43]), .B0(d2[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[44]), .B1(d2[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15825), .COUT(n15826), .S0(n162_adj_5182), .S1(n159_adj_5181));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_8 (.A0(d3[41]), .B0(d2[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[42]), .B1(d2[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15824), .COUT(n15825), .S0(n168_adj_5184), .S1(n165_adj_5183));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_6 (.A0(d3[39]), .B0(d2[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[40]), .B1(d2[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15823), .COUT(n15824), .S0(n174_adj_5186), .S1(n171_adj_5185));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_4 (.A0(d3[37]), .B0(d2[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[38]), .B1(d2[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15822), .COUT(n15823), .S0(n180_adj_5188), .S1(n177_adj_5187));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1532_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1532_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[36]), .B1(d2[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15822), .S1(n183_adj_5189));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1532_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1532_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1532_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1532_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_37 (.A0(d8[70]), .B0(cout_adj_5461), .C0(n81_adj_4574), 
          .D0(n3_adj_4616), .A1(d8[71]), .B1(cout_adj_5461), .C1(n78_adj_4575), 
          .D1(n2_adj_4617), .CIN(n15812), .S0(d9_71__N_1675[70]), .S1(d9_71__N_1675[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_35 (.A0(d8[68]), .B0(cout_adj_5461), .C0(n87_adj_4572), 
          .D0(n5_adj_4614), .A1(d8[69]), .B1(cout_adj_5461), .C1(n84_adj_4573), 
          .D1(n4_adj_4615), .CIN(n15811), .COUT(n15812), .S0(d9_71__N_1675[68]), 
          .S1(d9_71__N_1675[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_33 (.A0(d8[66]), .B0(cout_adj_5461), .C0(n93_adj_4570), 
          .D0(n7_adj_4612), .A1(d8[67]), .B1(cout_adj_5461), .C1(n90_adj_4571), 
          .D1(n6_adj_4613), .CIN(n15810), .COUT(n15811), .S0(d9_71__N_1675[66]), 
          .S1(d9_71__N_1675[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_31 (.A0(d8[64]), .B0(cout_adj_5461), .C0(n99_adj_4568), 
          .D0(n9_adj_4610), .A1(d8[65]), .B1(cout_adj_5461), .C1(n96_adj_4569), 
          .D1(n8_adj_4611), .CIN(n15809), .COUT(n15810), .S0(d9_71__N_1675[64]), 
          .S1(d9_71__N_1675[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_29 (.A0(d8[62]), .B0(cout_adj_5461), .C0(n105_adj_4566), 
          .D0(n11_adj_4608), .A1(d8[63]), .B1(cout_adj_5461), .C1(n102_adj_4567), 
          .D1(n10_adj_4609), .CIN(n15808), .COUT(n15809), .S0(d9_71__N_1675[62]), 
          .S1(d9_71__N_1675[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_27 (.A0(d8[60]), .B0(cout_adj_5461), .C0(n111_adj_4564), 
          .D0(n13_adj_4606), .A1(d8[61]), .B1(cout_adj_5461), .C1(n108_adj_4565), 
          .D1(n12_adj_4607), .CIN(n15807), .COUT(n15808), .S0(d9_71__N_1675[60]), 
          .S1(d9_71__N_1675[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_25 (.A0(d8[58]), .B0(cout_adj_5461), .C0(n117_adj_4562), 
          .D0(n15_adj_4604), .A1(d8[59]), .B1(cout_adj_5461), .C1(n114_adj_4563), 
          .D1(n14_adj_4605), .CIN(n15806), .COUT(n15807), .S0(d9_71__N_1675[58]), 
          .S1(d9_71__N_1675[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_23 (.A0(d8[56]), .B0(cout_adj_5461), .C0(n123), 
          .D0(n17_adj_4602), .A1(d8[57]), .B1(cout_adj_5461), .C1(n120_adj_4561), 
          .D1(n16_adj_4603), .CIN(n15805), .COUT(n15806), .S0(d9_71__N_1675[56]), 
          .S1(d9_71__N_1675[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_21 (.A0(d8[54]), .B0(cout_adj_5461), .C0(n129), 
          .D0(n19_adj_4600), .A1(d8[55]), .B1(cout_adj_5461), .C1(n126), 
          .D1(n18_adj_4601), .CIN(n15804), .COUT(n15805), .S0(d9_71__N_1675[54]), 
          .S1(d9_71__N_1675[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_19 (.A0(d8[52]), .B0(cout_adj_5461), .C0(n135), 
          .D0(n21_adj_4598), .A1(d8[53]), .B1(cout_adj_5461), .C1(n132), 
          .D1(n20_adj_4599), .CIN(n15803), .COUT(n15804), .S0(d9_71__N_1675[52]), 
          .S1(d9_71__N_1675[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_17 (.A0(d8[50]), .B0(cout_adj_5461), .C0(n141), 
          .D0(n23_adj_4596), .A1(d8[51]), .B1(cout_adj_5461), .C1(n138), 
          .D1(n22_adj_4597), .CIN(n15802), .COUT(n15803), .S0(d9_71__N_1675[50]), 
          .S1(d9_71__N_1675[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_15 (.A0(d8[48]), .B0(cout_adj_5461), .C0(n147), 
          .D0(n25_adj_4593), .A1(d8[49]), .B1(cout_adj_5461), .C1(n144), 
          .D1(n24_adj_4594), .CIN(n15801), .COUT(n15802), .S0(d9_71__N_1675[48]), 
          .S1(d9_71__N_1675[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_13 (.A0(d8[46]), .B0(cout_adj_5461), .C0(n153), 
          .D0(n27_adj_4591), .A1(d8[47]), .B1(cout_adj_5461), .C1(n150), 
          .D1(n26_adj_4592), .CIN(n15800), .COUT(n15801), .S0(d9_71__N_1675[46]), 
          .S1(d9_71__N_1675[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_11 (.A0(d8[44]), .B0(cout_adj_5461), .C0(n159), 
          .D0(n29_adj_4589), .A1(d8[45]), .B1(cout_adj_5461), .C1(n156), 
          .D1(n28_adj_4590), .CIN(n15799), .COUT(n15800), .S0(d9_71__N_1675[44]), 
          .S1(d9_71__N_1675[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_9 (.A0(d8[42]), .B0(cout_adj_5461), .C0(n165), 
          .D0(n31_adj_4587), .A1(d8[43]), .B1(cout_adj_5461), .C1(n162), 
          .D1(n30_adj_4588), .CIN(n15798), .COUT(n15799), .S0(d9_71__N_1675[42]), 
          .S1(d9_71__N_1675[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_7 (.A0(d8[40]), .B0(cout_adj_5461), .C0(n171), 
          .D0(n33_adj_4585), .A1(d8[41]), .B1(cout_adj_5461), .C1(n168), 
          .D1(n32_adj_4586), .CIN(n15797), .COUT(n15798), .S0(d9_71__N_1675[40]), 
          .S1(d9_71__N_1675[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_5 (.A0(d8[38]), .B0(cout_adj_5461), .C0(n177), 
          .D0(n35_adj_4583), .A1(d8[39]), .B1(cout_adj_5461), .C1(n174), 
          .D1(n34_adj_4584), .CIN(n15796), .COUT(n15797), .S0(d9_71__N_1675[38]), 
          .S1(d9_71__N_1675[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_3 (.A0(d8[36]), .B0(cout_adj_5461), .C0(n183), 
          .D0(n37_adj_4581), .A1(d8[37]), .B1(cout_adj_5461), .C1(n180), 
          .D1(n36_adj_4582), .CIN(n15795), .COUT(n15796), .S0(d9_71__N_1675[36]), 
          .S1(d9_71__N_1675[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1427_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1427_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5461), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15795));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1427_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1427_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1427_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15791), .S0(cout_adj_5206));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1386_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1386_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_36 (.A0(d4_adj_5713[34]), .B0(d3_adj_5712[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[35]), .B1(d3_adj_5712[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15790), .COUT(n15791), .S0(d4_71__N_634_adj_5729[34]), 
          .S1(d4_71__N_634_adj_5729[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_34 (.A0(d4_adj_5713[32]), .B0(d3_adj_5712[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[33]), .B1(d3_adj_5712[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15789), .COUT(n15790), .S0(d4_71__N_634_adj_5729[32]), 
          .S1(d4_71__N_634_adj_5729[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_32 (.A0(d4_adj_5713[30]), .B0(d3_adj_5712[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[31]), .B1(d3_adj_5712[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15788), .COUT(n15789), .S0(d4_71__N_634_adj_5729[30]), 
          .S1(d4_71__N_634_adj_5729[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_30 (.A0(d4_adj_5713[28]), .B0(d3_adj_5712[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[29]), .B1(d3_adj_5712[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15787), .COUT(n15788), .S0(d4_71__N_634_adj_5729[28]), 
          .S1(d4_71__N_634_adj_5729[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_28 (.A0(d4_adj_5713[26]), .B0(d3_adj_5712[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[27]), .B1(d3_adj_5712[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15786), .COUT(n15787), .S0(d4_71__N_634_adj_5729[26]), 
          .S1(d4_71__N_634_adj_5729[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_26 (.A0(d4_adj_5713[24]), .B0(d3_adj_5712[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[25]), .B1(d3_adj_5712[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15785), .COUT(n15786), .S0(d4_71__N_634_adj_5729[24]), 
          .S1(d4_71__N_634_adj_5729[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_24 (.A0(d4_adj_5713[22]), .B0(d3_adj_5712[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[23]), .B1(d3_adj_5712[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15784), .COUT(n15785), .S0(d4_71__N_634_adj_5729[22]), 
          .S1(d4_71__N_634_adj_5729[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_22 (.A0(d4_adj_5713[20]), .B0(d3_adj_5712[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[21]), .B1(d3_adj_5712[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15783), .COUT(n15784), .S0(d4_71__N_634_adj_5729[20]), 
          .S1(d4_71__N_634_adj_5729[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_20 (.A0(d4_adj_5713[18]), .B0(d3_adj_5712[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[19]), .B1(d3_adj_5712[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15782), .COUT(n15783), .S0(d4_71__N_634_adj_5729[18]), 
          .S1(d4_71__N_634_adj_5729[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_18 (.A0(d4_adj_5713[16]), .B0(d3_adj_5712[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[17]), .B1(d3_adj_5712[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15781), .COUT(n15782), .S0(d4_71__N_634_adj_5729[16]), 
          .S1(d4_71__N_634_adj_5729[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_16 (.A0(d4_adj_5713[14]), .B0(d3_adj_5712[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[15]), .B1(d3_adj_5712[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15780), .COUT(n15781), .S0(d4_71__N_634_adj_5729[14]), 
          .S1(d4_71__N_634_adj_5729[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_14 (.A0(d4_adj_5713[12]), .B0(d3_adj_5712[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[13]), .B1(d3_adj_5712[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15779), .COUT(n15780), .S0(d4_71__N_634_adj_5729[12]), 
          .S1(d4_71__N_634_adj_5729[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_12 (.A0(d4_adj_5713[10]), .B0(d3_adj_5712[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[11]), .B1(d3_adj_5712[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15778), .COUT(n15779), .S0(d4_71__N_634_adj_5729[10]), 
          .S1(d4_71__N_634_adj_5729[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_10 (.A0(d4_adj_5713[8]), .B0(d3_adj_5712[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[9]), .B1(d3_adj_5712[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15777), .COUT(n15778), .S0(d4_71__N_634_adj_5729[8]), 
          .S1(d4_71__N_634_adj_5729[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_8 (.A0(d4_adj_5713[6]), .B0(d3_adj_5712[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[7]), .B1(d3_adj_5712[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15776), .COUT(n15777), .S0(d4_71__N_634_adj_5729[6]), 
          .S1(d4_71__N_634_adj_5729[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_6 (.A0(d4_adj_5713[4]), .B0(d3_adj_5712[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[5]), .B1(d3_adj_5712[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15775), .COUT(n15776), .S0(d4_71__N_634_adj_5729[4]), 
          .S1(d4_71__N_634_adj_5729[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_4 (.A0(d4_adj_5713[2]), .B0(d3_adj_5712[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[3]), .B1(d3_adj_5712[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15774), .COUT(n15775), .S0(d4_71__N_634_adj_5729[2]), 
          .S1(d4_71__N_634_adj_5729[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1386_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1386_add_4_2 (.A0(d4_adj_5713[0]), .B0(d3_adj_5712[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5713[1]), .B1(d3_adj_5712[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15774), .S1(d4_71__N_634_adj_5729[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1386_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1386_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1386_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1386_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1377_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15772), .S0(n36_adj_2807));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1377_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1377_add_4_17.INIT1 = 16'h0000;
    defparam _add_1_1377_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1377_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1377_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15771), .COUT(n15772), .S0(n42_adj_2805), 
          .S1(n39_adj_2806));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1377_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1377_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1377_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1377_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1377_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15770), .COUT(n15771), .S0(n48_adj_2803), 
          .S1(n45_adj_2804));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1377_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1377_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1377_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1377_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1377_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15769), .COUT(n15770), .S0(n54_adj_2801), 
          .S1(n51_adj_2802));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1377_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1377_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1377_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1377_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1377_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15768), .COUT(n15769), .S0(n60_adj_2799), .S1(n57_adj_2800));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1377_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1377_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1377_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1377_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1377_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15767), .COUT(n15768), .S0(n66), .S1(n63));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1377_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1377_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1377_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1377_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1377_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15766), .COUT(n15767), .S0(n72), .S1(n69));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1377_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1377_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1377_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1377_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1377_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15765), .COUT(n15766), .S0(n78), .S1(n75));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1377_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1377_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1377_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1377_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1377_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15765), .S1(n81));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1377_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1377_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1377_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1377_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15764), .S0(cout_adj_5207));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1389_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1389_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_36 (.A0(d5_adj_5714[34]), .B0(d4_adj_5713[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[35]), .B1(d4_adj_5713[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15763), .COUT(n15764), .S0(d5_71__N_706_adj_5730[34]), 
          .S1(d5_71__N_706_adj_5730[35]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_34 (.A0(d5_adj_5714[32]), .B0(d4_adj_5713[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[33]), .B1(d4_adj_5713[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15762), .COUT(n15763), .S0(d5_71__N_706_adj_5730[32]), 
          .S1(d5_71__N_706_adj_5730[33]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_32 (.A0(d5_adj_5714[30]), .B0(d4_adj_5713[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[31]), .B1(d4_adj_5713[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15761), .COUT(n15762), .S0(d5_71__N_706_adj_5730[30]), 
          .S1(d5_71__N_706_adj_5730[31]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_30 (.A0(d5_adj_5714[28]), .B0(d4_adj_5713[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[29]), .B1(d4_adj_5713[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15760), .COUT(n15761), .S0(d5_71__N_706_adj_5730[28]), 
          .S1(d5_71__N_706_adj_5730[29]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_28 (.A0(d5_adj_5714[26]), .B0(d4_adj_5713[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[27]), .B1(d4_adj_5713[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15759), .COUT(n15760), .S0(d5_71__N_706_adj_5730[26]), 
          .S1(d5_71__N_706_adj_5730[27]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_26 (.A0(d5_adj_5714[24]), .B0(d4_adj_5713[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[25]), .B1(d4_adj_5713[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15758), .COUT(n15759), .S0(d5_71__N_706_adj_5730[24]), 
          .S1(d5_71__N_706_adj_5730[25]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_24 (.A0(d5_adj_5714[22]), .B0(d4_adj_5713[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[23]), .B1(d4_adj_5713[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15757), .COUT(n15758), .S0(d5_71__N_706_adj_5730[22]), 
          .S1(d5_71__N_706_adj_5730[23]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_22 (.A0(d5_adj_5714[20]), .B0(d4_adj_5713[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[21]), .B1(d4_adj_5713[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15756), .COUT(n15757), .S0(d5_71__N_706_adj_5730[20]), 
          .S1(d5_71__N_706_adj_5730[21]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_20 (.A0(d5_adj_5714[18]), .B0(d4_adj_5713[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[19]), .B1(d4_adj_5713[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15755), .COUT(n15756), .S0(d5_71__N_706_adj_5730[18]), 
          .S1(d5_71__N_706_adj_5730[19]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_18 (.A0(d5_adj_5714[16]), .B0(d4_adj_5713[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[17]), .B1(d4_adj_5713[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15754), .COUT(n15755), .S0(d5_71__N_706_adj_5730[16]), 
          .S1(d5_71__N_706_adj_5730[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_16 (.A0(d5_adj_5714[14]), .B0(d4_adj_5713[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[15]), .B1(d4_adj_5713[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15753), .COUT(n15754), .S0(d5_71__N_706_adj_5730[14]), 
          .S1(d5_71__N_706_adj_5730[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_14 (.A0(d5_adj_5714[12]), .B0(d4_adj_5713[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[13]), .B1(d4_adj_5713[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15752), .COUT(n15753), .S0(d5_71__N_706_adj_5730[12]), 
          .S1(d5_71__N_706_adj_5730[13]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_12 (.A0(d5_adj_5714[10]), .B0(d4_adj_5713[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[11]), .B1(d4_adj_5713[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15751), .COUT(n15752), .S0(d5_71__N_706_adj_5730[10]), 
          .S1(d5_71__N_706_adj_5730[11]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_10 (.A0(d5_adj_5714[8]), .B0(d4_adj_5713[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[9]), .B1(d4_adj_5713[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15750), .COUT(n15751), .S0(d5_71__N_706_adj_5730[8]), 
          .S1(d5_71__N_706_adj_5730[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_8 (.A0(d5_adj_5714[6]), .B0(d4_adj_5713[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[7]), .B1(d4_adj_5713[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15749), .COUT(n15750), .S0(d5_71__N_706_adj_5730[6]), 
          .S1(d5_71__N_706_adj_5730[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_6 (.A0(d5_adj_5714[4]), .B0(d4_adj_5713[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[5]), .B1(d4_adj_5713[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15748), .COUT(n15749), .S0(d5_71__N_706_adj_5730[4]), 
          .S1(d5_71__N_706_adj_5730[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_4 (.A0(d5_adj_5714[2]), .B0(d4_adj_5713[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[3]), .B1(d4_adj_5713[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15747), .COUT(n15748), .S0(d5_71__N_706_adj_5730[2]), 
          .S1(d5_71__N_706_adj_5730[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1389_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1389_add_4_2 (.A0(d5_adj_5714[0]), .B0(d4_adj_5713[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[1]), .B1(d4_adj_5713[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15747), .S1(d5_71__N_706_adj_5730[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1389_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1389_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1389_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1389_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_37 (.A0(d7[70]), .B0(cout_adj_5575), .C0(n81_adj_5646), 
          .D0(n3_adj_4652), .A1(d7[71]), .B1(cout_adj_5575), .C1(n78_adj_5645), 
          .D1(n2_adj_4653), .CIN(n15744), .S0(d8_71__N_1603[70]), .S1(d8_71__N_1603[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_35 (.A0(d7[68]), .B0(cout_adj_5575), .C0(n87_adj_5648), 
          .D0(n5_adj_4650), .A1(d7[69]), .B1(cout_adj_5575), .C1(n84_adj_5647), 
          .D1(n4_adj_4651), .CIN(n15743), .COUT(n15744), .S0(d8_71__N_1603[68]), 
          .S1(d8_71__N_1603[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_33 (.A0(d7[66]), .B0(cout_adj_5575), .C0(n93_adj_5650), 
          .D0(n7_adj_4648), .A1(d7[67]), .B1(cout_adj_5575), .C1(n90_adj_5649), 
          .D1(n6_adj_4649), .CIN(n15742), .COUT(n15743), .S0(d8_71__N_1603[66]), 
          .S1(d8_71__N_1603[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_31 (.A0(d7[64]), .B0(cout_adj_5575), .C0(n99_adj_5652), 
          .D0(n9_adj_4646), .A1(d7[65]), .B1(cout_adj_5575), .C1(n96_adj_5651), 
          .D1(n8_adj_4647), .CIN(n15741), .COUT(n15742), .S0(d8_71__N_1603[64]), 
          .S1(d8_71__N_1603[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_29 (.A0(d7[62]), .B0(cout_adj_5575), .C0(n105_adj_5654), 
          .D0(n11_adj_4644), .A1(d7[63]), .B1(cout_adj_5575), .C1(n102_adj_5653), 
          .D1(n10_adj_4645), .CIN(n15740), .COUT(n15741), .S0(d8_71__N_1603[62]), 
          .S1(d8_71__N_1603[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_27 (.A0(d7[60]), .B0(cout_adj_5575), .C0(n111_adj_5656), 
          .D0(n13_adj_4642), .A1(d7[61]), .B1(cout_adj_5575), .C1(n108_adj_5655), 
          .D1(n12_adj_4643), .CIN(n15739), .COUT(n15740), .S0(d8_71__N_1603[60]), 
          .S1(d8_71__N_1603[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_25 (.A0(d7[58]), .B0(cout_adj_5575), .C0(n117_adj_5658), 
          .D0(n15_adj_4640), .A1(d7[59]), .B1(cout_adj_5575), .C1(n114_adj_5657), 
          .D1(n14_adj_4641), .CIN(n15738), .COUT(n15739), .S0(d8_71__N_1603[58]), 
          .S1(d8_71__N_1603[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_23 (.A0(d7[56]), .B0(cout_adj_5575), .C0(n123_adj_5660), 
          .D0(n17_adj_4638), .A1(d7[57]), .B1(cout_adj_5575), .C1(n120_adj_5659), 
          .D1(n16_adj_4639), .CIN(n15737), .COUT(n15738), .S0(d8_71__N_1603[56]), 
          .S1(d8_71__N_1603[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_21 (.A0(d7[54]), .B0(cout_adj_5575), .C0(n129_adj_5662), 
          .D0(n19_adj_4636), .A1(d7[55]), .B1(cout_adj_5575), .C1(n126_adj_5661), 
          .D1(n18_adj_4637), .CIN(n15736), .COUT(n15737), .S0(d8_71__N_1603[54]), 
          .S1(d8_71__N_1603[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_19 (.A0(d7[52]), .B0(cout_adj_5575), .C0(n135_adj_5664), 
          .D0(n21_adj_4634), .A1(d7[53]), .B1(cout_adj_5575), .C1(n132_adj_5663), 
          .D1(n20_adj_4635), .CIN(n15735), .COUT(n15736), .S0(d8_71__N_1603[52]), 
          .S1(d8_71__N_1603[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_17 (.A0(d7[50]), .B0(cout_adj_5575), .C0(n141_adj_5666), 
          .D0(n23_adj_4632), .A1(d7[51]), .B1(cout_adj_5575), .C1(n138_adj_5665), 
          .D1(n22_adj_4633), .CIN(n15734), .COUT(n15735), .S0(d8_71__N_1603[50]), 
          .S1(d8_71__N_1603[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_15 (.A0(d7[48]), .B0(cout_adj_5575), .C0(n147_adj_5668), 
          .D0(n25_adj_4630), .A1(d7[49]), .B1(cout_adj_5575), .C1(n144_adj_5667), 
          .D1(n24_adj_4631), .CIN(n15733), .COUT(n15734), .S0(d8_71__N_1603[48]), 
          .S1(d8_71__N_1603[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_13 (.A0(d7[46]), .B0(cout_adj_5575), .C0(n153_adj_5670), 
          .D0(n27_adj_4628), .A1(d7[47]), .B1(cout_adj_5575), .C1(n150_adj_5669), 
          .D1(n26_adj_4629), .CIN(n15732), .COUT(n15733), .S0(d8_71__N_1603[46]), 
          .S1(d8_71__N_1603[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_11 (.A0(d7[44]), .B0(cout_adj_5575), .C0(n159_adj_5672), 
          .D0(n29_adj_4626), .A1(d7[45]), .B1(cout_adj_5575), .C1(n156_adj_5671), 
          .D1(n28_adj_4627), .CIN(n15731), .COUT(n15732), .S0(d8_71__N_1603[44]), 
          .S1(d8_71__N_1603[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_9 (.A0(d7[42]), .B0(cout_adj_5575), .C0(n165_adj_5674), 
          .D0(n31_adj_4624), .A1(d7[43]), .B1(cout_adj_5575), .C1(n162_adj_5673), 
          .D1(n30_adj_4625), .CIN(n15730), .COUT(n15731), .S0(d8_71__N_1603[42]), 
          .S1(d8_71__N_1603[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_7 (.A0(d7[40]), .B0(cout_adj_5575), .C0(n171_adj_5676), 
          .D0(n33_adj_4622), .A1(d7[41]), .B1(cout_adj_5575), .C1(n168_adj_5675), 
          .D1(n32_adj_4623), .CIN(n15729), .COUT(n15730), .S0(d8_71__N_1603[40]), 
          .S1(d8_71__N_1603[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_5 (.A0(d7[38]), .B0(cout_adj_5575), .C0(n177_adj_5678), 
          .D0(n35_adj_4620), .A1(d7[39]), .B1(cout_adj_5575), .C1(n174_adj_5677), 
          .D1(n34_adj_4621), .CIN(n15728), .COUT(n15729), .S0(d8_71__N_1603[38]), 
          .S1(d8_71__N_1603[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_3 (.A0(d7[36]), .B0(cout_adj_5575), .C0(n183_adj_5680), 
          .D0(n37_adj_4618), .A1(d7[37]), .B1(cout_adj_5575), .C1(n180_adj_5679), 
          .D1(n36_adj_4619), .CIN(n15727), .COUT(n15728), .S0(d8_71__N_1603[36]), 
          .S1(d8_71__N_1603[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1430_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1430_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5575), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15727));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1430_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1430_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1430_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1392_add_4_17 (.A0(count_adj_5725[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15723), .S0(n36_adj_5208));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1392_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1392_add_4_17.INIT1 = 16'h0000;
    defparam _add_1_1392_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1392_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1392_add_4_15 (.A0(count_adj_5725[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5725[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15722), .COUT(n15723), .S0(n42_adj_5210), 
          .S1(n39_adj_5209));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1392_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1392_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1392_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1392_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1392_add_4_13 (.A0(count_adj_5725[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5725[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15721), .COUT(n15722), .S0(n48_adj_5212), 
          .S1(n45_adj_5211));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1392_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1392_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1392_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1392_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1392_add_4_11 (.A0(count_adj_5725[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5725[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15720), .COUT(n15721), .S0(n54_adj_5214), 
          .S1(n51_adj_5213));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1392_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1392_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1392_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1392_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1392_add_4_9 (.A0(count_adj_5725[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5725[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15719), .COUT(n15720), .S0(n60_adj_5216), 
          .S1(n57_adj_5215));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1392_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1392_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1392_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1392_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1392_add_4_7 (.A0(count_adj_5725[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5725[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15718), .COUT(n15719), .S0(n66_adj_5218), 
          .S1(n63_adj_5217));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1392_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1392_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1392_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1392_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1392_add_4_5 (.A0(count_adj_5725[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5725[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15717), .COUT(n15718), .S0(n72_adj_5220), 
          .S1(n69_adj_5219));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1392_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1392_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1392_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1392_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1392_add_4_3 (.A0(count_adj_5725[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5725[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15716), .COUT(n15717), .S0(n78_adj_5222), 
          .S1(n75_adj_5221));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1392_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1392_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1392_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1392_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1392_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_adj_5725[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15716), .S1(n81_adj_5223));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1392_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1392_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1392_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1392_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_37 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n81_adj_5083), .D0(d1[70]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n78_adj_5082), .D1(d1[71]), .CIN(n15714), .S0(d1_71__N_418[70]), 
          .S1(d1_71__N_418[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_35 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n87_adj_5085), .D0(d1[68]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n84_adj_5084), .D1(d1[69]), .CIN(n15713), .COUT(n15714), 
          .S0(d1_71__N_418[68]), .S1(d1_71__N_418[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_33 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n93_adj_5087), .D0(d1[66]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n90_adj_5086), .D1(d1[67]), .CIN(n15712), .COUT(n15713), 
          .S0(d1_71__N_418[66]), .S1(d1_71__N_418[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_31 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n99_adj_5089), .D0(d1[64]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n96_adj_5088), .D1(d1[65]), .CIN(n15711), .COUT(n15712), 
          .S0(d1_71__N_418[64]), .S1(d1_71__N_418[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_29 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n105_adj_5091), .D0(d1[62]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n102_adj_5090), .D1(d1[63]), .CIN(n15710), .COUT(n15711), 
          .S0(d1_71__N_418[62]), .S1(d1_71__N_418[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_27 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n111_adj_5093), .D0(d1[60]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n108_adj_5092), .D1(d1[61]), .CIN(n15709), .COUT(n15710), 
          .S0(d1_71__N_418[60]), .S1(d1_71__N_418[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_25 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n117_adj_5095), .D0(d1[58]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n114_adj_5094), .D1(d1[59]), .CIN(n15708), .COUT(n15709), 
          .S0(d1_71__N_418[58]), .S1(d1_71__N_418[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_23 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n123_adj_5097), .D0(d1[56]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n120_adj_5096), .D1(d1[57]), .CIN(n15707), .COUT(n15708), 
          .S0(d1_71__N_418[56]), .S1(d1_71__N_418[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_21 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n129_adj_5099), .D0(d1[54]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n126_adj_5098), .D1(d1[55]), .CIN(n15706), .COUT(n15707), 
          .S0(d1_71__N_418[54]), .S1(d1_71__N_418[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_19 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n135_adj_5101), .D0(d1[52]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n132_adj_5100), .D1(d1[53]), .CIN(n15705), .COUT(n15706), 
          .S0(d1_71__N_418[52]), .S1(d1_71__N_418[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_17 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n141_adj_5103), .D0(d1[50]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n138_adj_5102), .D1(d1[51]), .CIN(n15704), .COUT(n15705), 
          .S0(d1_71__N_418[50]), .S1(d1_71__N_418[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_17.INJECT1_1 = "NO";
    CCU2C add_3667_7 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(n84_adj_5406), .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(d_out_d_11__N_1884[17]), .C1(n81_adj_5405), .D1(VCC_net), 
          .CIN(n16446), .COUT(n16447), .S0(n81_adj_5604), .S1(n78_adj_5603));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3667_7.INIT0 = 16'h9696;
    defparam add_3667_7.INIT1 = 16'h9696;
    defparam add_3667_7.INJECT1_0 = "NO";
    defparam add_3667_7.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_18 (.A0(d_d6_adj_5716[15]), .B0(d6_adj_5715[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[16]), .B1(d6_adj_5715[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16254), .COUT(n16255), .S0(d7_71__N_1531_adj_5743[15]), 
          .S1(d7_71__N_1531_adj_5743[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_16 (.A0(d_d6_adj_5716[13]), .B0(d6_adj_5715[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[14]), .B1(d6_adj_5715[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16253), .COUT(n16254), .S0(d7_71__N_1531_adj_5743[13]), 
          .S1(d7_71__N_1531_adj_5743[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_15 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n147_adj_5105), .D0(d1[48]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n144_adj_5104), .D1(d1[49]), .CIN(n15703), .COUT(n15704), 
          .S0(d1_71__N_418[48]), .S1(d1_71__N_418[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_15.INJECT1_1 = "NO";
    CCU2C add_3667_5 (.A0(n90_adj_5408), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1882[17]), .B1(d_out_d_11__N_1884[17]), .C1(n87_adj_5407), 
          .D1(VCC_net), .CIN(n16445), .COUT(n16446), .S0(n87_adj_5606), 
          .S1(n84_adj_5605));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3667_5.INIT0 = 16'haaa0;
    defparam add_3667_5.INIT1 = 16'h9696;
    defparam add_3667_5.INJECT1_0 = "NO";
    defparam add_3667_5.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_14 (.A0(d_d6_adj_5716[11]), .B0(d6_adj_5715[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[12]), .B1(d6_adj_5715[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16252), .COUT(n16253), .S0(d7_71__N_1531_adj_5743[11]), 
          .S1(d7_71__N_1531_adj_5743[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_13 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n153_adj_5107), .D0(d1[46]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n150_adj_5106), .D1(d1[47]), .CIN(n15702), .COUT(n15703), 
          .S0(d1_71__N_418[46]), .S1(d1_71__N_418[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_13.INJECT1_1 = "NO";
    CCU2C add_3667_3 (.A0(d_out_d_11__N_1884[17]), .B0(ISquare[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16444), .COUT(n16445), .S1(n90_adj_5607));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3667_3.INIT0 = 16'h666a;
    defparam add_3667_3.INIT1 = 16'h555f;
    defparam add_3667_3.INJECT1_0 = "NO";
    defparam add_3667_3.INJECT1_1 = "NO";
    CCU2C add_3667_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1884[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16444));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3667_1.INIT0 = 16'h0000;
    defparam add_3667_1.INIT1 = 16'haaaf;
    defparam add_3667_1.INJECT1_0 = "NO";
    defparam add_3667_1.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_12 (.A0(d_d6_adj_5716[9]), .B0(d6_adj_5715[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[10]), .B1(d6_adj_5715[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16251), .COUT(n16252), .S0(d7_71__N_1531_adj_5743[9]), 
          .S1(d7_71__N_1531_adj_5743[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_10 (.A0(d_d6_adj_5716[7]), .B0(d6_adj_5715[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[8]), .B1(d6_adj_5715[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16250), .COUT(n16251), .S0(d7_71__N_1531_adj_5743[7]), 
          .S1(d7_71__N_1531_adj_5743[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_10.INJECT1_1 = "NO";
    CCU2C add_3660_65 (.A0(phase_inc_carrGen[62]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(phase_inc_carrGen[63]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16438), .S0(n137), .S1(n134));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_65.INIT0 = 16'haa6a;
    defparam add_3660_65.INIT1 = 16'haa6a;
    defparam add_3660_65.INJECT1_0 = "NO";
    defparam add_3660_65.INJECT1_1 = "NO";
    CCU2C add_3660_63 (.A0(phase_inc_carrGen[60]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(phase_inc_carrGen[61]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16437), .COUT(n16438), .S0(n143), .S1(n140));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_63.INIT0 = 16'haa6a;
    defparam add_3660_63.INIT1 = 16'haa6a;
    defparam add_3660_63.INJECT1_0 = "NO";
    defparam add_3660_63.INJECT1_1 = "NO";
    CCU2C add_3660_61 (.A0(phase_inc_carrGen[58]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(phase_inc_carrGen[59]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16436), .COUT(n16437), .S0(n149), .S1(n146));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_61.INIT0 = 16'haa6a;
    defparam add_3660_61.INIT1 = 16'haa6a;
    defparam add_3660_61.INJECT1_0 = "NO";
    defparam add_3660_61.INJECT1_1 = "NO";
    CCU2C add_3660_59 (.A0(phase_inc_carrGen[56]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(phase_inc_carrGen[57]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16435), .COUT(n16436), .S0(n155), .S1(n152));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_59.INIT0 = 16'haa6a;
    defparam add_3660_59.INIT1 = 16'haa6a;
    defparam add_3660_59.INJECT1_0 = "NO";
    defparam add_3660_59.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_8 (.A0(d_d6_adj_5716[5]), .B0(d6_adj_5715[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[6]), .B1(d6_adj_5715[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16249), .COUT(n16250), .S0(d7_71__N_1531_adj_5743[5]), 
          .S1(d7_71__N_1531_adj_5743[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_6 (.A0(d_d6_adj_5716[3]), .B0(d6_adj_5715[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[4]), .B1(d6_adj_5715[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16248), .COUT(n16249), .S0(d7_71__N_1531_adj_5743[3]), 
          .S1(d7_71__N_1531_adj_5743[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_6.INJECT1_1 = "NO";
    CCU2C add_3660_57 (.A0(phase_inc_carrGen[54]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(phase_inc_carrGen[55]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16434), .COUT(n16435), .S0(n161), .S1(n158));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_57.INIT0 = 16'haa6a;
    defparam add_3660_57.INIT1 = 16'haa6a;
    defparam add_3660_57.INJECT1_0 = "NO";
    defparam add_3660_57.INJECT1_1 = "NO";
    CCU2C add_3660_55 (.A0(phase_inc_carrGen[52]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(phase_inc_carrGen[53]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16433), .COUT(n16434), .S0(n167), .S1(n164));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_55.INIT0 = 16'haa6a;
    defparam add_3660_55.INIT1 = 16'haa6a;
    defparam add_3660_55.INJECT1_0 = "NO";
    defparam add_3660_55.INJECT1_1 = "NO";
    CCU2C add_3660_53 (.A0(phase_inc_carrGen[50]), .B0(led_c_4), .C0(n17820), 
          .D0(led_c_2), .A1(phase_inc_carrGen[51]), .B1(n17825), .C1(n12424), 
          .D1(led_c_4), .CIN(n16432), .COUT(n16433), .S0(n173), .S1(n170));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_53.INIT0 = 16'h959a;
    defparam add_3660_53.INIT1 = 16'haa6a;
    defparam add_3660_53.INJECT1_0 = "NO";
    defparam add_3660_53.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_4 (.A0(d_d6_adj_5716[1]), .B0(d6_adj_5715[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5716[2]), .B1(d6_adj_5715[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16247), .COUT(n16248), .S0(d7_71__N_1531_adj_5743[1]), 
          .S1(d7_71__N_1531_adj_5743[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1478_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_4.INJECT1_1 = "NO";
    CCU2C add_3660_51 (.A0(phase_inc_carrGen[48]), .B0(n18053), .C0(n17820), 
          .D0(led_c_2), .A1(phase_inc_carrGen[49]), .B1(n18053), .C1(n17820), 
          .D1(led_c_2), .CIN(n16431), .COUT(n16432), .S0(n179), .S1(n176));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_51.INIT0 = 16'h959a;
    defparam add_3660_51.INIT1 = 16'h959a;
    defparam add_3660_51.INJECT1_0 = "NO";
    defparam add_3660_51.INJECT1_1 = "NO";
    CCU2C add_3660_49 (.A0(n3728), .B0(phase_inc_carrGen[46]), .C0(GND_net), 
          .D0(VCC_net), .A1(n3728), .B1(phase_inc_carrGen[47]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16430), .COUT(n16431), .S0(n185), .S1(n182));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_49.INIT0 = 16'h9995;
    defparam add_3660_49.INIT1 = 16'h9995;
    defparam add_3660_49.INJECT1_0 = "NO";
    defparam add_3660_49.INJECT1_1 = "NO";
    CCU2C add_3660_47 (.A0(phase_inc_carrGen[44]), .B0(n17820), .C0(n18053), 
          .D0(led_c_2), .A1(phase_inc_carrGen[45]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16429), .COUT(n16430), .S0(n191), .S1(n188));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_47.INIT0 = 16'h596a;
    defparam add_3660_47.INIT1 = 16'haa6a;
    defparam add_3660_47.INJECT1_0 = "NO";
    defparam add_3660_47.INJECT1_1 = "NO";
    CCU2C _add_1_1478_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6_adj_5716[0]), .B1(d6_adj_5715[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16247), .S1(d7_71__N_1531_adj_5743[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1478_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1478_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1478_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1478_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_38 (.A0(d_d6[71]), .B0(d6[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16246), .S0(n78_adj_5465));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1559_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_38.INJECT1_1 = "NO";
    CCU2C add_3660_45 (.A0(phase_inc_carrGen[42]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(n18053), .B1(n17820), .C1(phase_inc_carrGen[43]), 
          .D1(VCC_net), .CIN(n16428), .COUT(n16429), .S0(n197), .S1(n194));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_45.INIT0 = 16'h6aaa;
    defparam add_3660_45.INIT1 = 16'h8787;
    defparam add_3660_45.INJECT1_0 = "NO";
    defparam add_3660_45.INJECT1_1 = "NO";
    CCU2C add_3660_43 (.A0(phase_inc_carrGen[40]), .B0(n18053), .C0(n17820), 
          .D0(led_c_2), .A1(n18053), .B1(n17820), .C1(phase_inc_carrGen[41]), 
          .D1(VCC_net), .CIN(n16427), .COUT(n16428), .S0(n203), .S1(n200));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_43.INIT0 = 16'h959a;
    defparam add_3660_43.INIT1 = 16'h8787;
    defparam add_3660_43.INJECT1_0 = "NO";
    defparam add_3660_43.INJECT1_1 = "NO";
    CCU2C add_3660_41 (.A0(phase_inc_carrGen[38]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(phase_inc_carrGen[39]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16426), .COUT(n16427), .S0(n209), .S1(n206));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_41.INIT0 = 16'haa6a;
    defparam add_3660_41.INIT1 = 16'haa6a;
    defparam add_3660_41.INJECT1_0 = "NO";
    defparam add_3660_41.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_36 (.A0(d_d6[69]), .B0(d6[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[70]), .B1(d6[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16245), .COUT(n16246), .S0(n84_adj_5467), .S1(n81_adj_5466));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_36.INJECT1_1 = "NO";
    CCU2C add_3660_39 (.A0(phase_inc_carrGen[36]), .B0(n17820), .C0(n18053), 
          .D0(led_c_2), .A1(n18053), .B1(n17820), .C1(phase_inc_carrGen[37]), 
          .D1(VCC_net), .CIN(n16425), .COUT(n16426), .S0(n215), .S1(n212));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_39.INIT0 = 16'h596a;
    defparam add_3660_39.INIT1 = 16'h4b4b;
    defparam add_3660_39.INJECT1_0 = "NO";
    defparam add_3660_39.INJECT1_1 = "NO";
    CCU2C add_3660_37 (.A0(phase_inc_carrGen[34]), .B0(n17820), .C0(n18053), 
          .D0(led_c_2), .A1(phase_inc_carrGen[35]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16424), .COUT(n16425), .S0(n221), .S1(n218));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_37.INIT0 = 16'h596a;
    defparam add_3660_37.INIT1 = 16'haa6a;
    defparam add_3660_37.INJECT1_0 = "NO";
    defparam add_3660_37.INJECT1_1 = "NO";
    CCU2C add_3660_35 (.A0(phase_inc_carrGen[32]), .B0(n18053), .C0(n17820), 
          .D0(led_c_2), .A1(n18053), .B1(n17820), .C1(phase_inc_carrGen[33]), 
          .D1(VCC_net), .CIN(n16423), .COUT(n16424), .S0(n227), .S1(n224));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_35.INIT0 = 16'h959a;
    defparam add_3660_35.INIT1 = 16'h4b4b;
    defparam add_3660_35.INJECT1_0 = "NO";
    defparam add_3660_35.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_34 (.A0(d_d6[67]), .B0(d6[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[68]), .B1(d6[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16244), .COUT(n16245), .S0(n90_adj_5469), .S1(n87_adj_5468));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_29 (.A0(d4[62]), .B0(cout_adj_2810), .C0(n105_adj_5294), 
          .D0(d5[62]), .A1(d4[63]), .B1(cout_adj_2810), .C1(n102_adj_5293), 
          .D1(d5[63]), .CIN(n16057), .COUT(n16058), .S0(d5_71__N_706[62]), 
          .S1(d5_71__N_706[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_29.INJECT1_1 = "NO";
    CCU2C add_3660_33 (.A0(phase_inc_carrGen[30]), .B0(n18053), .C0(n17820), 
          .D0(led_c_2), .A1(phase_inc_carrGen[31]), .B1(n17820), .C1(n18053), 
          .D1(n3674), .CIN(n16422), .COUT(n16423), .S0(n233), .S1(n230));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_33.INIT0 = 16'h959a;
    defparam add_3660_33.INIT1 = 16'h596a;
    defparam add_3660_33.INJECT1_0 = "NO";
    defparam add_3660_33.INJECT1_1 = "NO";
    CCU2C add_3660_31 (.A0(n18053), .B0(n17820), .C0(phase_inc_carrGen[28]), 
          .D0(VCC_net), .A1(phase_inc_carrGen[29]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16421), .COUT(n16422), .S0(n239), .S1(n236));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_31.INIT0 = 16'h8787;
    defparam add_3660_31.INIT1 = 16'h6aaa;
    defparam add_3660_31.INJECT1_0 = "NO";
    defparam add_3660_31.INJECT1_1 = "NO";
    CCU2C add_3660_29 (.A0(phase_inc_carrGen[26]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(n18053), .B1(n17820), .C1(phase_inc_carrGen[27]), 
          .D1(VCC_net), .CIN(n16420), .COUT(n16421), .S0(n245), .S1(n242));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_29.INIT0 = 16'haa6a;
    defparam add_3660_29.INIT1 = 16'h4b4b;
    defparam add_3660_29.INJECT1_0 = "NO";
    defparam add_3660_29.INJECT1_1 = "NO";
    CCU2C add_3660_27 (.A0(phase_inc_carrGen[24]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(phase_inc_carrGen[25]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16419), .COUT(n16420), .S0(n251), .S1(n248));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_27.INIT0 = 16'haa6a;
    defparam add_3660_27.INIT1 = 16'haa6a;
    defparam add_3660_27.INJECT1_0 = "NO";
    defparam add_3660_27.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_28 (.A0(d5_adj_5714[61]), .B0(d4_adj_5713[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[62]), .B1(d4_adj_5713[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16165), .COUT(n16166), .S0(n108_adj_5548), 
          .S1(n105_adj_5547));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_28.INJECT1_1 = "NO";
    CCU2C add_3660_25 (.A0(phase_inc_carrGen[22]), .B0(n17820), .C0(n18053), 
          .D0(led_c_2), .A1(phase_inc_carrGen[23]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16418), .COUT(n16419), .S0(n257), .S1(n254));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_25.INIT0 = 16'h596a;
    defparam add_3660_25.INIT1 = 16'h6aaa;
    defparam add_3660_25.INJECT1_0 = "NO";
    defparam add_3660_25.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_26 (.A0(d5_adj_5714[59]), .B0(d4_adj_5713[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[60]), .B1(d4_adj_5713[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16164), .COUT(n16165), .S0(n114_adj_5550), 
          .S1(n111_adj_5549));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_26.INJECT1_1 = "NO";
    CCU2C add_3660_23 (.A0(phase_inc_carrGen[20]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(phase_inc_carrGen[21]), .B1(n18053), .C1(n17820), 
          .D1(led_c_2), .CIN(n16417), .COUT(n16418), .S0(n263), .S1(n260));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_23.INIT0 = 16'haa6a;
    defparam add_3660_23.INIT1 = 16'h959a;
    defparam add_3660_23.INJECT1_0 = "NO";
    defparam add_3660_23.INJECT1_1 = "NO";
    CCU2C add_3660_21 (.A0(phase_inc_carrGen[18]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(n18053), .B1(n17820), .C1(phase_inc_carrGen[19]), 
          .D1(VCC_net), .CIN(n16416), .COUT(n16417), .S0(n269), .S1(n266));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_21.INIT0 = 16'h6aaa;
    defparam add_3660_21.INIT1 = 16'h4b4b;
    defparam add_3660_21.INJECT1_0 = "NO";
    defparam add_3660_21.INJECT1_1 = "NO";
    CCU2C add_3660_19 (.A0(phase_inc_carrGen[16]), .B0(n17820), .C0(n18053), 
          .D0(n3674), .A1(n3728), .B1(phase_inc_carrGen[17]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16415), .COUT(n16416), .S0(n275), .S1(n272));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_19.INIT0 = 16'h596a;
    defparam add_3660_19.INIT1 = 16'h9995;
    defparam add_3660_19.INJECT1_0 = "NO";
    defparam add_3660_19.INJECT1_1 = "NO";
    CCU2C add_3660_17 (.A0(phase_inc_carrGen[14]), .B0(n17820), .C0(n18053), 
          .D0(led_c_2), .A1(n18053), .B1(n17820), .C1(phase_inc_carrGen[15]), 
          .D1(VCC_net), .CIN(n16414), .COUT(n16415), .S0(n281), .S1(n278));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_17.INIT0 = 16'h596a;
    defparam add_3660_17.INIT1 = 16'h4b4b;
    defparam add_3660_17.INJECT1_0 = "NO";
    defparam add_3660_17.INJECT1_1 = "NO";
    CCU2C add_3660_15 (.A0(phase_inc_carrGen[12]), .B0(n17820), .C0(n18053), 
          .D0(led_c_2), .A1(phase_inc_carrGen[13]), .B1(n17820), .C1(n18053), 
          .D1(n3674), .CIN(n16413), .COUT(n16414), .S0(n287), .S1(n284));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_15.INIT0 = 16'h596a;
    defparam add_3660_15.INIT1 = 16'h596a;
    defparam add_3660_15.INJECT1_0 = "NO";
    defparam add_3660_15.INJECT1_1 = "NO";
    CCU2C add_3660_13 (.A0(phase_inc_carrGen[10]), .B0(n17820), .C0(n18053), 
          .D0(n3674), .A1(phase_inc_carrGen[11]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16412), .COUT(n16413), .S0(n293), .S1(n290));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_13.INIT0 = 16'h596a;
    defparam add_3660_13.INIT1 = 16'haa6a;
    defparam add_3660_13.INJECT1_0 = "NO";
    defparam add_3660_13.INJECT1_1 = "NO";
    CCU2C add_3660_11 (.A0(n18053), .B0(n17820), .C0(phase_inc_carrGen[8]), 
          .D0(VCC_net), .A1(phase_inc_carrGen[9]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16411), .COUT(n16412), .S0(n299), .S1(n296));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_11.INIT0 = 16'h8787;
    defparam add_3660_11.INIT1 = 16'h6aaa;
    defparam add_3660_11.INJECT1_0 = "NO";
    defparam add_3660_11.INJECT1_1 = "NO";
    CCU2C add_3660_9 (.A0(n18053), .B0(n17820), .C0(phase_inc_carrGen[6]), 
          .D0(VCC_net), .A1(phase_inc_carrGen[7]), .B1(n17825), .C1(n12424), 
          .D1(n18053), .CIN(n16410), .COUT(n16411), .S0(n305), .S1(n302));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_9.INIT0 = 16'h4b4b;
    defparam add_3660_9.INIT1 = 16'h6aaa;
    defparam add_3660_9.INJECT1_0 = "NO";
    defparam add_3660_9.INJECT1_1 = "NO";
    CCU2C add_3660_7 (.A0(n18053), .B0(n17820), .C0(phase_inc_carrGen[4]), 
          .D0(VCC_net), .A1(n18053), .B1(n17820), .C1(phase_inc_carrGen[5]), 
          .D1(VCC_net), .CIN(n16409), .COUT(n16410), .S0(n311), .S1(n308));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_7.INIT0 = 16'h4b4b;
    defparam add_3660_7.INIT1 = 16'h4b4b;
    defparam add_3660_7.INJECT1_0 = "NO";
    defparam add_3660_7.INJECT1_1 = "NO";
    CCU2C add_3660_5 (.A0(n3728), .B0(phase_inc_carrGen[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(n3728), .B1(phase_inc_carrGen[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16408), .COUT(n16409), .S0(n317), .S1(n314));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_5.INIT0 = 16'h9995;
    defparam add_3660_5.INIT1 = 16'h9995;
    defparam add_3660_5.INJECT1_0 = "NO";
    defparam add_3660_5.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_2810), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16044));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1454_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1454_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_1.INJECT1_1 = "NO";
    CCU2C add_3660_3 (.A0(phase_inc_carrGen[0]), .B0(n17825), .C0(n12424), 
          .D0(n18053), .A1(phase_inc_carrGen[1]), .B1(n17820), .C1(n18053), 
          .D1(n3674), .CIN(n16407), .COUT(n16408), .S0(n323), .S1(n320));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_3.INIT0 = 16'h6aaa;
    defparam add_3660_3.INIT1 = 16'h596a;
    defparam add_3660_3.INJECT1_0 = "NO";
    defparam add_3660_3.INJECT1_1 = "NO";
    CCU2C add_3660_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n17827), .B1(n18096), .C1(n12424), .D1(led_c_4), .COUT(n16407));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam add_3660_1.INIT0 = 16'h0000;
    defparam add_3660_1.INIT1 = 16'hff7f;
    defparam add_3660_1.INJECT1_0 = "NO";
    defparam add_3660_1.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_38 (.A0(d2_adj_5711[71]), .B0(d1_adj_5710[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16040), .S0(n78_adj_5608));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1544_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_38.INJECT1_1 = "NO";
    CCU2C add_3658_17 (.A0(d_out_d_11__N_1877), .B0(d_out_d_11__N_1878[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1877), .B1(d_out_d_11__N_1878[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16402), .S0(n41_adj_4837), 
          .S1(d_out_d_11__N_1880[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3658_17.INIT0 = 16'h666a;
    defparam add_3658_17.INIT1 = 16'h666a;
    defparam add_3658_17.INJECT1_0 = "NO";
    defparam add_3658_17.INJECT1_1 = "NO";
    CCU2C add_3658_15 (.A0(d_out_d_11__N_1878[17]), .B0(n40), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n37_adj_5681), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16401), .COUT(n16402), .S0(n47_adj_4839), 
          .S1(n44_adj_4838));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3658_15.INIT0 = 16'h9995;
    defparam add_3658_15.INIT1 = 16'h9995;
    defparam add_3658_15.INJECT1_0 = "NO";
    defparam add_3658_15.INJECT1_1 = "NO";
    CCU2C add_3658_13 (.A0(d_out_d_11__N_1878[17]), .B0(n46), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n43), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16400), .COUT(n16401), .S0(n53), .S1(n50_adj_4840));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3658_13.INIT0 = 16'h9995;
    defparam add_3658_13.INIT1 = 16'h9995;
    defparam add_3658_13.INJECT1_0 = "NO";
    defparam add_3658_13.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_32 (.A0(d_d6[65]), .B0(d6[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[66]), .B1(d6[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16243), .COUT(n16244), .S0(n96_adj_5471), .S1(n93_adj_5470));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_32.INJECT1_1 = "NO";
    CCU2C add_3658_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1878[17]), .C0(n52), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1878[17]), 
          .C1(n49), .D1(VCC_net), .CIN(n16399), .COUT(n16400), .S0(n59), 
          .S1(n56));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3658_11.INIT0 = 16'h6969;
    defparam add_3658_11.INIT1 = 16'h6969;
    defparam add_3658_11.INJECT1_0 = "NO";
    defparam add_3658_11.INJECT1_1 = "NO";
    CCU2C add_3658_9 (.A0(d_out_d_11__N_1878[17]), .B0(n58), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1878[17]), 
          .C1(n55), .D1(VCC_net), .CIN(n16398), .COUT(n16399), .S0(n65_adj_4841), 
          .S1(n62));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3658_9.INIT0 = 16'h9995;
    defparam add_3658_9.INIT1 = 16'h6969;
    defparam add_3658_9.INJECT1_0 = "NO";
    defparam add_3658_9.INJECT1_1 = "NO";
    CCU2C add_3658_7 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1878[17]), 
          .C0(n64), .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n17826), 
          .C1(n61), .D1(VCC_net), .CIN(n16397), .COUT(n16398), .S0(n71), 
          .S1(n68));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3658_7.INIT0 = 16'h9696;
    defparam add_3658_7.INIT1 = 16'h6969;
    defparam add_3658_7.INJECT1_0 = "NO";
    defparam add_3658_7.INJECT1_1 = "NO";
    CCU2C add_3658_5 (.A0(n70), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1876[17]), .B1(d_out_d_11__N_1878[17]), .C1(n67), 
          .D1(VCC_net), .CIN(n16396), .COUT(n16397), .S0(n77), .S1(n74));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3658_5.INIT0 = 16'haaa0;
    defparam add_3658_5.INIT1 = 16'h9696;
    defparam add_3658_5.INJECT1_0 = "NO";
    defparam add_3658_5.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_24 (.A0(d5_adj_5714[57]), .B0(d4_adj_5713[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[58]), .B1(d4_adj_5713[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16163), .COUT(n16164), .S0(n120_adj_5552), 
          .S1(n117_adj_5551));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_30 (.A0(d_d6[63]), .B0(d6[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[64]), .B1(d6[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16242), .COUT(n16243), .S0(n102_adj_5473), .S1(n99_adj_5472));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_30.INJECT1_1 = "NO";
    CCU2C add_3658_3 (.A0(d_out_d_11__N_1878[17]), .B0(ISquare[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16395), .COUT(n16396), .S1(n80));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3658_3.INIT0 = 16'h666a;
    defparam add_3658_3.INIT1 = 16'h555f;
    defparam add_3658_3.INJECT1_0 = "NO";
    defparam add_3658_3.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_28 (.A0(d_d6[61]), .B0(d6[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[62]), .B1(d6[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16241), .COUT(n16242), .S0(n108_adj_5475), .S1(n105_adj_5474));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_28.INJECT1_1 = "NO";
    CCU2C add_3658_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1878[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16395));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3658_1.INIT0 = 16'h0000;
    defparam add_3658_1.INIT1 = 16'haaaf;
    defparam add_3658_1.INJECT1_0 = "NO";
    defparam add_3658_1.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_6 (.A0(d_d_tmp[39]), .B0(d_tmp[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[40]), .B1(d_tmp[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16194), .COUT(n16195), .S0(n174_adj_5534), 
          .S1(n171_adj_5533));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_27 (.A0(d4[60]), .B0(cout_adj_2810), .C0(n111_adj_5296), 
          .D0(d5[60]), .A1(d4[61]), .B1(cout_adj_2810), .C1(n108_adj_5295), 
          .D1(d5[61]), .CIN(n16056), .COUT(n16057), .S0(d5_71__N_706[60]), 
          .S1(d5_71__N_706[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_27.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_78 (.A(led_c_0), .B(led_c_2), .Z(n16867)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_78.init = 16'h2222;
    CCU2C _add_1_1553_add_4_22 (.A0(d5_adj_5714[55]), .B0(d4_adj_5713[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[56]), .B1(d4_adj_5713[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16162), .COUT(n16163), .S0(n126_adj_5554), 
          .S1(n123_adj_5553));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_11 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n159_adj_5109), .D0(d1[44]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n156_adj_5108), .D1(d1[45]), .CIN(n15701), .COUT(n15702), 
          .S0(d1_71__N_418[44]), .S1(d1_71__N_418[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_11.INJECT1_1 = "NO";
    CCU2C add_3657_19 (.A0(d_out_d_11__N_1888[17]), .B0(n48_adj_5683), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n45_adj_5682), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16389), .S0(n45_adj_5445), 
          .S1(d_out_d_11__N_1890[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3657_19.INIT0 = 16'h9995;
    defparam add_3657_19.INIT1 = 16'h9995;
    defparam add_3657_19.INJECT1_0 = "NO";
    defparam add_3657_19.INJECT1_1 = "NO";
    CCU2C add_3657_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1888[17]), .C0(n54_adj_5685), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n51_adj_5684), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16388), .COUT(n16389), .S0(n51_adj_5447), 
          .S1(n48_adj_5446));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3657_17.INIT0 = 16'h6969;
    defparam add_3657_17.INIT1 = 16'h9995;
    defparam add_3657_17.INJECT1_0 = "NO";
    defparam add_3657_17.INJECT1_1 = "NO";
    CCU2C add_3657_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1888[17]), .C0(n60_adj_5687), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1888[17]), 
          .C1(n57_adj_5686), .D1(VCC_net), .CIN(n16387), .COUT(n16388), 
          .S0(n57_adj_5449), .S1(n54_adj_5448));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3657_15.INIT0 = 16'h6969;
    defparam add_3657_15.INIT1 = 16'h6969;
    defparam add_3657_15.INJECT1_0 = "NO";
    defparam add_3657_15.INJECT1_1 = "NO";
    CCU2C add_3657_13 (.A0(d_out_d_11__N_1888[17]), .B0(n17826), .C0(n66_adj_5689), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n63_adj_5688), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16386), .COUT(n16387), .S0(n63_adj_5451), 
          .S1(n60_adj_5450));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3657_13.INIT0 = 16'h6969;
    defparam add_3657_13.INIT1 = 16'h9995;
    defparam add_3657_13.INJECT1_0 = "NO";
    defparam add_3657_13.INJECT1_1 = "NO";
    CCU2C add_3657_11 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(n72_adj_5691), .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(n69_adj_5690), .D1(VCC_net), 
          .CIN(n16385), .COUT(n16386), .S0(n69_adj_5453), .S1(n66_adj_5452));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3657_11.INIT0 = 16'h9696;
    defparam add_3657_11.INIT1 = 16'h9696;
    defparam add_3657_11.INJECT1_0 = "NO";
    defparam add_3657_11.INJECT1_1 = "NO";
    CCU2C add_3657_9 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(n78_adj_5693), .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(n75_adj_5692), .D1(VCC_net), 
          .CIN(n16384), .COUT(n16385), .S0(n75_adj_5455), .S1(n72_adj_5454));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3657_9.INIT0 = 16'h9696;
    defparam add_3657_9.INIT1 = 16'h9696;
    defparam add_3657_9.INJECT1_0 = "NO";
    defparam add_3657_9.INJECT1_1 = "NO";
    CCU2C add_3657_7 (.A0(d_out_d_11__N_1884[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(n84_adj_5695), .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(n81_adj_5694), .D1(VCC_net), 
          .CIN(n16383), .COUT(n16384), .S0(n81_adj_5457), .S1(n78_adj_5456));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3657_7.INIT0 = 16'h9696;
    defparam add_3657_7.INIT1 = 16'h9696;
    defparam add_3657_7.INJECT1_0 = "NO";
    defparam add_3657_7.INJECT1_1 = "NO";
    CCU2C add_3657_5 (.A0(n90_adj_5697), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1886[17]), .B1(d_out_d_11__N_1888[17]), .C1(n87_adj_5696), 
          .D1(VCC_net), .CIN(n16382), .COUT(n16383), .S0(n87_adj_5459), 
          .S1(n84_adj_5458));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3657_5.INIT0 = 16'haaa0;
    defparam add_3657_5.INIT1 = 16'h9696;
    defparam add_3657_5.INJECT1_0 = "NO";
    defparam add_3657_5.INJECT1_1 = "NO";
    CCU2C add_3657_3 (.A0(d_out_d_11__N_1888[17]), .B0(ISquare[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16381), .COUT(n16382), .S1(n90_adj_5460));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3657_3.INIT0 = 16'h666a;
    defparam add_3657_3.INIT1 = 16'h555f;
    defparam add_3657_3.INJECT1_0 = "NO";
    defparam add_3657_3.INJECT1_1 = "NO";
    CCU2C add_3657_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1888[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16381));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3657_1.INIT0 = 16'h0000;
    defparam add_3657_1.INIT1 = 16'haaaf;
    defparam add_3657_1.INJECT1_0 = "NO";
    defparam add_3657_1.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_9 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n165_adj_5111), .D0(d1[42]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n162_adj_5110), .D1(d1[43]), .CIN(n15700), .COUT(n15701), 
          .S0(d1_71__N_418[42]), .S1(d1_71__N_418[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_9.INJECT1_1 = "NO";
    CCU2C add_3659_13 (.A0(d_out_d_11__N_1873), .B0(d_out_d_11__N_1874[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1873), .B1(d_out_d_11__N_1874[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16375), .S0(n33_adj_2796), 
          .S1(d_out_d_11__N_1876[17]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3659_13.INIT0 = 16'h666a;
    defparam add_3659_13.INIT1 = 16'h666a;
    defparam add_3659_13.INJECT1_0 = "NO";
    defparam add_3659_13.INJECT1_1 = "NO";
    CCU2C add_3659_11 (.A0(d_out_d_11__N_1874[17]), .B0(n32_adj_4743), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), .B1(n29_adj_4752), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16374), .COUT(n16375), .S0(n39), 
          .S1(n36_adj_2795));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3659_11.INIT0 = 16'h9995;
    defparam add_3659_11.INIT1 = 16'h9995;
    defparam add_3659_11.INJECT1_0 = "NO";
    defparam add_3659_11.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_12 (.A0(d2_adj_5711[45]), .B0(d1_adj_5710[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[46]), .B1(d1_adj_5710[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16027), .COUT(n16028), .S0(n156_adj_5634), 
          .S1(n153_adj_5633));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_7 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n171_adj_5113), .D0(d1[40]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n168_adj_5112), .D1(d1[41]), .CIN(n15699), .COUT(n15700), 
          .S0(d1_71__N_418[40]), .S1(d1_71__N_418[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_5 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n177_adj_5115), .D0(d1[38]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n174_adj_5114), .D1(d1[39]), .CIN(n15698), .COUT(n15699), 
          .S0(d1_71__N_418[38]), .S1(d1_71__N_418[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_3 (.A0(MixerOutSin[11]), .B0(cout_adj_5021), 
          .C0(n183_adj_5117), .D0(d1[36]), .A1(MixerOutSin[11]), .B1(cout_adj_5021), 
          .C1(n180_adj_5116), .D1(d1[37]), .CIN(n15697), .COUT(n15698), 
          .S0(d1_71__N_418[36]), .S1(d1_71__N_418[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1397_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1397_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1397_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5021), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15697));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1397_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1397_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1397_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1397_add_4_1.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_26 (.A0(MultResult2[23]), .B0(MultResult1[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15693), .S0(n54_adj_5224));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_26.INIT0 = 16'h666a;
    defparam ISquare_add_4_26.INIT1 = 16'h0000;
    defparam ISquare_add_4_26.INJECT1_0 = "NO";
    defparam ISquare_add_4_26.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_24 (.A0(MultResult2[22]), .B0(MultResult1[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[23]), .B1(MultResult1[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15692), .COUT(n15693), .S0(n60_adj_5226), 
          .S1(n57_adj_5225));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_24.INIT0 = 16'h666a;
    defparam ISquare_add_4_24.INIT1 = 16'h666a;
    defparam ISquare_add_4_24.INJECT1_0 = "NO";
    defparam ISquare_add_4_24.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_22 (.A0(MultResult2[20]), .B0(MultResult1[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[21]), .B1(MultResult1[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15691), .COUT(n15692), .S0(n66_adj_5228), 
          .S1(n63_adj_5227));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_22.INIT0 = 16'h666a;
    defparam ISquare_add_4_22.INIT1 = 16'h666a;
    defparam ISquare_add_4_22.INJECT1_0 = "NO";
    defparam ISquare_add_4_22.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_20 (.A0(MultResult2[18]), .B0(MultResult1[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[19]), .B1(MultResult1[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15690), .COUT(n15691), .S0(n72_adj_5230), 
          .S1(n69_adj_5229));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_20.INIT0 = 16'h666a;
    defparam ISquare_add_4_20.INIT1 = 16'h666a;
    defparam ISquare_add_4_20.INJECT1_0 = "NO";
    defparam ISquare_add_4_20.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_18 (.A0(MultResult2[16]), .B0(MultResult1[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[17]), .B1(MultResult1[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15689), .COUT(n15690), .S0(n78_adj_5232), 
          .S1(n75_adj_5231));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_18.INIT0 = 16'h666a;
    defparam ISquare_add_4_18.INIT1 = 16'h666a;
    defparam ISquare_add_4_18.INJECT1_0 = "NO";
    defparam ISquare_add_4_18.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_16 (.A0(MultResult2[14]), .B0(MultResult1[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[15]), .B1(MultResult1[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15688), .COUT(n15689), .S0(n84_adj_5234), 
          .S1(n81_adj_5233));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_16.INIT0 = 16'h666a;
    defparam ISquare_add_4_16.INIT1 = 16'h666a;
    defparam ISquare_add_4_16.INJECT1_0 = "NO";
    defparam ISquare_add_4_16.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_14 (.A0(MultResult2[12]), .B0(MultResult1[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[13]), .B1(MultResult1[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15687), .COUT(n15688), .S0(n90_adj_5236), 
          .S1(n87_adj_5235));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_14.INIT0 = 16'h666a;
    defparam ISquare_add_4_14.INIT1 = 16'h666a;
    defparam ISquare_add_4_14.INJECT1_0 = "NO";
    defparam ISquare_add_4_14.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_12 (.A0(MultResult2[10]), .B0(MultResult1[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[11]), .B1(MultResult1[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15686), .COUT(n15687), .S0(n96_adj_5238), 
          .S1(n93_adj_5237));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_12.INIT0 = 16'h666a;
    defparam ISquare_add_4_12.INIT1 = 16'h666a;
    defparam ISquare_add_4_12.INJECT1_0 = "NO";
    defparam ISquare_add_4_12.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_10 (.A0(MultResult2[8]), .B0(MultResult1[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[9]), .B1(MultResult1[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15685), .COUT(n15686), .S0(n102_adj_5240), 
          .S1(n99_adj_5239));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_10.INIT0 = 16'h666a;
    defparam ISquare_add_4_10.INIT1 = 16'h666a;
    defparam ISquare_add_4_10.INJECT1_0 = "NO";
    defparam ISquare_add_4_10.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_8 (.A0(MultResult2[6]), .B0(MultResult1[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[7]), .B1(MultResult1[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15684), .COUT(n15685), .S0(n108_adj_5242), 
          .S1(n105_adj_5241));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_8.INIT0 = 16'h666a;
    defparam ISquare_add_4_8.INIT1 = 16'h666a;
    defparam ISquare_add_4_8.INJECT1_0 = "NO";
    defparam ISquare_add_4_8.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_6 (.A0(MultResult2[4]), .B0(MultResult1[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[5]), .B1(MultResult1[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15683), .COUT(n15684), .S0(n114_adj_5244), 
          .S1(n111_adj_5243));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_6.INIT0 = 16'h666a;
    defparam ISquare_add_4_6.INIT1 = 16'h666a;
    defparam ISquare_add_4_6.INJECT1_0 = "NO";
    defparam ISquare_add_4_6.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_4 (.A0(MultResult2[2]), .B0(MultResult1[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[3]), .B1(MultResult1[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15682), .COUT(n15683), .S0(n120_adj_5246), 
          .S1(n117_adj_5245));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_4.INIT0 = 16'h666a;
    defparam ISquare_add_4_4.INIT1 = 16'h666a;
    defparam ISquare_add_4_4.INJECT1_0 = "NO";
    defparam ISquare_add_4_4.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_2 (.A0(MultResult2[0]), .B0(MultResult1[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[1]), .B1(MultResult1[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15682), .S1(n123_adj_5247));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_2.INIT0 = 16'h0008;
    defparam ISquare_add_4_2.INIT1 = 16'h666a;
    defparam ISquare_add_4_2.INJECT1_0 = "NO";
    defparam ISquare_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_37 (.A0(d6[70]), .B0(cout_adj_5644), .C0(n81_adj_5466), 
          .D0(n3_adj_4688), .A1(d6[71]), .B1(cout_adj_5644), .C1(n78_adj_5465), 
          .D1(n2_adj_4689), .CIN(n15679), .S0(d7_71__N_1531[70]), .S1(d7_71__N_1531[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_35 (.A0(d6[68]), .B0(cout_adj_5644), .C0(n87_adj_5468), 
          .D0(n5_adj_4686), .A1(d6[69]), .B1(cout_adj_5644), .C1(n84_adj_5467), 
          .D1(n4_adj_4687), .CIN(n15678), .COUT(n15679), .S0(d7_71__N_1531[68]), 
          .S1(d7_71__N_1531[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_33 (.A0(d6[66]), .B0(cout_adj_5644), .C0(n93_adj_5470), 
          .D0(n7_adj_4684), .A1(d6[67]), .B1(cout_adj_5644), .C1(n90_adj_5469), 
          .D1(n6_adj_4685), .CIN(n15677), .COUT(n15678), .S0(d7_71__N_1531[66]), 
          .S1(d7_71__N_1531[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_31 (.A0(d6[64]), .B0(cout_adj_5644), .C0(n99_adj_5472), 
          .D0(n9_adj_4682), .A1(d6[65]), .B1(cout_adj_5644), .C1(n96_adj_5471), 
          .D1(n8_adj_4683), .CIN(n15676), .COUT(n15677), .S0(d7_71__N_1531[64]), 
          .S1(d7_71__N_1531[65]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_29 (.A0(d6[62]), .B0(cout_adj_5644), .C0(n105_adj_5474), 
          .D0(n11_adj_4680), .A1(d6[63]), .B1(cout_adj_5644), .C1(n102_adj_5473), 
          .D1(n10_adj_4681), .CIN(n15675), .COUT(n15676), .S0(d7_71__N_1531[62]), 
          .S1(d7_71__N_1531[63]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_27 (.A0(d6[60]), .B0(cout_adj_5644), .C0(n111_adj_5476), 
          .D0(n13_adj_4678), .A1(d6[61]), .B1(cout_adj_5644), .C1(n108_adj_5475), 
          .D1(n12_adj_4679), .CIN(n15674), .COUT(n15675), .S0(d7_71__N_1531[60]), 
          .S1(d7_71__N_1531[61]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_25 (.A0(d6[58]), .B0(cout_adj_5644), .C0(n117_adj_5478), 
          .D0(n15_adj_4676), .A1(d6[59]), .B1(cout_adj_5644), .C1(n114_adj_5477), 
          .D1(n14_adj_4677), .CIN(n15673), .COUT(n15674), .S0(d7_71__N_1531[58]), 
          .S1(d7_71__N_1531[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_23 (.A0(d6[56]), .B0(cout_adj_5644), .C0(n123_adj_5480), 
          .D0(n17_adj_4674), .A1(d6[57]), .B1(cout_adj_5644), .C1(n120_adj_5479), 
          .D1(n16_adj_4675), .CIN(n15672), .COUT(n15673), .S0(d7_71__N_1531[56]), 
          .S1(d7_71__N_1531[57]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_21 (.A0(d6[54]), .B0(cout_adj_5644), .C0(n129_adj_5482), 
          .D0(n19_adj_4672), .A1(d6[55]), .B1(cout_adj_5644), .C1(n126_adj_5481), 
          .D1(n18_adj_4673), .CIN(n15671), .COUT(n15672), .S0(d7_71__N_1531[54]), 
          .S1(d7_71__N_1531[55]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_19 (.A0(d6[52]), .B0(cout_adj_5644), .C0(n135_adj_5484), 
          .D0(n21_adj_4670), .A1(d6[53]), .B1(cout_adj_5644), .C1(n132_adj_5483), 
          .D1(n20_adj_4671), .CIN(n15670), .COUT(n15671), .S0(d7_71__N_1531[52]), 
          .S1(d7_71__N_1531[53]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_17 (.A0(d6[50]), .B0(cout_adj_5644), .C0(n141_adj_5486), 
          .D0(n23_adj_4668), .A1(d6[51]), .B1(cout_adj_5644), .C1(n138_adj_5485), 
          .D1(n22_adj_4669), .CIN(n15669), .COUT(n15670), .S0(d7_71__N_1531[50]), 
          .S1(d7_71__N_1531[51]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_15 (.A0(d6[48]), .B0(cout_adj_5644), .C0(n147_adj_5488), 
          .D0(n25_adj_4666), .A1(d6[49]), .B1(cout_adj_5644), .C1(n144_adj_5487), 
          .D1(n24_adj_4667), .CIN(n15668), .COUT(n15669), .S0(d7_71__N_1531[48]), 
          .S1(d7_71__N_1531[49]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_13 (.A0(d6[46]), .B0(cout_adj_5644), .C0(n153_adj_5490), 
          .D0(n27_adj_4664), .A1(d6[47]), .B1(cout_adj_5644), .C1(n150_adj_5489), 
          .D1(n26_adj_4665), .CIN(n15667), .COUT(n15668), .S0(d7_71__N_1531[46]), 
          .S1(d7_71__N_1531[47]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_11 (.A0(d6[44]), .B0(cout_adj_5644), .C0(n159_adj_5492), 
          .D0(n29_adj_4662), .A1(d6[45]), .B1(cout_adj_5644), .C1(n156_adj_5491), 
          .D1(n28_adj_4663), .CIN(n15666), .COUT(n15667), .S0(d7_71__N_1531[44]), 
          .S1(d7_71__N_1531[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_9 (.A0(d6[42]), .B0(cout_adj_5644), .C0(n165_adj_5494), 
          .D0(n31_adj_4660), .A1(d6[43]), .B1(cout_adj_5644), .C1(n162_adj_5493), 
          .D1(n30_adj_4661), .CIN(n15665), .COUT(n15666), .S0(d7_71__N_1531[42]), 
          .S1(d7_71__N_1531[43]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_7 (.A0(d6[40]), .B0(cout_adj_5644), .C0(n171_adj_5496), 
          .D0(n33_adj_4658), .A1(d6[41]), .B1(cout_adj_5644), .C1(n168_adj_5495), 
          .D1(n32_adj_4659), .CIN(n15664), .COUT(n15665), .S0(d7_71__N_1531[40]), 
          .S1(d7_71__N_1531[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_5 (.A0(d6[38]), .B0(cout_adj_5644), .C0(n177_adj_5498), 
          .D0(n35_adj_4656), .A1(d6[39]), .B1(cout_adj_5644), .C1(n174_adj_5497), 
          .D1(n34_adj_4657), .CIN(n15663), .COUT(n15664), .S0(d7_71__N_1531[38]), 
          .S1(d7_71__N_1531[39]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_3 (.A0(d6[36]), .B0(cout_adj_5644), .C0(n183_adj_5500), 
          .D0(n37_adj_4654), .A1(d6[37]), .B1(cout_adj_5644), .C1(n180_adj_5499), 
          .D1(n36_adj_4655), .CIN(n15662), .COUT(n15663), .S0(d7_71__N_1531[36]), 
          .S1(d7_71__N_1531[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1433_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1433_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5644), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15662));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1433_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1433_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1433_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_38 (.A0(d_d8_adj_5720[71]), .B0(d8_adj_5719[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15658), .S0(n78_adj_4950));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1592_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_36 (.A0(d_d8_adj_5720[69]), .B0(d8_adj_5719[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[70]), .B1(d8_adj_5719[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15657), .COUT(n15658), .S0(n84_adj_4952), 
          .S1(n81_adj_4951));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_34 (.A0(d_d8_adj_5720[67]), .B0(d8_adj_5719[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[68]), .B1(d8_adj_5719[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15656), .COUT(n15657), .S0(n90_adj_4954), 
          .S1(n87_adj_4953));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_32 (.A0(d_d8_adj_5720[65]), .B0(d8_adj_5719[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[66]), .B1(d8_adj_5719[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15655), .COUT(n15656), .S0(n96_adj_4956), 
          .S1(n93_adj_4955));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_30 (.A0(d_d8_adj_5720[63]), .B0(d8_adj_5719[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[64]), .B1(d8_adj_5719[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15654), .COUT(n15655), .S0(n102_adj_4958), 
          .S1(n99_adj_4957));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_28 (.A0(d_d8_adj_5720[61]), .B0(d8_adj_5719[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[62]), .B1(d8_adj_5719[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15653), .COUT(n15654), .S0(n108_adj_4960), 
          .S1(n105_adj_4959));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_26 (.A0(d_d8_adj_5720[59]), .B0(d8_adj_5719[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[60]), .B1(d8_adj_5719[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15652), .COUT(n15653), .S0(n114_adj_4962), 
          .S1(n111_adj_4961));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_24 (.A0(d_d8_adj_5720[57]), .B0(d8_adj_5719[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[58]), .B1(d8_adj_5719[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15651), .COUT(n15652), .S0(n120_adj_4964), 
          .S1(n117_adj_4963));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_22 (.A0(d_d8_adj_5720[55]), .B0(d8_adj_5719[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[56]), .B1(d8_adj_5719[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15650), .COUT(n15651), .S0(n126_adj_4966), 
          .S1(n123_adj_4965));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_20 (.A0(d_d8_adj_5720[53]), .B0(d8_adj_5719[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[54]), .B1(d8_adj_5719[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15649), .COUT(n15650), .S0(n132_adj_4968), 
          .S1(n129_adj_4967));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_18 (.A0(d_d8_adj_5720[51]), .B0(d8_adj_5719[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[52]), .B1(d8_adj_5719[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15648), .COUT(n15649), .S0(n138_adj_4970), 
          .S1(n135_adj_4969));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_16 (.A0(d_d8_adj_5720[49]), .B0(d8_adj_5719[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[50]), .B1(d8_adj_5719[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15647), .COUT(n15648), .S0(n144_adj_4972), 
          .S1(n141_adj_4971));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_14 (.A0(d_d8_adj_5720[47]), .B0(d8_adj_5719[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[48]), .B1(d8_adj_5719[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15646), .COUT(n15647), .S0(n150_adj_4974), 
          .S1(n147_adj_4973));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_12 (.A0(d_d8_adj_5720[45]), .B0(d8_adj_5719[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[46]), .B1(d8_adj_5719[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15645), .COUT(n15646), .S0(n156_adj_4976), 
          .S1(n153_adj_4975));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_10 (.A0(d_d8_adj_5720[43]), .B0(d8_adj_5719[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[44]), .B1(d8_adj_5719[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15644), .COUT(n15645), .S0(n162_adj_4978), 
          .S1(n159_adj_4977));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_8 (.A0(d_d8_adj_5720[41]), .B0(d8_adj_5719[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[42]), .B1(d8_adj_5719[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15643), .COUT(n15644), .S0(n168_adj_4980), 
          .S1(n165_adj_4979));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_6 (.A0(d_d8_adj_5720[39]), .B0(d8_adj_5719[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[40]), .B1(d8_adj_5719[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15642), .COUT(n15643), .S0(n174_adj_4982), 
          .S1(n171_adj_4981));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_4 (.A0(d_d8_adj_5720[37]), .B0(d8_adj_5719[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5720[38]), .B1(d8_adj_5719[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15641), .COUT(n15642), .S0(n180_adj_4984), 
          .S1(n177_adj_4983));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1592_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1592_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8_adj_5720[36]), .B1(d8_adj_5719[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15641), .S1(n183_adj_4985));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1592_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1592_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1592_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1592_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_38 (.A0(d_d9_adj_5722[71]), .B0(d9_adj_5721[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15640), .S0(n78_adj_4986));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1595_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_36 (.A0(d_d9_adj_5722[69]), .B0(d9_adj_5721[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[70]), .B1(d9_adj_5721[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15639), .COUT(n15640), .S0(n84_adj_4988), 
          .S1(n81_adj_4987));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_34 (.A0(d_d9_adj_5722[67]), .B0(d9_adj_5721[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[68]), .B1(d9_adj_5721[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15638), .COUT(n15639), .S0(n90_adj_4990), 
          .S1(n87_adj_4989));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_32 (.A0(d_d9_adj_5722[65]), .B0(d9_adj_5721[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[66]), .B1(d9_adj_5721[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15637), .COUT(n15638), .S0(n96_adj_4992), 
          .S1(n93_adj_4991));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_30 (.A0(d_d9_adj_5722[63]), .B0(d9_adj_5721[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[64]), .B1(d9_adj_5721[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15636), .COUT(n15637), .S0(n102_adj_4994), 
          .S1(n99_adj_4993));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_28 (.A0(d_d9_adj_5722[61]), .B0(d9_adj_5721[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[62]), .B1(d9_adj_5721[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15635), .COUT(n15636), .S0(n108_adj_4996), 
          .S1(n105_adj_4995));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_26 (.A0(d_d9_adj_5722[59]), .B0(d9_adj_5721[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[60]), .B1(d9_adj_5721[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15634), .COUT(n15635), .S0(n114_adj_4998), 
          .S1(n111_adj_4997));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_24 (.A0(d_d9_adj_5722[57]), .B0(d9_adj_5721[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[58]), .B1(d9_adj_5721[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15633), .COUT(n15634), .S0(n120_adj_5000), 
          .S1(n117_adj_4999));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_22 (.A0(d_d9_adj_5722[55]), .B0(d9_adj_5721[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[56]), .B1(d9_adj_5721[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15632), .COUT(n15633));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_20 (.A0(d_d9_adj_5722[53]), .B0(d9_adj_5721[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[54]), .B1(d9_adj_5721[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15631), .COUT(n15632));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_18 (.A0(d_d9_adj_5722[51]), .B0(d9_adj_5721[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[52]), .B1(d9_adj_5721[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15630), .COUT(n15631));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_16 (.A0(d_d9_adj_5722[49]), .B0(d9_adj_5721[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[50]), .B1(d9_adj_5721[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15629), .COUT(n15630));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_14 (.A0(d_d9_adj_5722[47]), .B0(d9_adj_5721[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[48]), .B1(d9_adj_5721[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15628), .COUT(n15629));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_12 (.A0(d_d9_adj_5722[45]), .B0(d9_adj_5721[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[46]), .B1(d9_adj_5721[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15627), .COUT(n15628));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_10 (.A0(d_d9_adj_5722[43]), .B0(d9_adj_5721[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[44]), .B1(d9_adj_5721[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15626), .COUT(n15627));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_8 (.A0(d_d9_adj_5722[41]), .B0(d9_adj_5721[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[42]), .B1(d9_adj_5721[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15625), .COUT(n15626));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_6 (.A0(d_d9_adj_5722[39]), .B0(d9_adj_5721[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[40]), .B1(d9_adj_5721[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15624), .COUT(n15625));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_4 (.A0(d_d9_adj_5722[37]), .B0(d9_adj_5721[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5722[38]), .B1(d9_adj_5721[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15623), .COUT(n15624));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1595_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1595_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9_adj_5722[36]), .B1(d9_adj_5721[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15623));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1595_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1595_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1595_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1595_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1601_add_4_38 (.A0(d_d_tmp[35]), .B0(d_tmp[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15622), .S0(d6_71__N_1459[35]), .S1(cout_adj_5001));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1601_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1601_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1601_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1601_add_4_38.INJECT1_1 = "NO";
    LUT4 i3178_4_lut_4_lut (.A(led_c_4), .B(n17817), .C(n205), .D(n199_adj_5047), 
         .Z(n2607)) /* synthesis lut_function=(A (C)+!A !(B+!(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3178_4_lut_4_lut.init = 16'hb1a0;
    LUT4 i5964_4_lut (.A(n16829), .B(led_c_1), .C(n17832), .D(led_c_0), 
         .Z(n16842)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i5964_4_lut.init = 16'h0040;
    LUT4 i2357_3_lut (.A(led_c_1), .B(n160), .C(n18053), .Z(n12260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2357_3_lut.init = 16'hcaca;
    LUT4 i2355_3_lut (.A(led_c_1), .B(n175), .C(led_c_4), .Z(n12258)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2355_3_lut.init = 16'hc5c5;
    LUT4 i2353_3_lut (.A(led_c_1), .B(n199), .C(led_c_4), .Z(n12256)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2353_3_lut.init = 16'hc5c5;
    LUT4 i2690_3_lut (.A(n188), .B(n2668), .C(n12538), .Z(n12595)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2690_3_lut.init = 16'hacac;
    LUT4 mux_339_i46_4_lut (.A(n3906), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2668)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i46_4_lut.init = 16'hc0ca;
    LUT4 mux_843_i45_3_lut (.A(n178_adj_5040), .B(n184), .C(led_c_4), 
         .Z(n3906)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i45_3_lut.init = 16'hcaca;
    LUT4 i2706_4_lut (.A(n158), .B(n12007), .C(n12538), .D(n17813), 
         .Z(n12611)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2706_4_lut.init = 16'hafac;
    LUT4 i3162_4_lut_4_lut (.A(led_c_4), .B(n17817), .C(n307), .D(n301_adj_5081), 
         .Z(n2641)) /* synthesis lut_function=(A (C)+!A !(B+!(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3162_4_lut_4_lut.init = 16'hb1a0;
    LUT4 i3179_4_lut_4_lut (.A(n18053), .B(n17817), .C(n202), .D(n196_adj_5046), 
         .Z(n2606)) /* synthesis lut_function=(A (C)+!A !(B+!(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3179_4_lut_4_lut.init = 16'hb1a0;
    LUT4 mux_843_i31_3_lut (.A(n220_adj_5054), .B(n226), .C(n18053), .Z(n3920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i31_3_lut.init = 16'hcaca;
    LUT4 i2113_3_lut (.A(n12006), .B(n154), .C(n18053), .Z(n12007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2113_3_lut.init = 16'hcaca;
    LUT4 i2672_3_lut (.A(n236), .B(n2684), .C(n12538), .Z(n12577)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2672_3_lut.init = 16'hacac;
    LUT4 mux_339_i30_4_lut (.A(n3922), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i30_4_lut.init = 16'hcfca;
    LUT4 i5065_2_lut (.A(d2_adj_5711[0]), .B(d1_adj_5710[0]), .Z(d2_71__N_490_adj_5727[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5065_2_lut.init = 16'h6666;
    LUT4 i5064_2_lut (.A(d3_adj_5712[0]), .B(d2_adj_5711[0]), .Z(d3_71__N_562_adj_5728[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5064_2_lut.init = 16'h6666;
    LUT4 i5045_2_lut (.A(d4[0]), .B(d3[0]), .Z(d4_71__N_634[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5045_2_lut.init = 16'h6666;
    LUT4 mux_843_i29_3_lut (.A(n226_adj_5056), .B(n232), .C(n18053), .Z(n3922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i29_3_lut.init = 16'hcaca;
    LUT4 i5044_2_lut (.A(d5[0]), .B(d4[0]), .Z(d5_71__N_706[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5044_2_lut.init = 16'h6666;
    LUT4 i2704_3_lut (.A(n161), .B(n2659), .C(n12538), .Z(n12609)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2704_3_lut.init = 16'hacac;
    LUT4 mux_339_i55_4_lut (.A(n3897), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2659)) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i55_4_lut.init = 16'h3f3a;
    LUT4 i2090_3_lut_4_lut (.A(n17823), .B(n16869), .C(led_c_0), .D(n232_adj_5058), 
         .Z(n11984)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i2090_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_843_i54_3_lut (.A(n151_adj_5031), .B(n157), .C(led_c_4), 
         .Z(n3897)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i54_3_lut.init = 16'hcaca;
    LUT4 i2070_3_lut_4_lut (.A(n17823), .B(n16869), .C(led_c_0), .D(n292_adj_5078), 
         .Z(n11964)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i2070_3_lut_4_lut.init = 16'hf780;
    LUT4 i2670_4_lut (.A(n239), .B(n2617), .C(n12538), .D(n17813), .Z(n12575)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2670_4_lut.init = 16'hafac;
    LUT4 i2664_4_lut (.A(n254), .B(n2622), .C(n12538), .D(n17813), .Z(n12569)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2664_4_lut.init = 16'hafac;
    LUT4 i5074_2_lut (.A(d4_adj_5713[0]), .B(d3_adj_5712[0]), .Z(d4_71__N_634_adj_5729[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5074_2_lut.init = 16'h6666;
    LUT4 i5073_2_lut (.A(d5_adj_5714[0]), .B(d4_adj_5713[0]), .Z(d5_71__N_706_adj_5730[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5073_2_lut.init = 16'h6666;
    LUT4 i2700_4_lut (.A(n170), .B(n2594), .C(n12538), .D(n17813), .Z(n12605)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2700_4_lut.init = 16'hafac;
    LUT4 i2660_4_lut (.A(n263), .B(n11977), .C(n12538), .D(n17813), 
         .Z(n12565)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2660_4_lut.init = 16'hafac;
    LUT4 i2083_3_lut (.A(n11976), .B(n259), .C(led_c_4), .Z(n11977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2083_3_lut.init = 16'hcaca;
    LUT4 i3171_4_lut_4_lut (.A(led_c_4), .B(n17817), .C(n235), .D(n229_adj_5057), 
         .Z(n2617)) /* synthesis lut_function=(A (C)+!A !(B+!(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3171_4_lut_4_lut.init = 16'hb1a0;
    LUT4 i3184_4_lut_4_lut (.A(n18053), .B(n17817), .C(n166), .D(n160_adj_5034), 
         .Z(n2594)) /* synthesis lut_function=(A (C)+!A !(B+!(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3184_4_lut_4_lut.init = 16'hb1a0;
    LUT4 i5063_2_lut (.A(d2[0]), .B(d1[0]), .Z(d2_71__N_490[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5063_2_lut.init = 16'h6666;
    LUT4 i2658_3_lut (.A(n269), .B(n2695), .C(n12538), .Z(n12563)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2658_3_lut.init = 16'hacac;
    LUT4 i3189_4_lut_4_lut (.A(led_c_4), .B(n17817), .C(n139), .D(n133_adj_5025), 
         .Z(n2585)) /* synthesis lut_function=(A (C)+!A (B+(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3189_4_lut_4_lut.init = 16'hf5e4;
    LUT4 i2080_3_lut_4_lut (.A(n17823), .B(n16869), .C(led_c_0), .D(n268_adj_5070), 
         .Z(n11974)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i2080_3_lut_4_lut.init = 16'hf780;
    LUT4 i5046_2_lut (.A(d1[0]), .B(MixerOutSin[0]), .Z(d1_71__N_418[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5046_2_lut.init = 16'h6666;
    LUT4 i3188_4_lut_4_lut (.A(n18053), .B(n17817), .C(n142), .D(n136_adj_5026), 
         .Z(n2586)) /* synthesis lut_function=(A (C)+!A (B+(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3188_4_lut_4_lut.init = 16'hf5e4;
    LUT4 i2698_3_lut (.A(n173), .B(n2663), .C(n12538), .Z(n12603)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2698_3_lut.init = 16'hacac;
    LUT4 i3166_4_lut_4_lut (.A(led_c_4), .B(n17817), .C(n271), .D(n265_adj_5069), 
         .Z(n2629)) /* synthesis lut_function=(A (C)+!A !(B+!(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3166_4_lut_4_lut.init = 16'hb1a0;
    LUT4 mux_339_i51_4_lut (.A(n3901), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2663)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i51_4_lut.init = 16'h303a;
    LUT4 mux_843_i50_3_lut (.A(n163_adj_5035), .B(n169), .C(n18053), .Z(n3901)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i50_3_lut.init = 16'hcaca;
    LUT4 i2696_4_lut (.A(n176), .B(n12003), .C(n12538), .D(n17813), 
         .Z(n12601)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2696_4_lut.init = 16'hafac;
    LUT4 i2109_3_lut (.A(n12002), .B(n172), .C(n18053), .Z(n12003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2109_3_lut.init = 16'hcaca;
    LUT4 i2692_4_lut (.A(n185), .B(n11999), .C(n12538), .D(n17813), 
         .Z(n12597)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2692_4_lut.init = 16'hafac;
    LUT4 mux_339_i19_4_lut (.A(n3933), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2695)) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i19_4_lut.init = 16'h3f3a;
    LUT4 mux_843_i18_3_lut (.A(n259_adj_5067), .B(n265), .C(led_c_4), 
         .Z(n3933)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i18_3_lut.init = 16'hcaca;
    LUT4 i2105_3_lut (.A(n11998), .B(n181), .C(n18053), .Z(n11999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2105_3_lut.init = 16'hcaca;
    LUT4 i2102_3_lut_4_lut (.A(n17823), .B(n16869), .C(led_c_0), .D(n181_adj_5041), 
         .Z(n11996)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i2102_3_lut_4_lut.init = 16'hf780;
    LUT4 i2344_3_lut (.A(n12246), .B(n299), .C(n12538), .Z(n12247)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2344_3_lut.init = 16'hcaca;
    LUT4 i2656_3_lut (.A(n272), .B(n2696), .C(n12538), .Z(n12561)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2656_3_lut.init = 16'hacac;
    LUT4 mux_339_i18_4_lut (.A(n3934), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2696)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i18_4_lut.init = 16'h303a;
    LUT4 i2346_3_lut (.A(n12248), .B(n281), .C(n12538), .Z(n12249)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2346_3_lut.init = 16'hcaca;
    LUT4 mux_843_i17_3_lut (.A(n262_adj_5068), .B(n268), .C(n18053), .Z(n3934)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i17_3_lut.init = 16'hcaca;
    LUT4 i2348_3_lut (.A(n12250), .B(n257), .C(n12538), .Z(n12251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2348_3_lut.init = 16'hcaca;
    LUT4 i2350_3_lut (.A(n12252), .B(n248), .C(n12538), .Z(n12253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2350_3_lut.init = 16'hcaca;
    LUT4 i5043_2_lut (.A(d1_adj_5710[0]), .B(MixerOutCos[0]), .Z(d1_71__N_418_adj_5726[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5043_2_lut.init = 16'h6666;
    LUT4 i5047_2_lut (.A(phase_inc_carrGen1[0]), .B(phase_accum_adj_5702[0]), 
         .Z(n321)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5047_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_adj_79 (.A(led_c_2), .B(led_c_1), .Z(n16869)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_79.init = 16'h8888;
    LUT4 i2352_3_lut (.A(n12254), .B(n242), .C(n12538), .Z(n12255)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2352_3_lut.init = 16'hcaca;
    LUT4 i3182_4_lut_4_lut (.A(n18053), .B(n17817), .C(n178), .D(n172_adj_5038), 
         .Z(n2598)) /* synthesis lut_function=(A (C)+!A (B+(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3182_4_lut_4_lut.init = 16'hf5e4;
    LUT4 i3180_4_lut_4_lut (.A(n18053), .B(n17817), .C(n190), .D(n184_adj_5042), 
         .Z(n2602)) /* synthesis lut_function=(A (C)+!A (B+(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3180_4_lut_4_lut.init = 16'hf5e4;
    LUT4 i5062_2_lut (.A(d3[0]), .B(d2[0]), .Z(d3_71__N_562[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5062_2_lut.init = 16'h6666;
    LUT4 mux_339_i14_4_lut (.A(n3938), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2700)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i14_4_lut.init = 16'h303a;
    CCU2C _add_1_1374_add_4_2 (.A0(d1_adj_5710[0]), .B0(MixerOutCos[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5710[1]), .B1(MixerOutCos[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14993), .S1(d1_71__N_418_adj_5726[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1374_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1374_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1374_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1374_add_4_2.INJECT1_1 = "NO";
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 mux_843_i13_3_lut (.A(n274_adj_5072), .B(n280), .C(n18053), .Z(n3938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i13_3_lut.init = 16'hcaca;
    LUT4 i2349_3_lut (.A(led_c_1), .B(n244), .C(n18053), .Z(n12252)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2349_3_lut.init = 16'hc5c5;
    LUT4 i2650_3_lut (.A(n284), .B(n2700), .C(n12538), .Z(n12555)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2650_3_lut.init = 16'hacac;
    CCU2C add_3659_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1874[17]), .C0(n38), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1874[17]), 
          .C1(n35_adj_4742), .D1(VCC_net), .CIN(n16373), .COUT(n16374), 
          .S0(n45), .S1(n42));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3659_9.INIT0 = 16'h6969;
    defparam add_3659_9.INIT1 = 16'h6969;
    defparam add_3659_9.INJECT1_0 = "NO";
    defparam add_3659_9.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_26 (.A0(d_d6[59]), .B0(d6[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[60]), .B1(d6[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16240), .COUT(n16241), .S0(n114_adj_5477), .S1(n111_adj_5476));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_24 (.A0(d_d6[57]), .B0(d6[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[58]), .B1(d6[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16239), .COUT(n16240), .S0(n120_adj_5479), .S1(n117_adj_5478));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_22 (.A0(d_d6[55]), .B0(d6[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[56]), .B1(d6[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16238), .COUT(n16239), .S0(n126_adj_5481), .S1(n123_adj_5480));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_20 (.A0(d_d6[53]), .B0(d6[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[54]), .B1(d6[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16237), .COUT(n16238), .S0(n132_adj_5483), .S1(n129_adj_5482));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_20.INJECT1_1 = "NO";
    LUT4 i2347_3_lut (.A(led_c_1), .B(n253), .C(led_c_4), .Z(n12250)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2347_3_lut.init = 16'hc5c5;
    CCU2C _add_1_1559_add_4_18 (.A0(d_d6[51]), .B0(d6[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[52]), .B1(d6[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16236), .COUT(n16237), .S0(n138_adj_5485), .S1(n135_adj_5484));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_16 (.A0(d_d6[49]), .B0(d6[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[50]), .B1(d6[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16235), .COUT(n16236), .S0(n144_adj_5487), .S1(n141_adj_5486));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_16.INJECT1_1 = "NO";
    FD1S3AX o_Rx_Byte_i1 (.D(o_Rx_Byte1[0]), .CK(clk_80mhz), .Q(led_c_0));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    CCU2C _add_1_1559_add_4_14 (.A0(d_d6[47]), .B0(d6[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[48]), .B1(d6[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16234), .COUT(n16235), .S0(n150_adj_5489), .S1(n147_adj_5488));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_14.INJECT1_1 = "NO";
    LUT4 mux_305_i1_4_lut (.A(n323), .B(led_c_0), .C(n17815), .D(n17809), 
         .Z(n1994)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_305_i1_4_lut.init = 16'h0a3a;
    LUT4 i3223_2_lut_rep_210 (.A(n18053), .B(led_c_5), .Z(n17832)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3223_2_lut_rep_210.init = 16'h8888;
    CCU2C _add_1_1559_add_4_12 (.A0(d_d6[45]), .B0(d6[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[46]), .B1(d6[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16233), .COUT(n16234), .S0(n156_adj_5491), .S1(n153_adj_5490));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_12.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_212 (.A(led_c_2), .B(led_c_1), .C(led_c_0), .Z(n17834)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i1_3_lut_rep_212.init = 16'h1414;
    LUT4 i2341_3_lut_4_lut_4_lut (.A(led_c_2), .B(led_c_1), .C(led_c_0), 
         .D(n17823), .Z(n12701)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B !((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i2341_3_lut_4_lut_4_lut.init = 16'he4f0;
    CCU2C _add_1_1559_add_4_10 (.A0(d_d6[43]), .B0(d6[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[44]), .B1(d6[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16232), .COUT(n16233), .S0(n162_adj_5493), .S1(n159_adj_5492));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_10.INJECT1_1 = "NO";
    LUT4 i2072_3_lut_4_lut_4_lut (.A(led_c_0), .B(n289_adj_5077), .C(n16869), 
         .D(n17823), .Z(n11966)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;
    defparam i2072_3_lut_4_lut_4_lut.init = 16'h5ccc;
    LUT4 i3170_4_lut_4_lut (.A(led_c_4), .B(n17817), .C(n247), .D(n241_adj_5061), 
         .Z(n2621)) /* synthesis lut_function=(A (C)+!A (B+(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3170_4_lut_4_lut.init = 16'hf5e4;
    LUT4 i2106_3_lut_4_lut_4_lut (.A(led_c_0), .B(n169_adj_5037), .C(n16869), 
         .D(n17823), .Z(n12000)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;
    defparam i2106_3_lut_4_lut_4_lut.init = 16'h5ccc;
    LUT4 i2094_3_lut_4_lut_4_lut (.A(led_c_0), .B(n211_adj_5051), .C(n16869), 
         .D(n17823), .Z(n11988)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;
    defparam i2094_3_lut_4_lut_4_lut.init = 16'h5ccc;
    CCU2C _add_1_1559_add_4_8 (.A0(d_d6[41]), .B0(d6[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[42]), .B1(d6[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16231), .COUT(n16232), .S0(n168_adj_5495), .S1(n165_adj_5494));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_6 (.A0(d_d6[39]), .B0(d6[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[40]), .B1(d6[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16230), .COUT(n16231), .S0(n174_adj_5497), .S1(n171_adj_5496));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1559_add_4_4 (.A0(d_d6[37]), .B0(d6[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[38]), .B1(d6[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16229), .COUT(n16230), .S0(n180_adj_5499), .S1(n177_adj_5498));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1559_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_4.INJECT1_1 = "NO";
    LUT4 i2112_3_lut_4_lut_4_lut (.A(led_c_0), .B(n148_adj_5030), .C(n16869), 
         .D(n17823), .Z(n12006)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;
    defparam i2112_3_lut_4_lut_4_lut.init = 16'h5ccc;
    LUT4 i2108_3_lut_4_lut_4_lut (.A(led_c_0), .B(n166_adj_5036), .C(n16869), 
         .D(n17823), .Z(n12002)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;
    defparam i2108_3_lut_4_lut_4_lut.init = 16'h5ccc;
    PLL PLL_inst (.clk_25mhz_c(clk_25mhz_c), .clk_80mhz(clk_80mhz), .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(97[8] 100[5])
    LUT4 i2088_3_lut_4_lut_4_lut (.A(led_c_0), .B(n235_adj_5059), .C(n16869), 
         .D(n17823), .Z(n11982)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;
    defparam i2088_3_lut_4_lut_4_lut.init = 16'h5ccc;
    LUT4 i2092_3_lut_4_lut_4_lut (.A(led_c_0), .B(n223_adj_5055), .C(n16869), 
         .D(n17823), .Z(n11986)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;
    defparam i2092_3_lut_4_lut_4_lut.init = 16'h5ccc;
    LUT4 i1_4_lut_adj_80 (.A(n16944), .B(n17827), .C(n18053), .D(n39_adj_4738), 
         .Z(n16837)) /* synthesis lut_function=(A (B)+!A !((C+!(D))+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i1_4_lut_adj_80.init = 16'h8c88;
    CCU2C _add_1_1559_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[36]), .B1(d6[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16229), .S1(n183_adj_5500));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1559_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1559_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1559_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1559_add_4_2.INJECT1_1 = "NO";
    LUT4 i2078_3_lut_4_lut_4_lut (.A(led_c_0), .B(n271_adj_5071), .C(n16869), 
         .D(n17823), .Z(n11972)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;
    defparam i2078_3_lut_4_lut_4_lut.init = 16'h5ccc;
    LUT4 i2068_3_lut_4_lut_4_lut (.A(led_c_0), .B(n298_adj_5080), .C(n16869), 
         .D(n17823), .Z(n11962)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;
    defparam i2068_3_lut_4_lut_4_lut.init = 16'h5ccc;
    LUT4 i1_4_lut_adj_81 (.A(led_c_2), .B(n17523), .C(led_c_4), .D(led_c_0), 
         .Z(n16944)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(200[9] 212[17])
    defparam i1_4_lut_adj_81.init = 16'h1110;
    LUT4 i2100_3_lut_4_lut_4_lut (.A(led_c_0), .B(n187_adj_5043), .C(n16869), 
         .D(n17823), .Z(n11994)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;
    defparam i2100_3_lut_4_lut_4_lut.init = 16'h5ccc;
    LUT4 i2686_4_lut (.A(n206), .B(n2606), .C(n12538), .D(n17813), .Z(n12591)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2686_4_lut.init = 16'hafac;
    CCU2C _add_1_1475_add_4_38 (.A0(d_d7_adj_5718[35]), .B0(d7_adj_5717[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16228), .S0(d8_71__N_1603_adj_5744[35]), 
          .S1(cout_adj_5501));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1475_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_38.INJECT1_1 = "NO";
    LUT4 i3103_rep_99_2_lut (.A(led_c_1), .B(led_c_3), .Z(n17523)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3103_rep_99_2_lut.init = 16'heeee;
    LUT4 i2086_3_lut_4_lut_4_lut (.A(led_c_0), .B(n238_adj_5060), .C(n16869), 
         .D(n17823), .Z(n11980)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;
    defparam i2086_3_lut_4_lut_4_lut.init = 16'h5ccc;
    CCU2C _add_1_1475_add_4_36 (.A0(d_d7_adj_5718[33]), .B0(d7_adj_5717[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[34]), .B1(d7_adj_5717[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16227), .COUT(n16228), .S0(d8_71__N_1603_adj_5744[33]), 
          .S1(d8_71__N_1603_adj_5744[34]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_36.INJECT1_1 = "NO";
    LUT4 i2684_4_lut (.A(n209), .B(n2607), .C(n12538), .D(n17813), .Z(n12589)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2684_4_lut.init = 16'hafac;
    LUT4 i2682_4_lut (.A(n212), .B(n11991), .C(n12538), .D(n17813), 
         .Z(n12587)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2682_4_lut.init = 16'hafac;
    LUT4 i5949_3_lut_4_lut_4_lut (.A(led_c_0), .B(n16829), .C(led_c_5), 
         .D(led_c_4), .Z(n17032)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i5949_3_lut_4_lut_4_lut.init = 16'h2000;
    LUT4 i2097_3_lut (.A(n11990), .B(n208), .C(n18053), .Z(n11991)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2097_3_lut.init = 16'hcaca;
    LUT4 i2076_3_lut_4_lut_4_lut (.A(led_c_0), .B(n277_adj_5073), .C(n16869), 
         .D(n17823), .Z(n11970)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;
    defparam i2076_3_lut_4_lut_4_lut.init = 16'h5ccc;
    LUT4 i2680_4_lut (.A(n215), .B(n2609), .C(n12538), .D(n17813), .Z(n12585)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2680_4_lut.init = 16'hafac;
    LUT4 i1_2_lut_rep_213 (.A(led_c_6), .B(led_c_7), .Z(n17835)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_213.init = 16'h2222;
    FD1S3AX o_Rx_DV_40_rep_258 (.D(o_Rx_DV1), .CK(clk_80mhz), .Q(clk_80mhz_enable_1411));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam o_Rx_DV_40_rep_258.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_205_3_lut (.A(led_c_6), .B(led_c_7), .C(led_c_5), 
         .Z(n17827)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_rep_205_3_lut.init = 16'h2020;
    LUT4 i3174_4_lut_4_lut (.A(led_c_4), .B(n17817), .C(n223), .D(n217_adj_5053), 
         .Z(n2613)) /* synthesis lut_function=(A (C)+!A (B+(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam i3174_4_lut_4_lut.init = 16'hf5e4;
    LUT4 i2520_4_lut_then_4_lut (.A(led_c_2), .B(led_c_4), .C(led_c_3), 
         .D(led_c_1), .Z(n17837)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(44[22:25])
    defparam i2520_4_lut_then_4_lut.init = 16'h2000;
    LUT4 i2520_4_lut_else_4_lut (.A(led_c_2), .B(led_c_4), .C(led_c_3), 
         .D(led_c_1), .Z(n17836)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(44[22:25])
    defparam i2520_4_lut_else_4_lut.init = 16'h0004;
    LUT4 i2678_3_lut (.A(n218), .B(n2678), .C(n12538), .Z(n12583)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2678_3_lut.init = 16'hacac;
    FD1S3AX o_Rx_DV_40_rep_257 (.D(o_Rx_DV1), .CK(clk_80mhz), .Q(n18096));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam o_Rx_DV_40_rep_257.GSR = "ENABLED";
    LUT4 mux_339_i36_4_lut (.A(n3916), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2678)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i36_4_lut.init = 16'hc0ca;
    LUT4 i1_2_lut_rep_203_3_lut_4_lut (.A(led_c_6), .B(led_c_7), .C(n18096), 
         .D(led_c_5), .Z(n17825)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_rep_203_3_lut_4_lut.init = 16'h2000;
    LUT4 mux_843_i35_3_lut (.A(n208_adj_5050), .B(n214), .C(n18053), .Z(n3916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i35_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut (.A(led_c_6), .B(led_c_7), .C(n18096), .Z(n17075)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i2676_3_lut (.A(n224), .B(n2680), .C(n12538), .Z(n12581)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2676_3_lut.init = 16'hacac;
    LUT4 mux_339_i34_4_lut (.A(n3918), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2680)) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i34_4_lut.init = 16'h3f3a;
    VLO i1 (.Z(GND_net));
    LUT4 i2710_3_lut (.A(n149), .B(n2655), .C(n12538), .Z(n12615)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2710_3_lut.init = 16'hacac;
    LUT4 mux_339_i59_4_lut (.A(n3893), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2655)) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i59_4_lut.init = 16'h3f3a;
    LUT4 mux_843_i58_3_lut (.A(n139_adj_5027), .B(n145), .C(led_c_4), 
         .Z(n3893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i58_3_lut.init = 16'hcaca;
    LUT4 i2708_3_lut (.A(n155), .B(n2657), .C(n12538), .Z(n12613)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2708_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_4_lut (.A(n17823), .B(n16869), .C(n17834), .D(n18053), 
         .Z(n17081)) /* synthesis lut_function=(A (B+(C+(D)))+!A (D)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i1_2_lut_4_lut.init = 16'hffa8;
    LUT4 mux_339_i57_4_lut (.A(n3895), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i57_4_lut.init = 16'hcfca;
    LUT4 mux_843_i33_3_lut (.A(n214_adj_5052), .B(n220), .C(n18053), .Z(n3918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i33_3_lut.init = 16'hcaca;
    CCU2C _add_1_1475_add_4_34 (.A0(d_d7_adj_5718[31]), .B0(d7_adj_5717[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[32]), .B1(d7_adj_5717[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16226), .COUT(n16227), .S0(d8_71__N_1603_adj_5744[31]), 
          .S1(d8_71__N_1603_adj_5744[32]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_34.INJECT1_1 = "NO";
    FD1P3IX CICGain__i2 (.D(n16842), .SP(clk_80mhz_enable_1411), .CD(n12710), 
            .CK(clk_80mhz), .Q(CICGain[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam CICGain__i2.GSR = "ENABLED";
    CCU2C _add_1_1475_add_4_32 (.A0(d_d7_adj_5718[29]), .B0(d7_adj_5717[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[30]), .B1(d7_adj_5717[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16225), .COUT(n16226), .S0(d8_71__N_1603_adj_5744[29]), 
          .S1(d8_71__N_1603_adj_5744[30]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_32.INJECT1_1 = "NO";
    FD1S3AX o_Rx_Byte_i5_rep_214 (.D(o_Rx_Byte1[4]), .CK(clk_80mhz), .Q(n18053));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam o_Rx_Byte_i5_rep_214.GSR = "ENABLED";
    CCU2C _add_1_1475_add_4_30 (.A0(d_d7_adj_5718[27]), .B0(d7_adj_5717[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[28]), .B1(d7_adj_5717[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16224), .COUT(n16225), .S0(d8_71__N_1603_adj_5744[27]), 
          .S1(d8_71__N_1603_adj_5744[28]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_28 (.A0(d_d7_adj_5718[25]), .B0(d7_adj_5717[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[26]), .B1(d7_adj_5717[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16223), .COUT(n16224), .S0(d8_71__N_1603_adj_5744[25]), 
          .S1(d8_71__N_1603_adj_5744[26]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_28.INJECT1_1 = "NO";
    LUT4 mux_843_i56_3_lut (.A(n145_adj_5029), .B(n151), .C(led_c_4), 
         .Z(n3895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i56_3_lut.init = 16'hcaca;
    CCU2C _add_1_1475_add_4_26 (.A0(d_d7_adj_5718[23]), .B0(d7_adj_5717[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[24]), .B1(d7_adj_5717[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16222), .COUT(n16223), .S0(d8_71__N_1603_adj_5744[23]), 
          .S1(d8_71__N_1603_adj_5744[24]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_24 (.A0(d_d7_adj_5718[21]), .B0(d7_adj_5717[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[22]), .B1(d7_adj_5717[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16221), .COUT(n16222), .S0(d8_71__N_1603_adj_5744[21]), 
          .S1(d8_71__N_1603_adj_5744[22]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_22 (.A0(d_d7_adj_5718[19]), .B0(d7_adj_5717[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[20]), .B1(d7_adj_5717[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16220), .COUT(n16221), .S0(d8_71__N_1603_adj_5744[19]), 
          .S1(d8_71__N_1603_adj_5744[20]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_20 (.A0(d_d7_adj_5718[17]), .B0(d7_adj_5717[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[18]), .B1(d7_adj_5717[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16219), .COUT(n16220), .S0(d8_71__N_1603_adj_5744[17]), 
          .S1(d8_71__N_1603_adj_5744[18]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_18 (.A0(d_d7_adj_5718[15]), .B0(d7_adj_5717[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[16]), .B1(d7_adj_5717[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16218), .COUT(n16219), .S0(d8_71__N_1603_adj_5744[15]), 
          .S1(d8_71__N_1603_adj_5744[16]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_16 (.A0(d_d7_adj_5718[13]), .B0(d7_adj_5717[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[14]), .B1(d7_adj_5717[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16217), .COUT(n16218), .S0(d8_71__N_1603_adj_5744[13]), 
          .S1(d8_71__N_1603_adj_5744[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_14 (.A0(d_d7_adj_5718[11]), .B0(d7_adj_5717[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[12]), .B1(d7_adj_5717[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16216), .COUT(n16217), .S0(d8_71__N_1603_adj_5744[11]), 
          .S1(d8_71__N_1603_adj_5744[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_12 (.A0(d_d7_adj_5718[9]), .B0(d7_adj_5717[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[10]), .B1(d7_adj_5717[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16215), .COUT(n16216), .S0(d8_71__N_1603_adj_5744[9]), 
          .S1(d8_71__N_1603_adj_5744[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_12.INJECT1_1 = "NO";
    LUT4 i2674_3_lut (.A(n230), .B(n2682), .C(n12538), .Z(n12579)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2674_3_lut.init = 16'hacac;
    CCU2C _add_1_1475_add_4_10 (.A0(d_d7_adj_5718[7]), .B0(d7_adj_5717[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[8]), .B1(d7_adj_5717[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16214), .COUT(n16215), .S0(d8_71__N_1603_adj_5744[7]), 
          .S1(d8_71__N_1603_adj_5744[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_8 (.A0(d_d7_adj_5718[5]), .B0(d7_adj_5717[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[6]), .B1(d7_adj_5717[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16213), .COUT(n16214), .S0(d8_71__N_1603_adj_5744[5]), 
          .S1(d8_71__N_1603_adj_5744[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_8.INJECT1_1 = "NO";
    LUT4 i2648_4_lut (.A(n287), .B(n11971), .C(n12538), .D(n17813), 
         .Z(n12553)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2648_4_lut.init = 16'hafac;
    CCU2C _add_1_1454_add_4_7 (.A0(d4[40]), .B0(cout_adj_2810), .C0(n171_adj_5316), 
          .D0(d5[40]), .A1(d4[41]), .B1(cout_adj_2810), .C1(n168_adj_5315), 
          .D1(d5[41]), .CIN(n16046), .COUT(n16047), .S0(d5_71__N_706[40]), 
          .S1(d5_71__N_706[41]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_6 (.A0(d_d7_adj_5718[3]), .B0(d7_adj_5717[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[4]), .B1(d7_adj_5717[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16212), .COUT(n16213), .S0(d8_71__N_1603_adj_5744[3]), 
          .S1(d8_71__N_1603_adj_5744[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_4 (.A0(d_d7_adj_5718[1]), .B0(d7_adj_5717[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5718[2]), .B1(d7_adj_5717[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16211), .COUT(n16212), .S0(d8_71__N_1603_adj_5744[1]), 
          .S1(d8_71__N_1603_adj_5744[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1475_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_35 (.A0(d6_adj_5715[68]), .B0(cout_adj_5464), 
          .C0(n87_adj_4881), .D0(n5_adj_4759), .A1(d6_adj_5715[69]), .B1(cout_adj_5464), 
          .C1(n84_adj_4880), .D1(n4_adj_4760), .CIN(n16190), .COUT(n16191), 
          .S0(d7_71__N_1531_adj_5743[68]), .S1(d7_71__N_1531_adj_5743[69]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_4 (.A0(d_d_tmp[37]), .B0(d_tmp[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[38]), .B1(d_tmp[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16193), .COUT(n16194), .S0(n180_adj_5536), 
          .S1(n177_adj_5535));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1475_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7_adj_5718[0]), .B1(d7_adj_5717[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16211), .S1(d8_71__N_1603_adj_5744[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1475_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1475_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1475_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1475_add_4_2.INJECT1_1 = "NO";
    PFUMX i2702 (.BLUT(n12004), .ALUT(n12261), .C0(n17389), .Z(n12607));
    CCU2C _add_1_1556_add_4_38 (.A0(d_d_tmp[71]), .B0(d_tmp[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16210), .S0(n78_adj_5502));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1556_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_38.INJECT1_1 = "NO";
    LUT4 mux_305_i64_4_lut_4_lut (.A(n17822), .B(n12538), .C(n8_adj_4728), 
         .D(n134), .Z(n1931)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam mux_305_i64_4_lut_4_lut.init = 16'h5410;
    CCU2C _add_1_1556_add_4_36 (.A0(d_d_tmp[69]), .B0(d_tmp[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[70]), .B1(d_tmp[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16209), .COUT(n16210), .S0(n84_adj_5504), 
          .S1(n81_adj_5503));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_34 (.A0(d_d_tmp[67]), .B0(d_tmp[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[68]), .B1(d_tmp[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16208), .COUT(n16209), .S0(n90_adj_5506), 
          .S1(n87_adj_5505));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_32 (.A0(d_d_tmp[65]), .B0(d_tmp[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[66]), .B1(d_tmp[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16207), .COUT(n16208), .S0(n96_adj_5508), 
          .S1(n93_adj_5507));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_32.INJECT1_1 = "NO";
    LUT4 mux_305_i63_4_lut_4_lut (.A(n17822), .B(n12538), .C(n8_adj_4727), 
         .D(n137), .Z(n1932)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam mux_305_i63_4_lut_4_lut.init = 16'h5410;
    CCU2C _add_1_1556_add_4_30 (.A0(d_d_tmp[63]), .B0(d_tmp[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[64]), .B1(d_tmp[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16206), .COUT(n16207), .S0(n102_adj_5510), 
          .S1(n99_adj_5509));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_30.INJECT1_1 = "NO";
    PFUMX i2694 (.BLUT(n12000), .ALUT(n12259), .C0(n17389), .Z(n12599));
    CCU2C _add_1_1556_add_4_28 (.A0(d_d_tmp[61]), .B0(d_tmp[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[62]), .B1(d_tmp[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16205), .COUT(n16206), .S0(n108_adj_5512), 
          .S1(n105_adj_5511));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_33 (.A0(d6_adj_5715[66]), .B0(cout_adj_5464), 
          .C0(n93_adj_4883), .D0(n7_adj_4757), .A1(d6_adj_5715[67]), .B1(cout_adj_5464), 
          .C1(n90_adj_4882), .D1(n6_adj_4758), .CIN(n16189), .COUT(n16190), 
          .S0(d7_71__N_1531_adj_5743[66]), .S1(d7_71__N_1531_adj_5743[67]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[36]), .B1(d_tmp[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16193), .S1(n183_adj_5537));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1556_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_26 (.A0(d_d_tmp[59]), .B0(d_tmp[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[60]), .B1(d_tmp[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16204), .COUT(n16205), .S0(n114_adj_5514), 
          .S1(n111_adj_5513));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_24 (.A0(d_d_tmp[57]), .B0(d_tmp[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[58]), .B1(d_tmp[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16203), .COUT(n16204), .S0(n120_adj_5516), 
          .S1(n117_adj_5515));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_24.INJECT1_1 = "NO";
    LUT4 mux_305_i62_4_lut_4_lut (.A(n17822), .B(n12538), .C(n8_adj_4730), 
         .D(n140), .Z(n1933)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam mux_305_i62_4_lut_4_lut.init = 16'h5410;
    CCU2C _add_1_1556_add_4_22 (.A0(d_d_tmp[55]), .B0(d_tmp[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[56]), .B1(d_tmp[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16202), .COUT(n16203), .S0(n126_adj_5518), 
          .S1(n123_adj_5517));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1544_add_4_36 (.A0(d2_adj_5711[69]), .B0(d1_adj_5710[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5711[70]), .B1(d1_adj_5710[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16039), .COUT(n16040), .S0(n84_adj_5610), 
          .S1(n81_adj_5609));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1544_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1544_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1544_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1544_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1454_add_4_25 (.A0(d4[58]), .B0(cout_adj_2810), .C0(n117_adj_5298), 
          .D0(d5[58]), .A1(d4[59]), .B1(cout_adj_2810), .C1(n114_adj_5297), 
          .D1(d5[59]), .CIN(n16055), .COUT(n16056), .S0(d5_71__N_706[58]), 
          .S1(d5_71__N_706[59]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_25.INJECT1_1 = "NO";
    CCU2C add_3659_7 (.A0(d_out_d_11__N_1874[17]), .B0(n44), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1874[17]), 
          .C1(n41), .D1(VCC_net), .CIN(n16372), .COUT(n16373), .S0(n51), 
          .S1(n48));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3659_7.INIT0 = 16'h9995;
    defparam add_3659_7.INIT1 = 16'h6969;
    defparam add_3659_7.INJECT1_0 = "NO";
    defparam add_3659_7.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_20 (.A0(d_d_tmp[53]), .B0(d_tmp[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[54]), .B1(d_tmp[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16201), .COUT(n16202), .S0(n132_adj_5520), 
          .S1(n129_adj_5519));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_18 (.A0(d_d_tmp[51]), .B0(d_tmp[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[52]), .B1(d_tmp[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16200), .COUT(n16201), .S0(n138_adj_5522), 
          .S1(n135_adj_5521));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_16 (.A0(d_d_tmp[49]), .B0(d_tmp[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[50]), .B1(d_tmp[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16199), .COUT(n16200), .S0(n144_adj_5524), 
          .S1(n141_adj_5523));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_14 (.A0(d_d_tmp[47]), .B0(d_tmp[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[48]), .B1(d_tmp[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16198), .COUT(n16199), .S0(n150_adj_5526), 
          .S1(n147_adj_5525));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_12 (.A0(d_d_tmp[45]), .B0(d_tmp[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[46]), .B1(d_tmp[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16197), .COUT(n16198), .S0(n156_adj_5528), 
          .S1(n153_adj_5527));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_10 (.A0(d_d_tmp[43]), .B0(d_tmp[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[44]), .B1(d_tmp[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16196), .COUT(n16197), .S0(n162_adj_5530), 
          .S1(n159_adj_5529));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_10.INJECT1_1 = "NO";
    PFUMX i2688 (.BLUT(n11992), .ALUT(n12257), .C0(n17389), .Z(n12593));
    CCU2C _add_1_1418_add_4_37 (.A0(d6_adj_5715[70]), .B0(cout_adj_5464), 
          .C0(n81_adj_4879), .D0(n3_adj_4761), .A1(d6_adj_5715[71]), .B1(cout_adj_5464), 
          .C1(n78_adj_4878), .D1(n2_adj_4762), .CIN(n16191), .S0(d7_71__N_1531_adj_5743[70]), 
          .S1(d7_71__N_1531_adj_5743[71]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1418_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1418_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1418_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1556_add_4_8 (.A0(d_d_tmp[41]), .B0(d_tmp[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[42]), .B1(d_tmp[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16195), .COUT(n16196), .S0(n168_adj_5532), 
          .S1(n165_adj_5531));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1556_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1556_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1556_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1556_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1553_add_4_14 (.A0(d5_adj_5714[47]), .B0(d4_adj_5713[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5714[48]), .B1(d4_adj_5713[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16158), .COUT(n16159), .S0(n150_adj_5562), 
          .S1(n147_adj_5561));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1553_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1553_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1553_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1553_add_4_14.INJECT1_1 = "NO";
    FD1P3IX phase_inc_carrGen_i0_i45 (.D(n12595), .SP(clk_80mhz_enable_1411), 
            .CD(n17822), .CK(clk_80mhz), .Q(phase_inc_carrGen[45]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(186[11] 214[6])
    defparam phase_inc_carrGen_i0_i45.GSR = "ENABLED";
    nco_sig nco_sig_inst (.\phase_accum[63] (phase_accum[63]), .sinGen_c(sinGen_c)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(114[4] 120[5])
    \CIC(WIDTH=72,DECIMATION_RATIO=4096)  CIC_cos_inst (.d_tmp({d_tmp_adj_5708}), 
            .clk_80mhz(clk_80mhz), .d5({d5_adj_5714}), .d_d_tmp({d_d_tmp_adj_5709}), 
            .d2({d2_adj_5711}), .d2_71__N_490({d2_71__N_490_adj_5727}), 
            .d3({d3_adj_5712}), .d3_71__N_562({d3_71__N_562_adj_5728}), 
            .d4({d4_adj_5713}), .d4_71__N_634({d4_71__N_634_adj_5729}), 
            .d5_71__N_706({d5_71__N_706_adj_5730}), .d6({d6_adj_5715}), 
            .d6_71__N_1459({d6_71__N_1459_adj_5742}), .d_d6({d_d6_adj_5716}), 
            .d7({d7_adj_5717}), .d7_71__N_1531({d7_71__N_1531_adj_5743}), 
            .d_d7({d_d7_adj_5718}), .d8({d8_adj_5719}), .d8_71__N_1603({d8_71__N_1603_adj_5744}), 
            .d_d8({d_d8_adj_5720}), .d9({d9_adj_5721}), .d9_71__N_1675({d9_71__N_1675_adj_5745}), 
            .d_d9({d_d9_adj_5722}), .CIC1_outCos({CIC1_outCos}), .d1({d1_adj_5710}), 
            .d1_71__N_418({d1_71__N_418_adj_5726}), .count({count_adj_5725}), 
            .n87_adj_228({n36_adj_5208, n39_adj_5209, n42_adj_5210, n45_adj_5211, 
            n48_adj_5212, n51_adj_5213, n54_adj_5214, n57_adj_5215, 
            n60_adj_5216, n63_adj_5217, n66_adj_5218, n69_adj_5219, 
            n72_adj_5220, n75_adj_5221, n78_adj_5222, n81_adj_5223}), 
            .n23(n23_adj_4557), .n10(n10_adj_4771), .n35(n35_adj_4796), 
            .n10_adj_115(n10_adj_4754), .n22(n22_adj_4576), .n13(n13_adj_4744), 
            .n12(n12_adj_4751), .n15(n15_adj_2794), .n34(n34_adj_4795), 
            .n37(n37_adj_4798), .n14(n14_adj_4732), .n17(n17_adj_4595), 
            .n36_adj_116(n36_adj_4797), .n16(n16_adj_4731), .n3(n3_adj_4800), 
            .n2(n2_adj_4799), .n5(n5_adj_4802), .n4(n4_adj_4801), .n7(n7_adj_4804), 
            .n6(n6_adj_4803), .n9(n9_adj_4806), .n8(n8_adj_4805), .\CICGain[1] (CICGain[1]), 
            .\d10[60] (d10_adj_5723[60]), .\d10[59] (d10_adj_5723[59]), 
            .\d10[61] (d10_adj_5723[61]), .\d10[62] (d10_adj_5723[62]), 
            .\d10[63] (d10_adj_5723[63]), .\d10[64] (d10_adj_5723[64]), 
            .\d10[65] (d10_adj_5723[65]), .\d10[66] (d10_adj_5723[66]), 
            .\d10[67] (d10_adj_5723[67]), .\d10[68] (d10_adj_5723[68]), 
            .\d10[69] (d10_adj_5723[69]), .\d10[70] (d10_adj_5723[70]), 
            .\d10[71] (d10_adj_5723[71]), .\d_out_11__N_1819[2] (d_out_11__N_1819_adj_5748[2]), 
            .\d_out_11__N_1819[3] (d_out_11__N_1819_adj_5748[3]), .\d_out_11__N_1819[4] (d_out_11__N_1819_adj_5748[4]), 
            .\d_out_11__N_1819[5] (d_out_11__N_1819_adj_5748[5]), .\d_out_11__N_1819[6] (d_out_11__N_1819_adj_5748[6]), 
            .\d_out_11__N_1819[7] (d_out_11__N_1819_adj_5748[7]), .\d_out_11__N_1819[8] (d_out_11__N_1819_adj_5748[8]), 
            .\d_out_11__N_1819[9] (d_out_11__N_1819_adj_5748[9]), .\d_out_11__N_1819[10] (d_out_11__N_1819_adj_5748[10]), 
            .\d_out_11__N_1819[11] (d_out_11__N_1819_adj_5748[11]), .n11(n11_adj_4808), 
            .n17325(n17325), .n10_adj_117(n10_adj_4807), .n13_adj_118(n13_adj_4810), 
            .n12_adj_119(n12_adj_4809), .n15_adj_120(n15_adj_4812), .n14_adj_121(n14_adj_4811), 
            .n17_adj_122(n17_adj_4814), .n16_adj_123(n16_adj_4813), .n19(n19_adj_4816), 
            .n18(n18_adj_4815), .n21(n21_adj_4818), .n20(n20_adj_4817), 
            .n23_adj_124(n23_adj_4820), .n22_adj_125(n22_adj_4819), .n25(n25_adj_4822), 
            .n24(n24_adj_4821), .n27(n27_adj_4824), .n26(n26_adj_4823), 
            .n31(n31_adj_4746), .n30(n30_adj_4747), .n29(n29_adj_4826), 
            .n28(n28_adj_4825), .n17302(n17302), .n33(n33_adj_4733), .n31_adj_126(n31_adj_4828), 
            .n32(n32_adj_4745), .n30_adj_127(n30_adj_4827), .n33_adj_128(n33_adj_4830), 
            .n19_adj_129(n19_adj_4579), .n32_adj_130(n32_adj_4829), .n35_adj_131(n35_adj_4832), 
            .n35_adj_132(n35_adj_4735), .n34_adj_133(n34_adj_4734), .n18_adj_134(n18_adj_4580), 
            .n34_adj_135(n34_adj_4831), .n37_adj_136(n37_adj_4834), .n36_adj_137(n36_adj_4833), 
            .n3_adj_138(n3), .n2_adj_139(n2), .n5_adj_140(n5), .n37_adj_141(n37_adj_4737), 
            .n36_adj_142(n36_adj_4736), .n4_adj_143(n4), .n7_adj_144(n7), 
            .n6_adj_145(n6), .n9_adj_146(n9), .n8_adj_147(n8), .n11_adj_148(n11), 
            .n10_adj_149(n10), .n13_adj_150(n13), .n12_adj_151(n12), .n15_adj_152(n15), 
            .n14_adj_153(n14), .n17_adj_154(n17), .n16_adj_155(n16), .n19_adj_156(n19), 
            .n18_adj_157(n18), .n21_adj_158(n21), .n20_adj_159(n20), .n23_adj_160(n23), 
            .n22_adj_161(n22), .n25_adj_162(n25), .n24_adj_163(n24), .n27_adj_164(n27), 
            .n26_adj_165(n26), .n29_adj_166(n29), .n28_adj_167(n28), .n31_adj_168(n31), 
            .n30_adj_169(n30), .n33_adj_170(n33), .n5_adj_171(n5_adj_4759), 
            .n4_adj_172(n4_adj_4760), .n7_adj_173(n7_adj_4757), .n6_adj_174(n6_adj_4758), 
            .n3_adj_175(n3_adj_4761), .n2_adj_176(n2_adj_4762), .n3_adj_177(n3_adj_4764), 
            .n2_adj_178(n2_adj_4763), .n13_adj_179(n13_adj_4774), .n12_adj_180(n12_adj_4773), 
            .n15_adj_181(n15_adj_4776), .n14_adj_182(n14_adj_4775), .n32_adj_183(n32), 
            .n35_adj_184(n35), .n34_adj_185(n34), .n118(n118_adj_5591), 
            .n120(n120_adj_5000), .cout(cout_adj_2808), .n115(n115_adj_5590), 
            .n117(n117_adj_4999), .n112(n112_adj_5589), .n114(n114_adj_4998), 
            .n109(n109_adj_5588), .n111(n111_adj_4997), .n106(n106_adj_5587), 
            .n108(n108_adj_4996), .n17_adj_186(n17_adj_4778), .n103(n103_adj_5586), 
            .n105(n105_adj_4995), .n100(n100_adj_5585), .n102(n102_adj_4994), 
            .n97(n97_adj_5584), .n99(n99_adj_4993), .n94(n94_adj_5583), 
            .n96(n96_adj_4992), .n5_adj_187(n5_adj_4766), .n91(n91_adj_5582), 
            .n93(n93_adj_4991), .n16_adj_188(n16_adj_4777), .n19_adj_189(n19_adj_4780), 
            .n18_adj_190(n18_adj_4779), .n88(n88_adj_5581), .n90(n90_adj_4990), 
            .n21_adj_191(n21_adj_4782), .n20_adj_192(n20_adj_4781), .n23_adj_193(n23_adj_4784), 
            .n22_adj_194(n22_adj_4783), .n25_adj_195(n25_adj_4786), .n24_adj_196(n24_adj_4785), 
            .n27_adj_197(n27_adj_4788), .n26_adj_198(n26_adj_4787), .n25_adj_199(n25_adj_2798), 
            .n4_adj_200(n4_adj_4765), .n7_adj_201(n7_adj_4768), .n29_adj_202(n29_adj_4790), 
            .n21_adj_203(n21_adj_4577), .n28_adj_204(n28_adj_4789), .\CICGain[0] (CICGain[0]), 
            .n85(n85_adj_5580), .n87(n87_adj_4989), .n82(n82_adj_5579), 
            .n84(n84_adj_4988), .n20_adj_205(n20_adj_4578), .n31_adj_206(n31_adj_4792), 
            .n6_adj_207(n6_adj_4767), .n30_adj_208(n30_adj_4791), .n27_adj_209(n27_adj_4750), 
            .n26_adj_210(n26_adj_2797), .n29_adj_211(n29_adj_4748), .n28_adj_212(n28_adj_4749), 
            .n79(n79_adj_5578), .n81_adj_213(n81_adj_4987), .n9_adj_214(n9_adj_4770), 
            .n9_adj_215(n9_adj_4755), .n8_adj_216(n8_adj_4756), .n76(n76_adj_5577), 
            .n78_adj_217(n78_adj_4986), .n32_adj_218(n32_adj_4793), .n33_adj_219(n33_adj_4794), 
            .n63_adj_220(n63_adj_4740), .n11_adj_221(n11_adj_4753), .n17288(n17288), 
            .n65(n65), .n8_adj_222(n8_adj_4769), .n66_adj_223(n66_adj_4741), 
            .n11_adj_224(n11_adj_4772), .n37_adj_225(n37), .n36_adj_226(n36), 
            .n24_adj_227(n24_adj_4556)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(148[4] 154[5])
    PFUMX i2668 (.BLUT(n11984), .ALUT(n12255), .C0(n17389), .Z(n12573));
    LUT4 mux_339_i32_4_lut (.A(n3920), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2682)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i32_4_lut.init = 16'hc0ca;
    LUT4 i2077_3_lut (.A(n11970), .B(n283), .C(led_c_4), .Z(n11971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2077_3_lut.init = 16'hcaca;
    LUT4 mux_305_i58_4_lut_4_lut (.A(n17822), .B(n12538), .C(n8_adj_4726), 
         .D(n152), .Z(n1937)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam mux_305_i58_4_lut_4_lut.init = 16'h5410;
    LUT4 mux_305_i53_4_lut_4_lut (.A(n17822), .B(n12538), .C(n8_adj_4729), 
         .D(n167), .Z(n1942)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam mux_305_i53_4_lut_4_lut.init = 16'h5410;
    LUT4 i2646_3_lut (.A(n293), .B(n2703), .C(n12538), .Z(n12551)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2646_3_lut.init = 16'hacac;
    \CIC(WIDTH=72,DECIMATION_RATIO=4096)_U0  CIC_Sin_inst (.d_d7({d_d7}), 
            .n15(n15_adj_4640), .d_tmp({d_tmp}), .clk_80mhz(clk_80mhz), 
            .d5({d5}), .d_d_tmp({d_d_tmp}), .d2({d2}), .d2_71__N_490({d2_71__N_490}), 
            .n13(n13_adj_4714), .n12(n12_adj_4715), .n14(n14_adj_4641), 
            .d3({d3}), .d3_71__N_562({d3_71__N_562}), .count({count}), 
            .n87_adj_114({n36_adj_2807, n39_adj_2806, n42_adj_2805, n45_adj_2804, 
            n48_adj_2803, n51_adj_2802, n54_adj_2801, n57_adj_2800, 
            n60_adj_2799, n63, n66, n69, n72, n75, n78, n81}), 
            .d4({d4}), .d4_71__N_634({d4_71__N_634}), .d5_71__N_706({d5_71__N_706}), 
            .d6({d6}), .d6_71__N_1459({d6_71__N_1459}), .d_d6({d_d6}), 
            .CIC1_out_clkSin(CIC1_out_clkSin), .d7({d7}), .d7_71__N_1531({d7_71__N_1531}), 
            .d8({d8}), .d8_71__N_1603({d8_71__N_1603}), .d_d8({d_d8}), 
            .d9({d9}), .d9_71__N_1675({d9_71__N_1675}), .d_d9({d_d9}), 
            .n17(n17_adj_4638), .MultDataB({MultDataB}), .d1({d1}), .d1_71__N_418({d1_71__N_418}), 
            .n16(n16_adj_4639), .n15_adj_1(n15_adj_4712), .n19(n19_adj_4636), 
            .n14_adj_2(n14_adj_4713), .n17_adj_3(n17_adj_4710), .n16_adj_4(n16_adj_4711), 
            .n18(n18_adj_4637), .n19_adj_5(n19_adj_4708), .n21(n21_adj_4634), 
            .n20(n20_adj_4635), .n18_adj_6(n18_adj_4709), .n23(n23_adj_4632), 
            .n22(n22_adj_4633), .n21_adj_7(n21_adj_4706), .n25(n25_adj_4630), 
            .n24(n24_adj_4631), .n27(n27_adj_4628), .n20_adj_8(n20_adj_4707), 
            .n23_adj_9(n23_adj_4704), .n22_adj_10(n22_adj_4705), .n26(n26_adj_4629), 
            .n29(n29_adj_4626), .n25_adj_11(n25_adj_4702), .n28(n28_adj_4627), 
            .n24_adj_12(n24_adj_4703), .n27_adj_13(n27_adj_4700), .n26_adj_14(n26_adj_4701), 
            .n31(n31_adj_4624), .n29_adj_15(n29_adj_4698), .n28_adj_16(n28_adj_4699), 
            .n31_adj_17(n31_adj_4696), .n30(n30_adj_4697), .n30_adj_18(n30_adj_4625), 
            .n33(n33_adj_4622), .n32(n32_adj_4623), .n33_adj_19(n33_adj_4694), 
            .n32_adj_20(n32_adj_4695), .n35(n35_adj_4692), .n34(n34_adj_4693), 
            .n35_adj_21(n35_adj_4620), .n37(n37_adj_4690), .n36_adj_22(n36_adj_4691), 
            .n34_adj_23(n34_adj_4621), .n37_adj_24(n37_adj_4618), .n36_adj_25(n36_adj_4619), 
            .\CICGain[1] (CICGain[1]), .\CICGain[0] (CICGain[0]), .\d10[66] (d10_adj_5723[66]), 
            .\d10[67] (d10_adj_5723[67]), .\d10[69] (d10_adj_5723[69]), 
            .\d10[68] (d10_adj_5723[68]), .n3(n3_adj_4688), .n2(n2_adj_4689), 
            .\d10[65] (d10_adj_5723[65]), .n5(n5_adj_4686), .\d10[70] (d10_adj_5723[70]), 
            .n4(n4_adj_4687), .\d10[71] (d10_adj_5723[71]), .n7(n7_adj_4684), 
            .n6(n6_adj_4685), .n9(n9_adj_4682), .n8(n8_adj_4683), .n11(n11_adj_4680), 
            .n10(n10_adj_4681), .n13_adj_26(n13_adj_4678), .n118(n118), 
            .n120(n120), .cout(cout_adj_5462), .n115(n115), .n117(n117), 
            .n112(n112), .n114(n114), .n3_adj_27(n3_adj_4616), .n109(n109), 
            .n111(n111), .n2_adj_28(n2_adj_4617), .n5_adj_29(n5_adj_4614), 
            .n63_adj_30(n63_adj_4740), .\d_out_11__N_1819[2] (d_out_11__N_1819_adj_5748[2]), 
            .n4_adj_31(n4_adj_4615), .n12_adj_32(n12_adj_4679), .n7_adj_33(n7_adj_4612), 
            .n6_adj_34(n6_adj_4613), .n9_adj_35(n9_adj_4610), .n17288(n17288), 
            .\d_out_11__N_1819[3] (d_out_11__N_1819_adj_5748[3]), .n65(n65), 
            .\d_out_11__N_1819[4] (d_out_11__N_1819_adj_5748[4]), .n8_adj_36(n8_adj_4611), 
            .n66_adj_37(n66_adj_4741), .\d_out_11__N_1819[5] (d_out_11__N_1819_adj_5748[5]), 
            .n11_adj_38(n11_adj_4608), .\d_out_11__N_1819[6] (d_out_11__N_1819_adj_5748[6]), 
            .n10_adj_39(n10_adj_4609), .n13_adj_40(n13_adj_4606), .n12_adj_41(n12_adj_4607), 
            .n15_adj_42(n15_adj_4676), .n15_adj_43(n15_adj_4604), .n14_adj_44(n14_adj_4677), 
            .\d_out_11__N_1819[7] (d_out_11__N_1819_adj_5748[7]), .n14_adj_45(n14_adj_4605), 
            .n17_adj_46(n17_adj_4602), .n106(n106), .n108(n108), .n16_adj_47(n16_adj_4603), 
            .n17_adj_48(n17_adj_4674), .n16_adj_49(n16_adj_4675), .n19_adj_50(n19_adj_4672), 
            .n18_adj_51(n18_adj_4673), .n21_adj_52(n21_adj_4670), .n20_adj_53(n20_adj_4671), 
            .n23_adj_54(n23_adj_4668), .n22_adj_55(n22_adj_4669), .n25_adj_56(n25_adj_4666), 
            .n24_adj_57(n24_adj_4667), .n27_adj_58(n27_adj_4664), .n26_adj_59(n26_adj_4665), 
            .n29_adj_60(n29_adj_4662), .n28_adj_61(n28_adj_4663), .n31_adj_62(n31_adj_4660), 
            .n30_adj_63(n30_adj_4661), .n33_adj_64(n33_adj_4658), .n32_adj_65(n32_adj_4659), 
            .n35_adj_66(n35_adj_4656), .n34_adj_67(n34_adj_4657), .n37_adj_68(n37_adj_4654), 
            .n36_adj_69(n36_adj_4655), .n19_adj_70(n19_adj_4600), .n18_adj_71(n18_adj_4601), 
            .n21_adj_72(n21_adj_4598), .n20_adj_73(n20_adj_4599), .n23_adj_74(n23_adj_4596), 
            .n22_adj_75(n22_adj_4597), .n25_adj_76(n25_adj_4593), .n24_adj_77(n24_adj_4594), 
            .n27_adj_78(n27_adj_4591), .n26_adj_79(n26_adj_4592), .n29_adj_80(n29_adj_4589), 
            .n28_adj_81(n28_adj_4590), .n31_adj_82(n31_adj_4587), .n30_adj_83(n30_adj_4588), 
            .n33_adj_84(n33_adj_4585), .n32_adj_85(n32_adj_4586), .n35_adj_86(n35_adj_4583), 
            .n34_adj_87(n34_adj_4584), .n37_adj_88(n37_adj_4581), .n36_adj_89(n36_adj_4582), 
            .n103(n103), .n105(n105), .n3_adj_90(n3_adj_4652), .n2_adj_91(n2_adj_4653), 
            .n100(n100), .n102(n102), .n97(n97), .n99(n99), .n5_adj_92(n5_adj_4650), 
            .n4_adj_93(n4_adj_4651), .n7_adj_94(n7_adj_4648), .n6_adj_95(n6_adj_4649), 
            .n9_adj_96(n9_adj_4646), .n94(n94), .n96(n96), .n8_adj_97(n8_adj_4647), 
            .n91(n91), .n93(n93), .n11_adj_98(n11_adj_4644), .n10_adj_99(n10_adj_4645), 
            .n13_adj_100(n13_adj_4642), .n12_adj_101(n12_adj_4643), .n88(n88), 
            .n90(n90), .n85(n85), .n87(n87), .n82(n82), .n84(n84), 
            .n79(n79), .n81_adj_102(n81_adj_4559), .n76(n76), .n78_adj_103(n78_adj_4560), 
            .\d10[63] (d10_adj_5723[63]), .\d10[64] (d10_adj_5723[64]), 
            .\d10[62] (d10_adj_5723[62]), .n17325(n17325), .\d10[60] (d10_adj_5723[60]), 
            .\d10[61] (d10_adj_5723[61]), .n17302(n17302), .\d10[59] (d10_adj_5723[59]), 
            .\d_out_11__N_1819[10] (d_out_11__N_1819_adj_5748[10]), .\d_out_11__N_1819[11] (d_out_11__N_1819_adj_5748[11]), 
            .\d_out_11__N_1819[8] (d_out_11__N_1819_adj_5748[8]), .\d_out_11__N_1819[9] (d_out_11__N_1819_adj_5748[9]), 
            .n3_adj_104(n3_adj_4724), .n2_adj_105(n2_adj_4725), .n5_adj_106(n5_adj_4722), 
            .n4_adj_107(n4_adj_4723), .n7_adj_108(n7_adj_4720), .n6_adj_109(n6_adj_4721), 
            .n9_adj_110(n9_adj_4718), .n8_adj_111(n8_adj_4719), .n11_adj_112(n11_adj_4716), 
            .n10_adj_113(n10_adj_4717)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(136[4] 142[5])
    LUT4 mux_339_i11_4_lut (.A(n3941), .B(led_c_1), .C(n17813), .D(n17812), 
         .Z(n2703)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_339_i11_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1454_add_4_3 (.A0(d4[36]), .B0(cout_adj_2810), .C0(n183_adj_5320), 
          .D0(d5[36]), .A1(d4[37]), .B1(cout_adj_2810), .C1(n180_adj_5319), 
          .D1(d5[37]), .CIN(n16044), .COUT(n16045), .S0(d5_71__N_706[36]), 
          .S1(d5_71__N_706[37]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1454_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1454_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1454_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1454_add_4_3.INJECT1_1 = "NO";
    LUT4 mux_843_i10_3_lut (.A(n283_adj_5075), .B(n289), .C(led_c_4), 
         .Z(n3941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam mux_843_i10_3_lut.init = 16'hcaca;
    LUT4 i2644_4_lut (.A(n296), .B(n11969), .C(n12538), .D(n17813), 
         .Z(n12549)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2644_4_lut.init = 16'hafac;
    LUT4 i2075_3_lut (.A(n11968), .B(n292), .C(n18053), .Z(n11969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(191[6] 213[10])
    defparam i2075_3_lut.init = 16'hcaca;
    PFUMX i6094 (.BLUT(n17836), .ALUT(n17837), .C0(led_c_0), .Z(n12424));
    AMDemodulator AMDemodulator_inst (.\DataInReg_11__N_1856[0] (DataInReg_11__N_1856[0]), 
            .CIC1_out_clkSin(CIC1_out_clkSin), .CIC1_outCos({CIC1_outCos}), 
            .MultResult2({MultResult2}), .\d_out_d_11__N_1874[17] (d_out_d_11__N_1874[17]), 
            .d_out_d_11__N_1873(d_out_d_11__N_1873), .MultDataB({MultDataB}), 
            .MultResult1({MultResult1}), .VCC_net(VCC_net), .GND_net(GND_net), 
            .\DataInReg_11__N_1856[1] (DataInReg_11__N_1856[1]), .\DataInReg_11__N_1856[2] (DataInReg_11__N_1856[2]), 
            .\DataInReg_11__N_1856[3] (DataInReg_11__N_1856[3]), .\DataInReg_11__N_1856[4] (DataInReg_11__N_1856[4]), 
            .\DataInReg_11__N_1856[5] (DataInReg_11__N_1856[5]), .\DataInReg_11__N_1856[6] (DataInReg_11__N_1856[6]), 
            .\DataInReg_11__N_1856[7] (DataInReg_11__N_1856[7]), .\DataInReg_11__N_1856[8] (DataInReg_11__N_1856[8]), 
            .\DemodOut[9] (DemodOut[9]), .\ISquare[31] (ISquare[31]), .n213(n213), 
            .\d_out_d_11__N_1892[17] (d_out_d_11__N_1892[17]), .\d_out_d_11__N_1890[17] (d_out_d_11__N_1890[17]), 
            .\d_out_d_11__N_1888[17] (d_out_d_11__N_1888[17]), .\d_out_d_11__N_1886[17] (d_out_d_11__N_1886[17]), 
            .\d_out_d_11__N_1884[17] (d_out_d_11__N_1884[17]), .\d_out_d_11__N_1882[17] (d_out_d_11__N_1882[17]), 
            .\d_out_d_11__N_1878[17] (d_out_d_11__N_1878[17]), .d_out_d_11__N_1877(d_out_d_11__N_1877), 
            .\d_out_d_11__N_1876[17] (d_out_d_11__N_1876[17]), .d_out_d_11__N_1875(d_out_d_11__N_1875), 
            .d_out_d_11__N_1879(d_out_d_11__N_1879), .\d_out_d_11__N_2383[17] (d_out_d_11__N_2383[17]), 
            .\d_out_d_11__N_2401[17] (d_out_d_11__N_2401[17]), .\d_out_d_11__N_1880[17] (d_out_d_11__N_1880[17])) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(171[18] 176[5])
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=87) 
//

module \uart_rx(CLKS_PER_BIT=87)  (clk_80mhz, i_Rx_Serial_c, o_Rx_Byte1, 
            o_Rx_DV1, GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input clk_80mhz;
    input i_Rx_Serial_c;
    output [7:0]o_Rx_Byte1;
    output o_Rx_DV1;
    input GND_net;
    input VCC_net;
    
    wire [7:0]UartClk /* synthesis SET_AS_NETWORK=\uart_rx_inst/UartClk[2], is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(37[14:21])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(61[23:32])
    wire [2:0]r_SM_Main;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(43[17:26])
    
    wire n17344, r_Rx_DV_last, r_Rx_DV, r_Rx_Data_R, r_Rx_Data, UartClk_2_enable_27;
    wire [7:0]r_Rx_Byte;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(41[17:26])
    wire [15:0]r_Clock_Count;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(39[18:31])
    
    wire UartClk_2_enable_18, n12716;
    wire [15:0]n69;
    wire [2:0]r_Bit_Index;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(40[17:28])
    
    wire UartClk_2_enable_29, n17038, n17342, n17343;
    wire [2:0]n30;
    wire [2:0]n17;
    
    wire n16821, n13228, n17843, n17819, n17842, n17811, UartClk_2_enable_36, 
        UartClk_2_enable_20, n17123, n17824, UartClk_2_enable_21, n17844, 
        n17818, n13202, n17137, n17062, n17833, r_Rx_DV_N_2532, 
        n12714, r_Rx_DV_last_N_2531, n24, n17111, n16878, UartClk_2_enable_31, 
        n13004, UartClk_2_enable_30, n26, n16952, n15395, UartClk_2_enable_32, 
        UartClk_2_enable_33, n15821, n15820, n15819, n15818, n15817, 
        n15816, n15815, n15814, UartClk_2_enable_34, UartClk_2_enable_35, 
        n17113, n16570, n17101, n17103, n17095, n17099, n13208, 
        n17831, n16859;
    
    FD1S3IX r_SM_Main_i0 (.D(n17344), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i0.GSR = "ENABLED";
    FD1S3AX r_Rx_DV_last_60 (.D(r_Rx_DV), .CK(clk_80mhz), .Q(r_Rx_DV_last)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(47[11] 52[8])
    defparam r_Rx_DV_last_60.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_R_61 (.D(i_Rx_Serial_c), .CK(UartClk[2]), .Q(r_Rx_Data_R)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(57[11] 62[8])
    defparam r_Rx_Data_R_61.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_62 (.D(r_Rx_Data_R), .CK(UartClk[2]), .Q(r_Rx_Data)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(57[11] 62[8])
    defparam r_Rx_Data_62.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i0 (.D(r_Rx_Byte[0]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i0.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i0 (.D(n69[0]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i0.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i0 (.D(n17038), .SP(UartClk_2_enable_29), .CK(UartClk[2]), 
            .Q(r_Bit_Index[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i0.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i15 (.D(n69[15]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[15])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i15.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i14 (.D(n69[14]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[14])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i14.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i13 (.D(n69[13]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[13])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i13.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i12 (.D(n69[12]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[12])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i12.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i11 (.D(n69[11]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[11])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i11.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i10 (.D(n69[10]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[10])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i10.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i9 (.D(n69[9]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i9.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i8 (.D(n69[8]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i8.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i7 (.D(n69[7]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i7.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i6 (.D(n69[6]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i6.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i5 (.D(n69[5]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i5.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i4 (.D(n69[4]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i4.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i3 (.D(n69[3]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i3.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i2 (.D(n69[2]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i2.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_958__i1 (.D(n69[1]), .SP(UartClk_2_enable_18), 
            .CD(n12716), .CK(UartClk[2]), .Q(r_Clock_Count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958__i1.GSR = "ENABLED";
    PFUMX i5885 (.BLUT(n17342), .ALUT(n17343), .C0(r_SM_Main[1]), .Z(n17344));
    FD1S3AX UartClk_956_969__i0 (.D(n17[0]), .CK(clk_80mhz), .Q(n30[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_956_969__i0.GSR = "ENABLED";
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut (.A(r_SM_Main[0]), 
         .B(n16821), .C(n13228), .Z(n17843)) /* synthesis lut_function=(!(A (B+(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(69[7] 161[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut.init = 16'h5757;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut (.A(r_SM_Main[0]), 
         .B(n17819), .C(r_Rx_Data), .Z(n17842)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(69[7] 161[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut.init = 16'h0202;
    LUT4 i5969_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n17811), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_36)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(114[17:39])
    defparam i5969_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i5954_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n17811), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_20)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(114[17:39])
    defparam i5954_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i6029_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(n17819), 
         .D(n17123), .Z(UartClk_2_enable_18)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(69[7] 161[14])
    defparam i6029_4_lut.init = 16'h5455;
    LUT4 i1_2_lut (.A(r_Rx_Data), .B(r_SM_Main[0]), .Z(n17123)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(r_SM_Main[1]), .B(n17824), .C(r_Bit_Index[0]), 
         .D(r_SM_Main[0]), .Z(n17038)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0008;
    LUT4 i21_4_lut_4_lut (.A(r_SM_Main[1]), .B(n17824), .C(r_SM_Main[0]), 
         .D(r_SM_Main[2]), .Z(UartClk_2_enable_21)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (C))) */ ;
    defparam i21_4_lut_4_lut.init = 16'h0585;
    LUT4 i1_2_lut_rep_202 (.A(n13228), .B(n16821), .Z(n17824)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_202.init = 16'heeee;
    FD1S3IX r_SM_Main_i1 (.D(n17844), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i1.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i1 (.D(r_Rx_Byte[1]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    LUT4 i1_3_lut_rep_196_3_lut_4_lut (.A(n13228), .B(n16821), .C(r_SM_Main[1]), 
         .D(r_SM_Main[2]), .Z(n17818)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;
    defparam i1_3_lut_rep_196_3_lut_4_lut.init = 16'hff1f;
    LUT4 i5884_4_lut_3_lut_4_lut (.A(n13228), .B(n16821), .C(n13202), 
         .D(r_SM_Main[0]), .Z(n17343)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(D)))) */ ;
    defparam i5884_4_lut_3_lut_4_lut.init = 16'h11e0;
    LUT4 i1_3_lut_4_lut_adj_56 (.A(n13228), .B(n16821), .C(n13202), .D(n17137), 
         .Z(n17062)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i1_3_lut_4_lut_adj_56.init = 16'h0e00;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n13228), .B(n16821), .C(n17833), .D(r_SM_Main[0]), 
         .Z(r_Rx_DV_N_2532)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'he000;
    FD1S3IX o_Rx_DV_59 (.D(r_Rx_DV_last_N_2531), .CK(clk_80mhz), .CD(n12714), 
            .Q(o_Rx_DV1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(47[11] 52[8])
    defparam o_Rx_DV_59.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(r_SM_Main[2]), .B(n24), .C(n17824), .D(r_SM_Main[1]), 
         .Z(n12716)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i1_4_lut.init = 16'h5044;
    FD1P3AX r_Rx_Byte_i0 (.D(r_Rx_Data), .SP(UartClk_2_enable_20), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i0.GSR = "ENABLED";
    FD1P3AX r_Rx_DV_64 (.D(r_Rx_DV_N_2532), .SP(UartClk_2_enable_21), .CK(UartClk[2]), 
            .Q(r_Rx_DV)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_DV_64.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i2 (.D(r_Rx_Byte[2]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i3 (.D(r_Rx_Byte[3]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i4 (.D(r_Rx_Byte[4]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i5 (.D(r_Rx_Byte[5]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i6 (.D(r_Rx_Byte[6]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i7 (.D(r_Rx_Byte[7]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    LUT4 i5989_4_lut (.A(n17111), .B(n16821), .C(n13228), .D(r_SM_Main[1]), 
         .Z(UartClk_2_enable_29)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;
    defparam i5989_4_lut.init = 16'h5455;
    LUT4 i1_2_lut_adj_57 (.A(r_SM_Main[0]), .B(r_SM_Main[2]), .Z(n17111)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_57.init = 16'heeee;
    LUT4 i5982_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n17818), .C(n16878), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_31)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(114[17:39])
    defparam i5982_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i5984_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n17818), .C(n13004), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_30)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(114[17:39])
    defparam i5984_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_4_lut_adj_58 (.A(r_Bit_Index[2]), .B(r_SM_Main[0]), .C(n13004), 
         .D(r_SM_Main[1]), .Z(n17137)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_58.init = 16'h1200;
    LUT4 i3093_2_lut (.A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .Z(n13004)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3093_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_59 (.A(n26), .B(n17824), .C(r_SM_Main[0]), .D(r_SM_Main[1]), 
         .Z(n16952)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_59.init = 16'h0800;
    LUT4 i39_2_lut (.A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .Z(n26)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i39_2_lut.init = 16'h6666;
    CCU2C UartClk_956_969_add_4_3 (.A0(n30[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(UartClk[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15395), .S0(n17[1]), .S1(n17[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_956_969_add_4_3.INIT0 = 16'haaa0;
    defparam UartClk_956_969_add_4_3.INIT1 = 16'haaa0;
    defparam UartClk_956_969_add_4_3.INJECT1_0 = "NO";
    defparam UartClk_956_969_add_4_3.INJECT1_1 = "NO";
    CCU2C UartClk_956_969_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15395), .S1(n17[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_956_969_add_4_1.INIT0 = 16'h0000;
    defparam UartClk_956_969_add_4_1.INIT1 = 16'h555f;
    defparam UartClk_956_969_add_4_1.INJECT1_0 = "NO";
    defparam UartClk_956_969_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_60 (.A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .Z(n16878)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(114[17:39])
    defparam i1_2_lut_adj_60.init = 16'hbbbb;
    FD1P3AX r_Bit_Index_i2 (.D(n17062), .SP(UartClk_2_enable_29), .CK(UartClk[2]), 
            .Q(r_Bit_Index[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i2.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i1 (.D(n16952), .SP(UartClk_2_enable_29), .CK(UartClk[2]), 
            .Q(r_Bit_Index[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i1.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i7 (.D(r_Rx_Data), .SP(UartClk_2_enable_30), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i7.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i6 (.D(r_Rx_Data), .SP(UartClk_2_enable_31), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i5 (.D(r_Rx_Data), .SP(UartClk_2_enable_32), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i4 (.D(r_Rx_Data), .SP(UartClk_2_enable_33), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i4.GSR = "ENABLED";
    CCU2C r_Clock_Count_958_add_4_17 (.A0(r_Clock_Count[15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15821), .S0(n69[15]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958_add_4_17.INIT0 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_17.INIT1 = 16'h0000;
    defparam r_Clock_Count_958_add_4_17.INJECT1_0 = "NO";
    defparam r_Clock_Count_958_add_4_17.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_958_add_4_15 (.A0(r_Clock_Count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15820), .COUT(n15821), .S0(n69[13]), 
          .S1(n69[14]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958_add_4_15.INIT0 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_15.INIT1 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_15.INJECT1_0 = "NO";
    defparam r_Clock_Count_958_add_4_15.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_958_add_4_13 (.A0(r_Clock_Count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15819), .COUT(n15820), .S0(n69[11]), 
          .S1(n69[12]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958_add_4_13.INIT0 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_13.INIT1 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_13.INJECT1_0 = "NO";
    defparam r_Clock_Count_958_add_4_13.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_958_add_4_11 (.A0(r_Clock_Count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15818), .COUT(n15819), .S0(n69[9]), 
          .S1(n69[10]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958_add_4_11.INIT0 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_11.INIT1 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_11.INJECT1_0 = "NO";
    defparam r_Clock_Count_958_add_4_11.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_958_add_4_9 (.A0(r_Clock_Count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15817), .COUT(n15818), .S0(n69[7]), 
          .S1(n69[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958_add_4_9.INIT0 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_9.INIT1 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_9.INJECT1_0 = "NO";
    defparam r_Clock_Count_958_add_4_9.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_958_add_4_7 (.A0(r_Clock_Count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15816), .COUT(n15817), .S0(n69[5]), 
          .S1(n69[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958_add_4_7.INIT0 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_7.INIT1 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_7.INJECT1_0 = "NO";
    defparam r_Clock_Count_958_add_4_7.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_958_add_4_5 (.A0(r_Clock_Count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15815), .COUT(n15816), .S0(n69[3]), 
          .S1(n69[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958_add_4_5.INIT0 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_5.INIT1 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_5.INJECT1_0 = "NO";
    defparam r_Clock_Count_958_add_4_5.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_958_add_4_3 (.A0(r_Clock_Count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15814), .COUT(n15815), .S0(n69[1]), 
          .S1(n69[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958_add_4_3.INIT0 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_3.INIT1 = 16'haaa0;
    defparam r_Clock_Count_958_add_4_3.INJECT1_0 = "NO";
    defparam r_Clock_Count_958_add_4_3.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_958_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(r_Clock_Count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15814), .S1(n69[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_958_add_4_1.INIT0 = 16'h0000;
    defparam r_Clock_Count_958_add_4_1.INIT1 = 16'h555f;
    defparam r_Clock_Count_958_add_4_1.INJECT1_0 = "NO";
    defparam r_Clock_Count_958_add_4_1.INJECT1_1 = "NO";
    FD1P3AX r_Rx_Byte_i3 (.D(r_Rx_Data), .SP(UartClk_2_enable_34), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i3.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i2 (.D(r_Rx_Data), .SP(UartClk_2_enable_35), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i2.GSR = "ENABLED";
    FD1S3AX UartClk_956_969__i1 (.D(n17[1]), .CK(clk_80mhz), .Q(n30[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_956_969__i1.GSR = "ENABLED";
    FD1S3AX UartClk_956_969__i2 (.D(n17[2]), .CK(clk_80mhz), .Q(UartClk[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_956_969__i2.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(r_Bit_Index[1]), .B(r_Bit_Index[0]), .C(r_Bit_Index[2]), 
         .Z(n13202)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_61 (.A(r_Clock_Count[1]), .B(n16821), .C(n17113), 
         .D(r_Clock_Count[6]), .Z(n16570)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(85[17:52])
    defparam i1_4_lut_adj_61.init = 16'hfffd;
    LUT4 i1_2_lut_adj_62 (.A(r_Clock_Count[2]), .B(r_Clock_Count[4]), .Z(n17113)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_62.init = 16'heeee;
    LUT4 i1_4_lut_adj_63 (.A(n17101), .B(n17103), .C(n17095), .D(n17099), 
         .Z(n16821)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(85[17:52])
    defparam i1_4_lut_adj_63.init = 16'hfffe;
    LUT4 i1_2_lut_adj_64 (.A(r_Clock_Count[11]), .B(r_Clock_Count[15]), 
         .Z(n17101)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_64.init = 16'heeee;
    LUT4 i1_3_lut_adj_65 (.A(r_Clock_Count[13]), .B(r_Clock_Count[8]), .C(r_Clock_Count[7]), 
         .Z(n17103)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(85[17:52])
    defparam i1_3_lut_adj_65.init = 16'hfefe;
    LUT4 i1_2_lut_adj_66 (.A(r_Clock_Count[14]), .B(r_Clock_Count[10]), 
         .Z(n17095)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_66.init = 16'heeee;
    LUT4 i1_2_lut_adj_67 (.A(r_Clock_Count[9]), .B(r_Clock_Count[12]), .Z(n17099)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_67.init = 16'heeee;
    LUT4 i5979_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n17811), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_32)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(114[17:39])
    defparam i5979_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i3317_4_lut (.A(n13208), .B(r_Clock_Count[6]), .C(r_Clock_Count[5]), 
         .D(r_Clock_Count[4]), .Z(n13228)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i3317_4_lut.init = 16'hc8c0;
    LUT4 i3297_3_lut (.A(r_Clock_Count[1]), .B(r_Clock_Count[3]), .C(r_Clock_Count[2]), 
         .Z(n13208)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i3297_3_lut.init = 16'hecec;
    LUT4 i5977_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n17811), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_33)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(114[17:39])
    defparam i5977_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i2803_1_lut (.A(r_Rx_DV), .Z(n12714)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i2803_1_lut.init = 16'h5555;
    LUT4 r_Rx_DV_last_I_0_1_lut (.A(r_Rx_DV_last), .Z(r_Rx_DV_last_N_2531)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(50[30:43])
    defparam r_Rx_DV_last_I_0_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_rep_189_4_lut_4_lut (.A(n17824), .B(r_SM_Main[0]), .C(r_SM_Main[2]), 
         .D(r_SM_Main[1]), .Z(n17811)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i1_2_lut_rep_189_4_lut_4_lut.init = 16'hfdff;
    LUT4 i6031_2_lut_4_lut_4_lut (.A(n17824), .B(r_SM_Main[0]), .C(r_SM_Main[2]), 
         .D(r_SM_Main[1]), .Z(UartClk_2_enable_27)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i6031_2_lut_4_lut_4_lut.init = 16'h0800;
    LUT4 i5972_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n17818), .C(n16878), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_35)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(114[17:39])
    defparam i5972_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_3_lut_rep_209 (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), .C(r_Clock_Count[0]), 
         .Z(n17831)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_rep_209.init = 16'h8080;
    LUT4 i1_2_lut_rep_197_4_lut (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), 
         .C(r_Clock_Count[0]), .D(n16570), .Z(n17819)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_197_4_lut.init = 16'hff7f;
    LUT4 i5883_3_lut_4_lut_4_lut (.A(r_Rx_Data), .B(r_SM_Main[0]), .C(n16570), 
         .D(n17831), .Z(n17342)) /* synthesis lut_function=(A (B (C+!(D)))+!A ((C+!(D))+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(87[21:38])
    defparam i5883_3_lut_4_lut_4_lut.init = 16'hd1dd;
    LUT4 i1_4_lut_4_lut (.A(r_Rx_Data), .B(n17831), .C(n16570), .D(r_SM_Main[0]), 
         .Z(n24)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(87[21:38])
    defparam i1_4_lut_4_lut.init = 16'h04ff;
    LUT4 i1_2_lut_rep_211 (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .Z(n17833)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(69[7] 161[14])
    defparam i1_2_lut_rep_211.init = 16'h2222;
    LUT4 i5967_2_lut_3_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .Z(n16859)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(69[7] 161[14])
    defparam i5967_2_lut_3_lut.init = 16'hdfdf;
    LUT4 i5974_2_lut_3_lut_4_lut (.A(r_SM_Main[0]), .B(n17818), .C(n13004), 
         .D(r_Bit_Index[2]), .Z(UartClk_2_enable_34)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(114[17:39])
    defparam i5974_2_lut_3_lut_4_lut.init = 16'h0010;
    FD1P3AX r_Rx_Byte_i1 (.D(r_Rx_Data), .SP(UartClk_2_enable_36), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i1.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i2 (.D(n17824), .CK(UartClk[2]), .CD(n16859), .Q(r_SM_Main[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i2.GSR = "ENABLED";
    PFUMX i6098 (.BLUT(n17842), .ALUT(n17843), .C0(r_SM_Main[1]), .Z(n17844));
    
endmodule
//
// Verilog Description of module Mixer
//

module Mixer (MixerOutSin, clk_80mhz, DiffOut_c, MixerOutCos, RFIn_c, 
            \LOSine[1] , MixerOutSin_11__N_236, \LOCosine[1] , MixerOutCos_11__N_250, 
            \LOSine[6] , \LOSine[11] , \LOSine[10] , \LOSine[9] , \LOSine[5] , 
            \LOSine[4] , \LOSine[8] , \LOSine[7] , \LOSine[3] , \LOSine[2] , 
            \LOCosine[12] , \LOCosine[11] , \LOCosine[10] , \LOCosine[9] , 
            \LOCosine[8] , \LOCosine[7] , \LOCosine[6] , \LOCosine[5] , 
            \LOCosine[4] , \LOCosine[3] , \LOCosine[2] , \LOSine[12] ) /* synthesis syn_module_defined=1 */ ;
    output [11:0]MixerOutSin;
    input clk_80mhz;
    output DiffOut_c;
    output [11:0]MixerOutCos;
    input RFIn_c;
    input \LOSine[1] ;
    input [11:0]MixerOutSin_11__N_236;
    input \LOCosine[1] ;
    input [11:0]MixerOutCos_11__N_250;
    input \LOSine[6] ;
    input \LOSine[11] ;
    input \LOSine[10] ;
    input \LOSine[9] ;
    input \LOSine[5] ;
    input \LOSine[4] ;
    input \LOSine[8] ;
    input \LOSine[7] ;
    input \LOSine[3] ;
    input \LOSine[2] ;
    input \LOCosine[12] ;
    input \LOCosine[11] ;
    input \LOCosine[10] ;
    input \LOCosine[9] ;
    input \LOCosine[8] ;
    input \LOCosine[7] ;
    input \LOCosine[6] ;
    input \LOCosine[5] ;
    input \LOCosine[4] ;
    input \LOCosine[3] ;
    input \LOCosine[2] ;
    input \LOSine[12] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(61[23:32])
    wire [11:0]MixerOutSin_11__N_212;
    
    wire RFInR;
    wire [11:0]MixerOutCos_11__N_224;
    
    FD1S3AX MixerOutSin_i0 (.D(MixerOutSin_11__N_212[0]), .CK(clk_80mhz), 
            .Q(MixerOutSin[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i0.GSR = "ENABLED";
    FD1S3AY RFInR_14 (.D(DiffOut_c), .CK(clk_80mhz), .Q(RFInR)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(34[10] 37[6])
    defparam RFInR_14.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i0 (.D(MixerOutCos_11__N_224[0]), .CK(clk_80mhz), 
            .Q(MixerOutCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i0.GSR = "ENABLED";
    FD1S3AY RFInR1_13 (.D(RFIn_c), .CK(clk_80mhz), .Q(DiffOut_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(34[10] 37[6])
    defparam RFInR1_13.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i11 (.D(MixerOutCos_11__N_224[11]), .CK(clk_80mhz), 
            .Q(MixerOutCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i11.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i10 (.D(MixerOutCos_11__N_224[10]), .CK(clk_80mhz), 
            .Q(MixerOutCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i10.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i9 (.D(MixerOutCos_11__N_224[9]), .CK(clk_80mhz), 
            .Q(MixerOutCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i9.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i8 (.D(MixerOutCos_11__N_224[8]), .CK(clk_80mhz), 
            .Q(MixerOutCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i8.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i7 (.D(MixerOutCos_11__N_224[7]), .CK(clk_80mhz), 
            .Q(MixerOutCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i7.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i6 (.D(MixerOutCos_11__N_224[6]), .CK(clk_80mhz), 
            .Q(MixerOutCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i6.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i5 (.D(MixerOutCos_11__N_224[5]), .CK(clk_80mhz), 
            .Q(MixerOutCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i5.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i4 (.D(MixerOutCos_11__N_224[4]), .CK(clk_80mhz), 
            .Q(MixerOutCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i4.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i3 (.D(MixerOutCos_11__N_224[3]), .CK(clk_80mhz), 
            .Q(MixerOutCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i3.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i2 (.D(MixerOutCos_11__N_224[2]), .CK(clk_80mhz), 
            .Q(MixerOutCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i2.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i1 (.D(MixerOutCos_11__N_224[1]), .CK(clk_80mhz), 
            .Q(MixerOutCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i1.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i11 (.D(MixerOutSin_11__N_212[11]), .CK(clk_80mhz), 
            .Q(MixerOutSin[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i11.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i10 (.D(MixerOutSin_11__N_212[10]), .CK(clk_80mhz), 
            .Q(MixerOutSin[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i10.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i9 (.D(MixerOutSin_11__N_212[9]), .CK(clk_80mhz), 
            .Q(MixerOutSin[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i9.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i8 (.D(MixerOutSin_11__N_212[8]), .CK(clk_80mhz), 
            .Q(MixerOutSin[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i8.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i7 (.D(MixerOutSin_11__N_212[7]), .CK(clk_80mhz), 
            .Q(MixerOutSin[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i7.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i6 (.D(MixerOutSin_11__N_212[6]), .CK(clk_80mhz), 
            .Q(MixerOutSin[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i6.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i5 (.D(MixerOutSin_11__N_212[5]), .CK(clk_80mhz), 
            .Q(MixerOutSin[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i5.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i4 (.D(MixerOutSin_11__N_212[4]), .CK(clk_80mhz), 
            .Q(MixerOutSin[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i4.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i3 (.D(MixerOutSin_11__N_212[3]), .CK(clk_80mhz), 
            .Q(MixerOutSin[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i3.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i2 (.D(MixerOutSin_11__N_212[2]), .CK(clk_80mhz), 
            .Q(MixerOutSin[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i2.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i1 (.D(MixerOutSin_11__N_212[1]), .CK(clk_80mhz), 
            .Q(MixerOutSin[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i1.GSR = "ENABLED";
    LUT4 MixerOutSin_11__I_0_i1_3_lut (.A(\LOSine[1] ), .B(MixerOutSin_11__N_236[0]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i1_3_lut (.A(\LOCosine[1] ), .B(MixerOutCos_11__N_250[0]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i6_3_lut (.A(\LOSine[6] ), .B(MixerOutSin_11__N_236[5]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i11_3_lut (.A(\LOSine[11] ), .B(MixerOutSin_11__N_236[10]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i10_3_lut (.A(\LOSine[10] ), .B(MixerOutSin_11__N_236[9]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i9_3_lut (.A(\LOSine[9] ), .B(MixerOutSin_11__N_236[8]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i5_3_lut (.A(\LOSine[5] ), .B(MixerOutSin_11__N_236[4]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i4_3_lut (.A(\LOSine[4] ), .B(MixerOutSin_11__N_236[3]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i8_3_lut (.A(\LOSine[8] ), .B(MixerOutSin_11__N_236[7]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i7_3_lut (.A(\LOSine[7] ), .B(MixerOutSin_11__N_236[6]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i3_3_lut (.A(\LOSine[3] ), .B(MixerOutSin_11__N_236[2]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i2_3_lut (.A(\LOSine[2] ), .B(MixerOutSin_11__N_236[1]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i12_3_lut (.A(\LOCosine[12] ), .B(MixerOutCos_11__N_250[11]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i11_3_lut (.A(\LOCosine[11] ), .B(MixerOutCos_11__N_250[10]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i10_3_lut (.A(\LOCosine[10] ), .B(MixerOutCos_11__N_250[9]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i9_3_lut (.A(\LOCosine[9] ), .B(MixerOutCos_11__N_250[8]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i8_3_lut (.A(\LOCosine[8] ), .B(MixerOutCos_11__N_250[7]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i7_3_lut (.A(\LOCosine[7] ), .B(MixerOutCos_11__N_250[6]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i6_3_lut (.A(\LOCosine[6] ), .B(MixerOutCos_11__N_250[5]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i5_3_lut (.A(\LOCosine[5] ), .B(MixerOutCos_11__N_250[4]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i4_3_lut (.A(\LOCosine[4] ), .B(MixerOutCos_11__N_250[3]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i3_3_lut (.A(\LOCosine[3] ), .B(MixerOutCos_11__N_250[2]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i2_3_lut (.A(\LOCosine[2] ), .B(MixerOutCos_11__N_250[1]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i12_3_lut (.A(\LOSine[12] ), .B(MixerOutSin_11__N_236[11]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i12_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module PWM
//

module PWM (\DataInReg[0] , clk_80mhz, \DataInReg_11__N_1856[0] , counter, 
            GND_net, VCC_net, \DataInReg[1] , \DataInReg_11__N_1856[1] , 
            \DataInReg[2] , \DataInReg_11__N_1856[2] , \DataInReg[3] , 
            \DataInReg_11__N_1856[3] , \DataInReg[4] , \DataInReg_11__N_1856[4] , 
            \DataInReg[5] , \DataInReg_11__N_1856[5] , \DataInReg[6] , 
            \DataInReg_11__N_1856[6] , \DataInReg[7] , \DataInReg_11__N_1856[7] , 
            \DataInReg[8] , \DataInReg_11__N_1856[8] , \DataInReg[9] , 
            \DemodOut[9] ) /* synthesis syn_module_defined=1 */ ;
    output \DataInReg[0] ;
    input clk_80mhz;
    input \DataInReg_11__N_1856[0] ;
    output [9:0]counter;
    input GND_net;
    input VCC_net;
    output \DataInReg[1] ;
    input \DataInReg_11__N_1856[1] ;
    output \DataInReg[2] ;
    input \DataInReg_11__N_1856[2] ;
    output \DataInReg[3] ;
    input \DataInReg_11__N_1856[3] ;
    output \DataInReg[4] ;
    input \DataInReg_11__N_1856[4] ;
    output \DataInReg[5] ;
    input \DataInReg_11__N_1856[5] ;
    output \DataInReg[6] ;
    input \DataInReg_11__N_1856[6] ;
    output \DataInReg[7] ;
    input \DataInReg_11__N_1856[7] ;
    output \DataInReg[8] ;
    input \DataInReg_11__N_1856[8] ;
    output \DataInReg[9] ;
    input \DemodOut[9] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(61[23:32])
    
    wire clk_80mhz_enable_1365, n16089;
    wire [9:0]n45;
    
    wire n16088, n16087, n16086, n16085;
    wire [11:0]n4027;
    
    wire n17, n15, n11, n12;
    
    FD1P3AX DataInReg__i1 (.D(\DataInReg_11__N_1856[0] ), .SP(clk_80mhz_enable_1365), 
            .CK(clk_80mhz), .Q(\DataInReg[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(41[8] 52[7])
    defparam DataInReg__i1.GSR = "ENABLED";
    CCU2C counter_955_add_4_11 (.A0(counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16089), .S0(n45[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955_add_4_11.INIT0 = 16'haaa0;
    defparam counter_955_add_4_11.INIT1 = 16'h0000;
    defparam counter_955_add_4_11.INJECT1_0 = "NO";
    defparam counter_955_add_4_11.INJECT1_1 = "NO";
    CCU2C counter_955_add_4_9 (.A0(counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16088), .COUT(n16089), .S0(n45[7]), .S1(n45[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955_add_4_9.INIT0 = 16'haaa0;
    defparam counter_955_add_4_9.INIT1 = 16'haaa0;
    defparam counter_955_add_4_9.INJECT1_0 = "NO";
    defparam counter_955_add_4_9.INJECT1_1 = "NO";
    CCU2C counter_955_add_4_7 (.A0(counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16087), .COUT(n16088), .S0(n45[5]), .S1(n45[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955_add_4_7.INIT0 = 16'haaa0;
    defparam counter_955_add_4_7.INIT1 = 16'haaa0;
    defparam counter_955_add_4_7.INJECT1_0 = "NO";
    defparam counter_955_add_4_7.INJECT1_1 = "NO";
    CCU2C counter_955_add_4_5 (.A0(counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16086), .COUT(n16087), .S0(n45[3]), .S1(n45[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955_add_4_5.INIT0 = 16'haaa0;
    defparam counter_955_add_4_5.INIT1 = 16'haaa0;
    defparam counter_955_add_4_5.INJECT1_0 = "NO";
    defparam counter_955_add_4_5.INJECT1_1 = "NO";
    CCU2C counter_955_add_4_3 (.A0(counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16085), .COUT(n16086), .S0(n45[1]), .S1(n45[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955_add_4_3.INIT0 = 16'haaa0;
    defparam counter_955_add_4_3.INIT1 = 16'haaa0;
    defparam counter_955_add_4_3.INJECT1_0 = "NO";
    defparam counter_955_add_4_3.INJECT1_1 = "NO";
    CCU2C counter_955_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16085), .S1(n45[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955_add_4_1.INIT0 = 16'h0000;
    defparam counter_955_add_4_1.INIT1 = 16'h555f;
    defparam counter_955_add_4_1.INJECT1_0 = "NO";
    defparam counter_955_add_4_1.INJECT1_1 = "NO";
    FD1S3AX counter_955__i0 (.D(n45[0]), .CK(clk_80mhz), .Q(counter[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955__i0.GSR = "ENABLED";
    FD1P3AX DataInReg__i2 (.D(\DataInReg_11__N_1856[1] ), .SP(clk_80mhz_enable_1365), 
            .CK(clk_80mhz), .Q(\DataInReg[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(41[8] 52[7])
    defparam DataInReg__i2.GSR = "ENABLED";
    FD1P3AX DataInReg__i3 (.D(\DataInReg_11__N_1856[2] ), .SP(clk_80mhz_enable_1365), 
            .CK(clk_80mhz), .Q(\DataInReg[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(41[8] 52[7])
    defparam DataInReg__i3.GSR = "ENABLED";
    FD1P3AX DataInReg__i4 (.D(\DataInReg_11__N_1856[3] ), .SP(clk_80mhz_enable_1365), 
            .CK(clk_80mhz), .Q(\DataInReg[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(41[8] 52[7])
    defparam DataInReg__i4.GSR = "ENABLED";
    FD1P3AX DataInReg__i5 (.D(\DataInReg_11__N_1856[4] ), .SP(clk_80mhz_enable_1365), 
            .CK(clk_80mhz), .Q(\DataInReg[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(41[8] 52[7])
    defparam DataInReg__i5.GSR = "ENABLED";
    FD1P3AX DataInReg__i6 (.D(\DataInReg_11__N_1856[5] ), .SP(clk_80mhz_enable_1365), 
            .CK(clk_80mhz), .Q(\DataInReg[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(41[8] 52[7])
    defparam DataInReg__i6.GSR = "ENABLED";
    FD1P3AX DataInReg__i7 (.D(\DataInReg_11__N_1856[6] ), .SP(clk_80mhz_enable_1365), 
            .CK(clk_80mhz), .Q(\DataInReg[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(41[8] 52[7])
    defparam DataInReg__i7.GSR = "ENABLED";
    FD1P3AX DataInReg__i8 (.D(\DataInReg_11__N_1856[7] ), .SP(clk_80mhz_enable_1365), 
            .CK(clk_80mhz), .Q(\DataInReg[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(41[8] 52[7])
    defparam DataInReg__i8.GSR = "ENABLED";
    FD1P3AX DataInReg__i9 (.D(\DataInReg_11__N_1856[8] ), .SP(clk_80mhz_enable_1365), 
            .CK(clk_80mhz), .Q(\DataInReg[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(41[8] 52[7])
    defparam DataInReg__i9.GSR = "ENABLED";
    FD1P3AX DataInReg__i10 (.D(n4027[9]), .SP(clk_80mhz_enable_1365), .CK(clk_80mhz), 
            .Q(\DataInReg[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(41[8] 52[7])
    defparam DataInReg__i10.GSR = "ENABLED";
    FD1S3AX counter_955__i1 (.D(n45[1]), .CK(clk_80mhz), .Q(counter[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955__i1.GSR = "ENABLED";
    FD1S3AX counter_955__i2 (.D(n45[2]), .CK(clk_80mhz), .Q(counter[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955__i2.GSR = "ENABLED";
    FD1S3AX counter_955__i3 (.D(n45[3]), .CK(clk_80mhz), .Q(counter[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955__i3.GSR = "ENABLED";
    FD1S3AX counter_955__i4 (.D(n45[4]), .CK(clk_80mhz), .Q(counter[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955__i4.GSR = "ENABLED";
    FD1S3AX counter_955__i5 (.D(n45[5]), .CK(clk_80mhz), .Q(counter[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955__i5.GSR = "ENABLED";
    FD1S3AX counter_955__i6 (.D(n45[6]), .CK(clk_80mhz), .Q(counter[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955__i6.GSR = "ENABLED";
    FD1S3AX counter_955__i7 (.D(n45[7]), .CK(clk_80mhz), .Q(counter[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955__i7.GSR = "ENABLED";
    FD1S3AX counter_955__i8 (.D(n45[8]), .CK(clk_80mhz), .Q(counter[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955__i8.GSR = "ENABLED";
    FD1S3AX counter_955__i9 (.D(n45[9]), .CK(clk_80mhz), .Q(counter[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_955__i9.GSR = "ENABLED";
    LUT4 i6034_4_lut (.A(n17), .B(n15), .C(n11), .D(n12), .Z(clk_80mhz_enable_1365)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(44[11:23])
    defparam i6034_4_lut.init = 16'h0001;
    LUT4 i7_4_lut (.A(counter[3]), .B(counter[2]), .C(counter[1]), .D(counter[9]), 
         .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(44[11:23])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(counter[6]), .B(counter[4]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(44[11:23])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(counter[0]), .B(counter[5]), .Z(n11)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(44[11:23])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2_2_lut (.A(counter[7]), .B(counter[8]), .Z(n12)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(44[11:23])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1106_1_lut (.A(\DemodOut[9] ), .Z(n4027[9])) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/PWM.v(44[7] 46[10])
    defparam i1106_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module SinCos
//

module SinCos (clk_80mhz, VCC_net, GND_net, \phase_accum[57] , \phase_accum[58] , 
            \phase_accum[59] , \phase_accum[60] , \phase_accum[61] , \phase_accum[62] , 
            \phase_accum[63] , \LOSine[1] , \LOSine[2] , \LOSine[3] , 
            \LOSine[4] , \LOSine[5] , \LOSine[6] , \LOSine[7] , \LOSine[8] , 
            \LOSine[9] , \LOSine[10] , \LOSine[11] , \LOSine[12] , \LOCosine[1] , 
            \LOCosine[2] , \LOCosine[3] , \LOCosine[4] , \LOCosine[5] , 
            \LOCosine[6] , \LOCosine[7] , \LOCosine[8] , \LOCosine[9] , 
            \LOCosine[10] , \LOCosine[11] , \LOCosine[12] , \phase_accum[56] ) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk_80mhz;
    input VCC_net;
    input GND_net;
    input \phase_accum[57] ;
    input \phase_accum[58] ;
    input \phase_accum[59] ;
    input \phase_accum[60] ;
    input \phase_accum[61] ;
    input \phase_accum[62] ;
    input \phase_accum[63] ;
    output \LOSine[1] ;
    output \LOSine[2] ;
    output \LOSine[3] ;
    output \LOSine[4] ;
    output \LOSine[5] ;
    output \LOSine[6] ;
    output \LOSine[7] ;
    output \LOSine[8] ;
    output \LOSine[9] ;
    output \LOSine[10] ;
    output \LOSine[11] ;
    output \LOSine[12] ;
    output \LOCosine[1] ;
    output \LOCosine[2] ;
    output \LOCosine[3] ;
    output \LOCosine[4] ;
    output \LOCosine[5] ;
    output \LOCosine[6] ;
    output \LOCosine[7] ;
    output \LOCosine[8] ;
    output \LOCosine[9] ;
    output \LOCosine[10] ;
    output \LOCosine[11] ;
    output \LOCosine[12] ;
    input \phase_accum[56] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(61[23:32])
    
    wire rom_addr0_r_1, rom_addr0_r_1_inv, rom_addr0_r_2, rom_addr0_r_3, 
        rom_addr0_r_4, rom_addr0_r_5, mx_ctrl_r, mx_ctrl_r_1, rom_addr0_r, 
        rom_addr0_r_n, rom_addr0_r_6, rom_dout_11, rom_dout_11_ffin, 
        rom_dout_10, rom_dout_10_ffin, rom_dout_9, rom_dout_9_ffin, 
        rom_dout_8, rom_dout_8_ffin, rom_dout_7, rom_dout_7_ffin, rom_dout_6, 
        rom_dout_6_ffin, rom_dout_5, rom_dout_5_ffin, rom_dout_4, rom_dout_4_ffin, 
        rom_dout_3, rom_dout_3_ffin, rom_dout_2, rom_dout_2_ffin, rom_dout_1, 
        rom_dout_1_ffin, rom_dout, rom_dout_ffin, rom_dout_25, rom_dout_25_ffin, 
        rom_dout_24, rom_dout_24_ffin, rom_dout_23, rom_dout_23_ffin, 
        rom_dout_22, rom_dout_22_ffin, rom_dout_21, rom_dout_21_ffin, 
        rom_dout_20, rom_dout_20_ffin, rom_dout_19, rom_dout_19_ffin, 
        rom_dout_18, rom_dout_18_ffin, rom_dout_17, rom_dout_17_ffin, 
        rom_dout_16, rom_dout_16_ffin, rom_dout_15, rom_dout_15_ffin, 
        rom_dout_14, rom_dout_14_ffin, rom_dout_13, rom_dout_13_ffin, 
        cosromoutsel_i, cosromoutsel, sinromoutsel, sinout_pre_1, sinout_pre_2, 
        sinout_pre_3, sinout_pre_4, sinout_pre_5, sinout_pre_6, sinout_pre_7, 
        sinout_pre_8, sinout_pre_9, sinout_pre_10, sinout_pre_11, sinout_pre_12, 
        cosout_pre_1, cosout_pre_2, cosout_pre_3, cosout_pre_4, cosout_pre_5, 
        cosout_pre_6, cosout_pre_7, cosout_pre_8, cosout_pre_9, cosout_pre_10, 
        cosout_pre_11, cosout_pre_12, rom_addr0_r_inv, co0, rom_addr0_r_n_1, 
        rom_addr0_r_n_2, rom_addr0_r_2_inv, co1, rom_addr0_r_n_3, rom_addr0_r_n_4, 
        rom_addr0_r_4_inv, rom_addr0_r_3_inv, co2, rom_addr0_r_n_5, 
        rom_addr0_r_5_inv, rom_dout_12_ffin, rom_addr0_r_7, rom_addr0_r_8, 
        rom_addr0_r_9, rom_addr0_r_10, rom_addr0_r_11, rom_dout_s_n_1, 
        rom_dout_s_n_2, rom_dout_2_inv, rom_dout_1_inv, co0_1, co1_1, 
        rom_dout_s_n_3, rom_dout_s_n_4, rom_dout_4_inv, rom_dout_3_inv, 
        co2_1, rom_dout_s_n_5, rom_dout_s_n_6, rom_dout_6_inv, rom_dout_5_inv, 
        co3, rom_dout_s_n_7, rom_dout_s_n_8, rom_dout_8_inv, rom_dout_7_inv, 
        co4, rom_dout_s_n_9, rom_dout_s_n_10, rom_dout_10_inv, rom_dout_9_inv, 
        co5, rom_dout_s_n_11, rom_dout_s_n_12, rom_dout_12_inv, rom_dout_11_inv, 
        rom_dout_13_inv, co0_2, rom_dout_c_n_1, rom_dout_c_n_2, rom_dout_15_inv, 
        rom_dout_14_inv, co1_2, rom_dout_c_n_3, rom_dout_c_n_4, rom_dout_17_inv, 
        rom_dout_16_inv, co2_2, rom_dout_c_n_5, rom_dout_c_n_6, rom_dout_19_inv, 
        rom_dout_18_inv, co3_1, rom_dout_c_n_7, rom_dout_c_n_8, rom_dout_21_inv, 
        rom_dout_20_inv, co4_1, rom_dout_c_n_9, rom_dout_c_n_10, rom_dout_23_inv, 
        rom_dout_22_inv, co5_1, rom_dout_c_n_11, rom_dout_c_n_12, rom_dout_25_inv, 
        rom_dout_24_inv, rom_dout_12, rom_dout_inv, func_or_inet, lx_ne0, 
        lx_ne0_inv, out_sel_i, rom_dout_s_1, rom_dout_s_2, rom_dout_s_3, 
        rom_dout_s_4, rom_dout_s_5, rom_dout_s_6, rom_dout_s_7, rom_dout_s_8, 
        rom_dout_s_9, rom_dout_s_10, rom_dout_s_11, rom_dout_s_12, rom_dout_c_1, 
        rom_dout_c_2, rom_dout_c_3, rom_dout_c_4, rom_dout_c_5, rom_dout_c_6, 
        rom_dout_c_7, rom_dout_c_8, rom_dout_c_9, rom_dout_c_10, rom_dout_c_11, 
        rom_dout_c_12, out_sel;
    
    INV INV_29 (.A(rom_addr0_r_1), .Z(rom_addr0_r_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    FD1P3DX FF_61 (.D(\phase_accum[57] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(312[13:88])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(\phase_accum[58] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(315[13:88])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(\phase_accum[59] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(318[13:88])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(\phase_accum[60] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(321[13:88])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(\phase_accum[61] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(324[13:88])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(\phase_accum[62] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(mx_ctrl_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(327[13:84])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(\phase_accum[63] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(mx_ctrl_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(330[13:86])
    defparam FF_55.GSR = "ENABLED";
    MUX21 muxb_57 (.D0(rom_addr0_r), .D1(rom_addr0_r_n), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    FD1P3DX FF_53 (.D(rom_dout_11_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(355[13] 356[25])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rom_dout_10_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(359[13] 360[25])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(rom_dout_9_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(363[13] 364[24])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(rom_dout_8_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(367[13] 368[24])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(rom_dout_7_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(371[13] 372[24])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(rom_dout_6_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(375[13] 376[24])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(rom_dout_5_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(379[13] 380[24])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(rom_dout_4_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(383[13] 384[24])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(rom_dout_3_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(387[13] 388[24])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(rom_dout_2_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(391[13] 392[24])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(rom_dout_1_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(395[13] 396[24])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(rom_dout_ffin), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(rom_dout)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(399[13] 400[22])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(rom_dout_25_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_25)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(403[13] 404[25])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(rom_dout_24_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_24)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(407[13] 408[25])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(rom_dout_23_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(411[13] 412[25])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(rom_dout_22_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(415[13] 416[25])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(rom_dout_21_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(419[13] 420[25])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(rom_dout_20_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(423[13] 424[25])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(rom_dout_19_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(427[13] 428[25])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(rom_dout_18_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(431[13] 432[25])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(rom_dout_17_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(435[13] 436[25])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(rom_dout_16_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(439[13] 440[25])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(rom_dout_15_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(443[13] 444[25])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(rom_dout_14_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(447[13] 448[25])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(rom_dout_13_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(451[13] 452[25])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(cosromoutsel_i), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(cosromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(455[13] 456[26])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(mx_ctrl_r_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(sinromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(459[13] 460[26])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(sinout_pre_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(599[13] 600[21])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(sinout_pre_2), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(603[13] 604[21])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(sinout_pre_3), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(607[13] 608[21])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(sinout_pre_4), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(611[13] 612[21])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(sinout_pre_5), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(615[13] 616[21])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(sinout_pre_6), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(619[13] 620[21])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(sinout_pre_7), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(623[13] 624[21])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(sinout_pre_8), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(627[13] 628[21])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(sinout_pre_9), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(631[13] 632[21])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(sinout_pre_10), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(635[13] 636[22])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(sinout_pre_11), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(639[13] 640[22])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(sinout_pre_12), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(643[13] 644[22])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(cosout_pre_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(650[13] 651[23])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(cosout_pre_2), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(654[13] 655[23])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(cosout_pre_3), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(658[13] 659[23])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(cosout_pre_4), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(662[13] 663[23])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(cosout_pre_5), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(666[13] 667[23])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(cosout_pre_6), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(670[13] 671[23])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(cosout_pre_7), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(674[13] 675[23])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(cosout_pre_8), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(678[13] 679[23])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(cosout_pre_9), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(682[13] 683[23])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(cosout_pre_10), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(686[13] 687[24])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(cosout_pre_11), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(690[13] 691[24])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(cosout_pre_12), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(694[13] 695[24])
    defparam FF_0.GSR = "ENABLED";
    CCU2C neg_rom_addr0_r_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0), .S1(rom_addr0_r_n)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(702[11] 704[71])
    defparam neg_rom_addr0_r_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_0.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_0.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_1 (.A0(rom_addr0_r_1_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_2_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0), .COUT(co1), .S0(rom_addr0_r_n_1), 
          .S1(rom_addr0_r_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(710[11] 713[42])
    defparam neg_rom_addr0_r_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_1.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_2 (.A0(rom_addr0_r_3_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_4_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1), .COUT(co2), .S0(rom_addr0_r_n_3), 
          .S1(rom_addr0_r_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(719[11] 722[42])
    defparam neg_rom_addr0_r_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_2.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_3 (.A0(rom_addr0_r_5_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co2), .S0(rom_addr0_r_n_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(728[11] 730[73])
    defparam neg_rom_addr0_r_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_3.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_3.INJECT1_1 = "NO";
    ROM64X1A triglut_1_0_25 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_12_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_25.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    CCU2C neg_rom_dout_s_n_1 (.A0(rom_dout_1_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_2_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0_1), .COUT(co1_1), .S0(rom_dout_s_n_1), 
          .S1(rom_dout_s_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(874[11] 877[43])
    defparam neg_rom_dout_s_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_1.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_2 (.A0(rom_dout_3_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_4_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1_1), .COUT(co2_1), .S0(rom_dout_s_n_3), 
          .S1(rom_dout_s_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(883[11] 886[43])
    defparam neg_rom_dout_s_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_2.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_3 (.A0(rom_dout_5_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_6_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co2_1), .COUT(co3), .S0(rom_dout_s_n_5), 
          .S1(rom_dout_s_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(892[11] 895[41])
    defparam neg_rom_dout_s_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_3.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_3.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_4 (.A0(rom_dout_7_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_8_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co3), .COUT(co4), .S0(rom_dout_s_n_7), 
          .S1(rom_dout_s_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(901[11] 904[41])
    defparam neg_rom_dout_s_n_4.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_4.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_4.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_4.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_5 (.A0(rom_dout_9_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_10_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co4), .COUT(co5), .S0(rom_dout_s_n_9), 
          .S1(rom_dout_s_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(910[11] 913[42])
    defparam neg_rom_dout_s_n_5.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_5.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_5.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_5.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_6 (.A0(rom_dout_11_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_12_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co5), .S0(rom_dout_s_n_11), .S1(rom_dout_s_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(919[11] 922[42])
    defparam neg_rom_dout_s_n_6.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_6.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_6.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_6.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_13_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(936[11] 938[72])
    defparam neg_rom_dout_c_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_0.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_0.INJECT1_1 = "NO";
    INV INV_30 (.A(rom_addr0_r_2), .Z(rom_addr0_r_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    CCU2C neg_rom_dout_c_n_1 (.A0(rom_dout_14_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_15_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0_2), .COUT(co1_2), .S0(rom_dout_c_n_1), 
          .S1(rom_dout_c_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(944[11] 947[43])
    defparam neg_rom_dout_c_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_1.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_2 (.A0(rom_dout_16_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_17_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1_2), .COUT(co2_2), .S0(rom_dout_c_n_3), 
          .S1(rom_dout_c_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(953[11] 956[43])
    defparam neg_rom_dout_c_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_2.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_3 (.A0(rom_dout_18_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_19_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co2_2), .COUT(co3_1), .S0(rom_dout_c_n_5), 
          .S1(rom_dout_c_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(962[11] 965[43])
    defparam neg_rom_dout_c_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_3.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_3.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_4 (.A0(rom_dout_20_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_21_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co3_1), .COUT(co4_1), .S0(rom_dout_c_n_7), 
          .S1(rom_dout_c_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(971[11] 974[43])
    defparam neg_rom_dout_c_n_4.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_4.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_4.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_4.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_5 (.A0(rom_dout_22_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_23_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co4_1), .COUT(co5_1), .S0(rom_dout_c_n_9), 
          .S1(rom_dout_c_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(980[11] 983[44])
    defparam neg_rom_dout_c_n_5.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_5.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_5.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_5.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_6 (.A0(rom_dout_24_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_25_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co5_1), .S0(rom_dout_c_n_11), .S1(rom_dout_c_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(989[11] 992[44])
    defparam neg_rom_dout_c_n_6.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_6.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_6.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_6.INJECT1_1 = "NO";
    INV INV_31 (.A(rom_addr0_r_3), .Z(rom_addr0_r_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_32 (.A(rom_addr0_r_4), .Z(rom_addr0_r_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_33 (.A(rom_addr0_r_5), .Z(rom_addr0_r_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_28 (.A(rom_addr0_r), .Z(rom_addr0_r_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    XOR2 XOR2_t1 (.A(mx_ctrl_r), .B(mx_ctrl_r_1), .Z(cosromoutsel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(241[10:70])
    INV INV_27 (.A(rom_dout_12), .Z(rom_dout_12_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_26 (.A(rom_dout_11), .Z(rom_dout_11_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_25 (.A(rom_dout_10), .Z(rom_dout_10_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_24 (.A(rom_dout_9), .Z(rom_dout_9_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_23 (.A(rom_dout_8), .Z(rom_dout_8_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_22 (.A(rom_dout_7), .Z(rom_dout_7_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_21 (.A(rom_dout_6), .Z(rom_dout_6_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_20 (.A(rom_dout_5), .Z(rom_dout_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_19 (.A(rom_dout_4), .Z(rom_dout_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_18 (.A(rom_dout_3), .Z(rom_dout_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_17 (.A(rom_dout_2), .Z(rom_dout_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_16 (.A(rom_dout_1), .Z(rom_dout_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_15 (.A(rom_dout), .Z(rom_dout_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_14 (.A(rom_dout_25), .Z(rom_dout_25_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_13 (.A(rom_dout_24), .Z(rom_dout_24_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_12 (.A(rom_dout_23), .Z(rom_dout_23_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_11 (.A(rom_dout_22), .Z(rom_dout_22_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_10 (.A(rom_dout_21), .Z(rom_dout_21_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_9 (.A(rom_dout_20), .Z(rom_dout_20_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_8 (.A(rom_dout_19), .Z(rom_dout_19_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_7 (.A(rom_dout_18), .Z(rom_dout_18_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_6 (.A(rom_dout_17), .Z(rom_dout_17_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_5 (.A(rom_dout_16), .Z(rom_dout_16_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_4 (.A(rom_dout_15), .Z(rom_dout_15_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_3 (.A(rom_dout_14), .Z(rom_dout_14_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_2 (.A(rom_dout_13), .Z(rom_dout_13_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    ROM16X1A LUT4_1 (.AD0(rom_addr0_r_9), .AD1(rom_addr0_r_8), .AD2(rom_addr0_r_7), 
            .AD3(rom_addr0_r_6), .DO0(func_or_inet)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam LUT4_1.initval = 16'b1111111111111110;
    ROM16X1A LUT4_0 (.AD0(GND_net), .AD1(rom_addr0_r_11), .AD2(rom_addr0_r_10), 
            .AD3(func_or_inet), .DO0(lx_ne0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam LUT4_0.initval = 16'b1111111111111110;
    INV INV_1 (.A(lx_ne0), .Z(lx_ne0_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    AND2 AND2_t0 (.A(mx_ctrl_r), .B(lx_ne0_inv), .Z(out_sel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(305[10:64])
    FD1P3DX FF_62 (.D(\phase_accum[56] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(309[13:86])
    defparam FF_62.GSR = "ENABLED";
    MUX21 muxb_56 (.D0(rom_addr0_r_1), .D1(rom_addr0_r_n_1), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_55 (.D0(rom_addr0_r_2), .D1(rom_addr0_r_n_2), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_54 (.D0(rom_addr0_r_3), .D1(rom_addr0_r_n_3), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_53 (.D0(rom_addr0_r_4), .D1(rom_addr0_r_n_4), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_52 (.D0(rom_addr0_r_5), .D1(rom_addr0_r_n_5), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    FD1P3DX FF_54 (.D(rom_dout_12_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(351[13] 352[25])
    defparam FF_54.GSR = "ENABLED";
    MUX21 muxb_50 (.D0(rom_dout_1), .D1(rom_dout_s_n_1), .SD(sinromoutsel), 
          .Z(rom_dout_s_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_49 (.D0(rom_dout_2), .D1(rom_dout_s_n_2), .SD(sinromoutsel), 
          .Z(rom_dout_s_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_48 (.D0(rom_dout_3), .D1(rom_dout_s_n_3), .SD(sinromoutsel), 
          .Z(rom_dout_s_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_47 (.D0(rom_dout_4), .D1(rom_dout_s_n_4), .SD(sinromoutsel), 
          .Z(rom_dout_s_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_46 (.D0(rom_dout_5), .D1(rom_dout_s_n_5), .SD(sinromoutsel), 
          .Z(rom_dout_s_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_45 (.D0(rom_dout_6), .D1(rom_dout_s_n_6), .SD(sinromoutsel), 
          .Z(rom_dout_s_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_44 (.D0(rom_dout_7), .D1(rom_dout_s_n_7), .SD(sinromoutsel), 
          .Z(rom_dout_s_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_43 (.D0(rom_dout_8), .D1(rom_dout_s_n_8), .SD(sinromoutsel), 
          .Z(rom_dout_s_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_42 (.D0(rom_dout_9), .D1(rom_dout_s_n_9), .SD(sinromoutsel), 
          .Z(rom_dout_s_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_41 (.D0(rom_dout_10), .D1(rom_dout_s_n_10), .SD(sinromoutsel), 
          .Z(rom_dout_s_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_40 (.D0(rom_dout_11), .D1(rom_dout_s_n_11), .SD(sinromoutsel), 
          .Z(rom_dout_s_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_39 (.D0(rom_dout_12), .D1(rom_dout_s_n_12), .SD(sinromoutsel), 
          .Z(rom_dout_s_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_37 (.D0(rom_dout_14), .D1(rom_dout_c_n_1), .SD(cosromoutsel), 
          .Z(rom_dout_c_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_36 (.D0(rom_dout_15), .D1(rom_dout_c_n_2), .SD(cosromoutsel), 
          .Z(rom_dout_c_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_35 (.D0(rom_dout_16), .D1(rom_dout_c_n_3), .SD(cosromoutsel), 
          .Z(rom_dout_c_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_34 (.D0(rom_dout_17), .D1(rom_dout_c_n_4), .SD(cosromoutsel), 
          .Z(rom_dout_c_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_33 (.D0(rom_dout_18), .D1(rom_dout_c_n_5), .SD(cosromoutsel), 
          .Z(rom_dout_c_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_32 (.D0(rom_dout_19), .D1(rom_dout_c_n_6), .SD(cosromoutsel), 
          .Z(rom_dout_c_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_31 (.D0(rom_dout_20), .D1(rom_dout_c_n_7), .SD(cosromoutsel), 
          .Z(rom_dout_c_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_30 (.D0(rom_dout_21), .D1(rom_dout_c_n_8), .SD(cosromoutsel), 
          .Z(rom_dout_c_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_29 (.D0(rom_dout_22), .D1(rom_dout_c_n_9), .SD(cosromoutsel), 
          .Z(rom_dout_c_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_28 (.D0(rom_dout_23), .D1(rom_dout_c_n_10), .SD(cosromoutsel), 
          .Z(rom_dout_c_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_27 (.D0(rom_dout_24), .D1(rom_dout_c_n_11), .SD(cosromoutsel), 
          .Z(rom_dout_c_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_26 (.D0(rom_dout_25), .D1(rom_dout_c_n_12), .SD(cosromoutsel), 
          .Z(rom_dout_c_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    FD1P3DX FF_26 (.D(out_sel_i), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(out_sel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(541[13:83])
    defparam FF_26.GSR = "ENABLED";
    MUX21 muxb_24 (.D0(rom_dout_s_1), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_23 (.D0(rom_dout_s_2), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_22 (.D0(rom_dout_s_3), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_21 (.D0(rom_dout_s_4), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_20 (.D0(rom_dout_s_5), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_19 (.D0(rom_dout_s_6), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_18 (.D0(rom_dout_s_7), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_17 (.D0(rom_dout_s_8), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_16 (.D0(rom_dout_s_9), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_15 (.D0(rom_dout_s_10), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_14 (.D0(rom_dout_s_11), .D1(VCC_net), .SD(out_sel), .Z(sinout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_13 (.D0(rom_dout_s_12), .D1(mx_ctrl_r_1), .SD(out_sel), 
          .Z(sinout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_11 (.D0(rom_dout_c_1), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_10 (.D0(rom_dout_c_2), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_9 (.D0(rom_dout_c_3), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_8 (.D0(rom_dout_c_4), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_7 (.D0(rom_dout_c_5), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_6 (.D0(rom_dout_c_6), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_5 (.D0(rom_dout_c_7), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_4 (.D0(rom_dout_c_8), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_3 (.D0(rom_dout_c_9), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_2 (.D0(rom_dout_c_10), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_1 (.D0(rom_dout_c_11), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_0 (.D0(rom_dout_c_12), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    ROM64X1A triglut_1_0_24 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_11_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_24.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_23 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_10_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_23.initval = 64'b1111111111111111111111111111111111111111110000000000000000000000;
    ROM64X1A triglut_1_0_22 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_9_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_22.initval = 64'b1111111111111111111111111111100000000000001111111111100000000000;
    ROM64X1A triglut_1_0_21 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_8_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_21.initval = 64'b1111111111111111111100000000011111110000001111110000011111000000;
    ROM64X1A triglut_1_0_20 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_7_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_20.initval = 64'b1111111111111100000011111000011110001110001110001110011100111000;
    ROM64X1A triglut_1_0_19 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_6_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_19.initval = 64'b1111111111000011100011100110011001001101101101001001011010110100;
    ROM64X1A triglut_1_0_18 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_5_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_18.initval = 64'b1111111000110011011010010101010100101001001001101100110001100110;
    ROM64X1A triglut_1_0_17 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_4_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_17.initval = 64'b1111100100101010110011000000000001110011011010110101010110101010;
    ROM64X1A triglut_1_0_16 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_3_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_16.initval = 64'b1110010110011100010101001111111101101010110011100000000011110000;
    ROM64X1A triglut_1_0_15 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_2_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_15.initval = 64'b1101000010100011001111010111110011001100010101100000000011001100;
    ROM64X1A triglut_1_0_14 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_1_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_14.initval = 64'b1111011011100010010110111011101001110011000000100111110010101010;
    ROM64X1A triglut_1_0_13 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_13.initval = 64'b1000100101001010011001010111111001010010011110001001001001111000;
    ROM64X1A triglut_1_0_12 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_25_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_12.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_11 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_24_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_11.initval = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    ROM64X1A triglut_1_0_10 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_23_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_10.initval = 64'b0000000000000000000001111111111111111111111111111111111111111110;
    ROM64X1A triglut_1_0_9 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_22_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_9.initval = 64'b0000000000111111111110000000000000111111111111111111111111111110;
    ROM64X1A triglut_1_0_8 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_21_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_8.initval = 64'b0000011111000001111110000001111111000000000111111111111111111110;
    ROM64X1A triglut_1_0_7 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_20_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_7.initval = 64'b0011100111001110001110001110001111000011111000000111111111111110;
    ROM64X1A triglut_1_0_6 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_19_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_6.initval = 64'b0101101011010010010110110110010011001100111000111000011111111110;
    ROM64X1A triglut_1_0_5 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_18_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_5.initval = 64'b1100110001100110110010010010100101010101001011011001100011111110;
    ROM64X1A triglut_1_0_4 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_17_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_4.initval = 64'b1010101101010101101011011001110000000000011001101010100100111110;
    ROM64X1A triglut_1_0_3 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_16_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_3.initval = 64'b0001111000000000111001101010110111111110010101000111001101001110;
    ROM64X1A triglut_1_0_2 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_15_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_2.initval = 64'b0110011000000000110101000110011001111101011110011000101000010110;
    ROM64X1A triglut_1_0_1 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_14_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_1.initval = 64'b1010101001111100100000011001110010111011101101001000111011011110;
    ROM64X1A triglut_1_0_0 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_13_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_0.initval = 64'b0011110010010010001111001001010011111101010011001010010100100010;
    CCU2C neg_rom_dout_s_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/IP/SinCos/SinCos.v(866[11] 868[72])
    defparam neg_rom_dout_s_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_0.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_0.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PLL
//

module PLL (clk_25mhz_c, clk_80mhz, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk_25mhz_c;
    output clk_80mhz;
    input GND_net;
    
    wire clk_25mhz_c /* synthesis is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(40[22:31])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(61[23:32])
    
    EHXPLLL PLLInst_0 (.CLKI(clk_25mhz_c), .CLKFB(clk_80mhz), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .PHASELOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .CLKOP(clk_80mhz)) /* synthesis FREQUENCY_PIN_CLKOP="83.333333", FREQUENCY_PIN_CLKI="25.000000", ICP_CURRENT="5", LPF_RESISTOR="16", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=97, LSE_RLINE=100 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(97[8] 100[5])
    defparam PLLInst_0.CLKI_DIV = 3;
    defparam PLLInst_0.CLKFB_DIV = 10;
    defparam PLLInst_0.CLKOP_DIV = 7;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 6;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.CLKOP_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.PLL_LOCK_DELAY = 200;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.REFIN_RESET = "DISABLED";
    defparam PLLInst_0.SYNC_ENABLE = "DISABLED";
    defparam PLLInst_0.INT_LOCK_STICKY = "ENABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module nco_sig
//

module nco_sig (\phase_accum[63] , sinGen_c) /* synthesis syn_module_defined=1 */ ;
    input \phase_accum[63] ;
    output sinGen_c;
    
    
    LUT4 phase_accum_63__I_0_13_1_lut (.A(\phase_accum[63] ), .Z(sinGen_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/NCO.v(34[22:66])
    defparam phase_accum_63__I_0_13_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module \CIC(WIDTH=72,DECIMATION_RATIO=4096) 
//

module \CIC(WIDTH=72,DECIMATION_RATIO=4096)  (d_tmp, clk_80mhz, d5, d_d_tmp, 
            d2, d2_71__N_490, d3, d3_71__N_562, d4, d4_71__N_634, 
            d5_71__N_706, d6, d6_71__N_1459, d_d6, d7, d7_71__N_1531, 
            d_d7, d8, d8_71__N_1603, d_d8, d9, d9_71__N_1675, d_d9, 
            CIC1_outCos, d1, d1_71__N_418, count, n87_adj_228, n23, 
            n10, n35, n10_adj_115, n22, n13, n12, n15, n34, 
            n37, n14, n17, n36_adj_116, n16, n3, n2, n5, n4, 
            n7, n6, n9, n8, \CICGain[1] , \d10[60] , \d10[59] , 
            \d10[61] , \d10[62] , \d10[63] , \d10[64] , \d10[65] , 
            \d10[66] , \d10[67] , \d10[68] , \d10[69] , \d10[70] , 
            \d10[71] , \d_out_11__N_1819[2] , \d_out_11__N_1819[3] , \d_out_11__N_1819[4] , 
            \d_out_11__N_1819[5] , \d_out_11__N_1819[6] , \d_out_11__N_1819[7] , 
            \d_out_11__N_1819[8] , \d_out_11__N_1819[9] , \d_out_11__N_1819[10] , 
            \d_out_11__N_1819[11] , n11, n17325, n10_adj_117, n13_adj_118, 
            n12_adj_119, n15_adj_120, n14_adj_121, n17_adj_122, n16_adj_123, 
            n19, n18, n21, n20, n23_adj_124, n22_adj_125, n25, 
            n24, n27, n26, n31, n30, n29, n28, n17302, n33, 
            n31_adj_126, n32, n30_adj_127, n33_adj_128, n19_adj_129, 
            n32_adj_130, n35_adj_131, n35_adj_132, n34_adj_133, n18_adj_134, 
            n34_adj_135, n37_adj_136, n36_adj_137, n3_adj_138, n2_adj_139, 
            n5_adj_140, n37_adj_141, n36_adj_142, n4_adj_143, n7_adj_144, 
            n6_adj_145, n9_adj_146, n8_adj_147, n11_adj_148, n10_adj_149, 
            n13_adj_150, n12_adj_151, n15_adj_152, n14_adj_153, n17_adj_154, 
            n16_adj_155, n19_adj_156, n18_adj_157, n21_adj_158, n20_adj_159, 
            n23_adj_160, n22_adj_161, n25_adj_162, n24_adj_163, n27_adj_164, 
            n26_adj_165, n29_adj_166, n28_adj_167, n31_adj_168, n30_adj_169, 
            n33_adj_170, n5_adj_171, n4_adj_172, n7_adj_173, n6_adj_174, 
            n3_adj_175, n2_adj_176, n3_adj_177, n2_adj_178, n13_adj_179, 
            n12_adj_180, n15_adj_181, n14_adj_182, n32_adj_183, n35_adj_184, 
            n34_adj_185, n118, n120, cout, n115, n117, n112, n114, 
            n109, n111, n106, n108, n17_adj_186, n103, n105, n100, 
            n102, n97, n99, n94, n96, n5_adj_187, n91, n93, 
            n16_adj_188, n19_adj_189, n18_adj_190, n88, n90, n21_adj_191, 
            n20_adj_192, n23_adj_193, n22_adj_194, n25_adj_195, n24_adj_196, 
            n27_adj_197, n26_adj_198, n25_adj_199, n4_adj_200, n7_adj_201, 
            n29_adj_202, n21_adj_203, n28_adj_204, \CICGain[0] , n85, 
            n87, n82, n84, n20_adj_205, n31_adj_206, n6_adj_207, 
            n30_adj_208, n27_adj_209, n26_adj_210, n29_adj_211, n28_adj_212, 
            n79, n81_adj_213, n9_adj_214, n9_adj_215, n8_adj_216, 
            n76, n78_adj_217, n32_adj_218, n33_adj_219, n63_adj_220, 
            n11_adj_221, n17288, n65, n8_adj_222, n66_adj_223, n11_adj_224, 
            n37_adj_225, n36_adj_226, n24_adj_227) /* synthesis syn_module_defined=1 */ ;
    output [71:0]d_tmp;
    input clk_80mhz;
    output [71:0]d5;
    output [71:0]d_d_tmp;
    output [71:0]d2;
    input [71:0]d2_71__N_490;
    output [71:0]d3;
    input [71:0]d3_71__N_562;
    output [71:0]d4;
    input [71:0]d4_71__N_634;
    input [71:0]d5_71__N_706;
    output [71:0]d6;
    input [71:0]d6_71__N_1459;
    output [71:0]d_d6;
    output [71:0]d7;
    input [71:0]d7_71__N_1531;
    output [71:0]d_d7;
    output [71:0]d8;
    input [71:0]d8_71__N_1603;
    output [71:0]d_d8;
    output [71:0]d9;
    input [71:0]d9_71__N_1675;
    output [71:0]d_d9;
    output [11:0]CIC1_outCos;
    output [71:0]d1;
    input [71:0]d1_71__N_418;
    output [15:0]count;
    input [15:0]n87_adj_228;
    output n23;
    output n10;
    output n35;
    output n10_adj_115;
    output n22;
    output n13;
    output n12;
    output n15;
    output n34;
    output n37;
    output n14;
    output n17;
    output n36_adj_116;
    output n16;
    output n3;
    output n2;
    output n5;
    output n4;
    output n7;
    output n6;
    output n9;
    output n8;
    input \CICGain[1] ;
    output \d10[60] ;
    output \d10[59] ;
    output \d10[61] ;
    output \d10[62] ;
    output \d10[63] ;
    output \d10[64] ;
    output \d10[65] ;
    output \d10[66] ;
    output \d10[67] ;
    output \d10[68] ;
    output \d10[69] ;
    output \d10[70] ;
    output \d10[71] ;
    input \d_out_11__N_1819[2] ;
    input \d_out_11__N_1819[3] ;
    input \d_out_11__N_1819[4] ;
    input \d_out_11__N_1819[5] ;
    input \d_out_11__N_1819[6] ;
    input \d_out_11__N_1819[7] ;
    input \d_out_11__N_1819[8] ;
    input \d_out_11__N_1819[9] ;
    input \d_out_11__N_1819[10] ;
    input \d_out_11__N_1819[11] ;
    output n11;
    output n17325;
    output n10_adj_117;
    output n13_adj_118;
    output n12_adj_119;
    output n15_adj_120;
    output n14_adj_121;
    output n17_adj_122;
    output n16_adj_123;
    output n19;
    output n18;
    output n21;
    output n20;
    output n23_adj_124;
    output n22_adj_125;
    output n25;
    output n24;
    output n27;
    output n26;
    output n31;
    output n30;
    output n29;
    output n28;
    output n17302;
    output n33;
    output n31_adj_126;
    output n32;
    output n30_adj_127;
    output n33_adj_128;
    output n19_adj_129;
    output n32_adj_130;
    output n35_adj_131;
    output n35_adj_132;
    output n34_adj_133;
    output n18_adj_134;
    output n34_adj_135;
    output n37_adj_136;
    output n36_adj_137;
    output n3_adj_138;
    output n2_adj_139;
    output n5_adj_140;
    output n37_adj_141;
    output n36_adj_142;
    output n4_adj_143;
    output n7_adj_144;
    output n6_adj_145;
    output n9_adj_146;
    output n8_adj_147;
    output n11_adj_148;
    output n10_adj_149;
    output n13_adj_150;
    output n12_adj_151;
    output n15_adj_152;
    output n14_adj_153;
    output n17_adj_154;
    output n16_adj_155;
    output n19_adj_156;
    output n18_adj_157;
    output n21_adj_158;
    output n20_adj_159;
    output n23_adj_160;
    output n22_adj_161;
    output n25_adj_162;
    output n24_adj_163;
    output n27_adj_164;
    output n26_adj_165;
    output n29_adj_166;
    output n28_adj_167;
    output n31_adj_168;
    output n30_adj_169;
    output n33_adj_170;
    output n5_adj_171;
    output n4_adj_172;
    output n7_adj_173;
    output n6_adj_174;
    output n3_adj_175;
    output n2_adj_176;
    output n3_adj_177;
    output n2_adj_178;
    output n13_adj_179;
    output n12_adj_180;
    output n15_adj_181;
    output n14_adj_182;
    output n32_adj_183;
    output n35_adj_184;
    output n34_adj_185;
    input n118;
    input n120;
    input cout;
    input n115;
    input n117;
    input n112;
    input n114;
    input n109;
    input n111;
    input n106;
    input n108;
    output n17_adj_186;
    input n103;
    input n105;
    input n100;
    input n102;
    input n97;
    input n99;
    input n94;
    input n96;
    output n5_adj_187;
    input n91;
    input n93;
    output n16_adj_188;
    output n19_adj_189;
    output n18_adj_190;
    input n88;
    input n90;
    output n21_adj_191;
    output n20_adj_192;
    output n23_adj_193;
    output n22_adj_194;
    output n25_adj_195;
    output n24_adj_196;
    output n27_adj_197;
    output n26_adj_198;
    output n25_adj_199;
    output n4_adj_200;
    output n7_adj_201;
    output n29_adj_202;
    output n21_adj_203;
    output n28_adj_204;
    input \CICGain[0] ;
    input n85;
    input n87;
    input n82;
    input n84;
    output n20_adj_205;
    output n31_adj_206;
    output n6_adj_207;
    output n30_adj_208;
    output n27_adj_209;
    output n26_adj_210;
    output n29_adj_211;
    output n28_adj_212;
    input n79;
    input n81_adj_213;
    output n9_adj_214;
    output n9_adj_215;
    output n8_adj_216;
    input n76;
    input n78_adj_217;
    output n32_adj_218;
    output n33_adj_219;
    output n63_adj_220;
    output n11_adj_221;
    output n17288;
    output n65;
    output n8_adj_222;
    output n66_adj_223;
    output n11_adj_224;
    output n37_adj_225;
    output n36_adj_226;
    output n24_adj_227;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(61[23:32])
    
    wire count_15__N_1458, clk_80mhz_enable_756, v_comb;
    wire [71:0]d_out_11__N_1819;
    
    wire n12783;
    wire [15:0]count_15__N_1442;
    wire [71:0]d10;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[68:71])
    
    wire n17858, clk_80mhz_enable_806, clk_80mhz_enable_856, clk_80mhz_enable_906, 
        clk_80mhz_enable_956, clk_80mhz_enable_1006, clk_80mhz_enable_1056, 
        clk_80mhz_enable_1106, clk_80mhz_enable_1156, clk_80mhz_enable_1206, 
        clk_80mhz_enable_1256, clk_80mhz_enable_1306, clk_80mhz_enable_1356;
    wire [71:0]d10_71__N_1747;
    
    wire n17857, n17191, n16826, n17876, n17875, n17193, n17268, 
        n17225, n17262, n17219, n17189, n17181, n17185;
    
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    FD1S3AX d2_i0 (.D(d2_71__N_490[0]), .CK(clk_80mhz), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i0.GSR = "ENABLED";
    FD1S3AX d3_i0 (.D(d3_71__N_562[0]), .CK(clk_80mhz), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_634[0]), .CK(clk_80mhz), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_706[0]), .CK(clk_80mhz), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1459[0]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1531[0]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1603[0]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1675[0]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1819[0]), .SP(clk_80mhz_enable_756), 
            .CK(clk_80mhz), .Q(CIC1_outCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_418[0]), .CK(clk_80mhz), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i0.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(n87_adj_228[1]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i1.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_15__N_1442[0]), .CK(clk_80mhz), .CD(count_15__N_1458), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i0.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i51_1_lut (.A(d_d6[50]), .Z(n23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i64_1_lut (.A(d_d7[63]), .Z(n10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i39_1_lut (.A(d_d7[38]), .Z(n35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i64_1_lut (.A(d_d6[63]), .Z(n10_adj_115)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i52_1_lut (.A(d_d6[51]), .Z(n22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i61_1_lut (.A(d_d6[60]), .Z(n13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i62_1_lut (.A(d_d6[61]), .Z(n12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i59_1_lut (.A(d_d6[58]), .Z(n15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i40_1_lut (.A(d_d7[39]), .Z(n34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i37_1_lut (.A(d_d7[36]), .Z(n37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i60_1_lut (.A(d_d6[59]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i57_1_lut (.A(d_d6[56]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i38_1_lut (.A(d_d7[37]), .Z(n36_adj_116)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i58_1_lut (.A(d_d6[57]), .Z(n16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i71_1_lut (.A(d_d8[70]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i72_1_lut (.A(d_d8[71]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i69_1_lut (.A(d_d8[68]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i70_1_lut (.A(d_d8[69]), .Z(n4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i67_1_lut (.A(d_d8[66]), .Z(n7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i68_1_lut (.A(d_d8[67]), .Z(n6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i65_1_lut (.A(d_d8[64]), .Z(n9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i66_1_lut (.A(d_d8[65]), .Z(n8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 i6080_then_3_lut (.A(\CICGain[1] ), .B(\d10[60] ), .C(d10[58]), 
         .Z(n17858)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6080_then_3_lut.init = 16'he4e4;
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(clk_80mhz_enable_756), .CK(clk_80mhz), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1S3AX d2_i1 (.D(d2_71__N_490[1]), .CK(clk_80mhz), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i1.GSR = "ENABLED";
    FD1S3AX d2_i2 (.D(d2_71__N_490[2]), .CK(clk_80mhz), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_490[3]), .CK(clk_80mhz), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_490[4]), .CK(clk_80mhz), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_490[5]), .CK(clk_80mhz), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_490[6]), .CK(clk_80mhz), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_490[7]), .CK(clk_80mhz), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_490[8]), .CK(clk_80mhz), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_490[9]), .CK(clk_80mhz), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_490[10]), .CK(clk_80mhz), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_490[11]), .CK(clk_80mhz), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_490[12]), .CK(clk_80mhz), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_490[13]), .CK(clk_80mhz), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_490[14]), .CK(clk_80mhz), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_490[15]), .CK(clk_80mhz), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_490[16]), .CK(clk_80mhz), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_490[17]), .CK(clk_80mhz), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_490[18]), .CK(clk_80mhz), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_490[19]), .CK(clk_80mhz), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_490[20]), .CK(clk_80mhz), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_490[21]), .CK(clk_80mhz), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_490[22]), .CK(clk_80mhz), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_490[23]), .CK(clk_80mhz), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_490[24]), .CK(clk_80mhz), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_490[25]), .CK(clk_80mhz), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_490[26]), .CK(clk_80mhz), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_490[27]), .CK(clk_80mhz), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_490[28]), .CK(clk_80mhz), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_490[29]), .CK(clk_80mhz), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_490[30]), .CK(clk_80mhz), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_490[31]), .CK(clk_80mhz), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_490[32]), .CK(clk_80mhz), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_490[33]), .CK(clk_80mhz), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_490[34]), .CK(clk_80mhz), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_490[35]), .CK(clk_80mhz), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_490[36]), .CK(clk_80mhz), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_490[37]), .CK(clk_80mhz), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_490[38]), .CK(clk_80mhz), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_490[39]), .CK(clk_80mhz), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_490[40]), .CK(clk_80mhz), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_490[41]), .CK(clk_80mhz), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_490[42]), .CK(clk_80mhz), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_490[43]), .CK(clk_80mhz), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_490[44]), .CK(clk_80mhz), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_490[45]), .CK(clk_80mhz), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_490[46]), .CK(clk_80mhz), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_490[47]), .CK(clk_80mhz), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_490[48]), .CK(clk_80mhz), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_490[49]), .CK(clk_80mhz), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_490[50]), .CK(clk_80mhz), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_490[51]), .CK(clk_80mhz), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_490[52]), .CK(clk_80mhz), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_490[53]), .CK(clk_80mhz), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_490[54]), .CK(clk_80mhz), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_490[55]), .CK(clk_80mhz), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_490[56]), .CK(clk_80mhz), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_490[57]), .CK(clk_80mhz), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_490[58]), .CK(clk_80mhz), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_490[59]), .CK(clk_80mhz), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_490[60]), .CK(clk_80mhz), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_490[61]), .CK(clk_80mhz), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_490[62]), .CK(clk_80mhz), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_490[63]), .CK(clk_80mhz), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_490[64]), .CK(clk_80mhz), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_490[65]), .CK(clk_80mhz), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_490[66]), .CK(clk_80mhz), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_490[67]), .CK(clk_80mhz), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_490[68]), .CK(clk_80mhz), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_490[69]), .CK(clk_80mhz), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_490[70]), .CK(clk_80mhz), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_490[71]), .CK(clk_80mhz), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_562[1]), .CK(clk_80mhz), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_562[2]), .CK(clk_80mhz), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_562[3]), .CK(clk_80mhz), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_562[4]), .CK(clk_80mhz), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_562[5]), .CK(clk_80mhz), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_562[6]), .CK(clk_80mhz), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_562[7]), .CK(clk_80mhz), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_562[8]), .CK(clk_80mhz), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_562[9]), .CK(clk_80mhz), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_562[10]), .CK(clk_80mhz), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_562[11]), .CK(clk_80mhz), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_562[12]), .CK(clk_80mhz), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_562[13]), .CK(clk_80mhz), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_562[14]), .CK(clk_80mhz), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_562[15]), .CK(clk_80mhz), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_562[16]), .CK(clk_80mhz), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_562[17]), .CK(clk_80mhz), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_562[18]), .CK(clk_80mhz), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_562[19]), .CK(clk_80mhz), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_562[20]), .CK(clk_80mhz), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_562[21]), .CK(clk_80mhz), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_562[22]), .CK(clk_80mhz), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_562[23]), .CK(clk_80mhz), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_562[24]), .CK(clk_80mhz), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_562[25]), .CK(clk_80mhz), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_562[26]), .CK(clk_80mhz), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_562[27]), .CK(clk_80mhz), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_562[28]), .CK(clk_80mhz), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_562[29]), .CK(clk_80mhz), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_562[30]), .CK(clk_80mhz), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_562[31]), .CK(clk_80mhz), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_562[32]), .CK(clk_80mhz), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_562[33]), .CK(clk_80mhz), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_562[34]), .CK(clk_80mhz), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_562[35]), .CK(clk_80mhz), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_562[36]), .CK(clk_80mhz), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_562[37]), .CK(clk_80mhz), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_562[38]), .CK(clk_80mhz), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_562[39]), .CK(clk_80mhz), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_562[40]), .CK(clk_80mhz), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_562[41]), .CK(clk_80mhz), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_562[42]), .CK(clk_80mhz), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_562[43]), .CK(clk_80mhz), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_562[44]), .CK(clk_80mhz), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_562[45]), .CK(clk_80mhz), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_562[46]), .CK(clk_80mhz), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_562[47]), .CK(clk_80mhz), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_562[48]), .CK(clk_80mhz), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_562[49]), .CK(clk_80mhz), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_562[50]), .CK(clk_80mhz), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_562[51]), .CK(clk_80mhz), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_562[52]), .CK(clk_80mhz), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_562[53]), .CK(clk_80mhz), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_562[54]), .CK(clk_80mhz), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_562[55]), .CK(clk_80mhz), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_562[56]), .CK(clk_80mhz), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_562[57]), .CK(clk_80mhz), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_562[58]), .CK(clk_80mhz), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_562[59]), .CK(clk_80mhz), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_562[60]), .CK(clk_80mhz), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_562[61]), .CK(clk_80mhz), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_562[62]), .CK(clk_80mhz), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_562[63]), .CK(clk_80mhz), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_562[64]), .CK(clk_80mhz), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_562[65]), .CK(clk_80mhz), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_562[66]), .CK(clk_80mhz), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_562[67]), .CK(clk_80mhz), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_562[68]), .CK(clk_80mhz), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_562[69]), .CK(clk_80mhz), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_562[70]), .CK(clk_80mhz), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_562[71]), .CK(clk_80mhz), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_634[1]), .CK(clk_80mhz), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_634[2]), .CK(clk_80mhz), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_634[3]), .CK(clk_80mhz), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_634[4]), .CK(clk_80mhz), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_634[5]), .CK(clk_80mhz), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_634[6]), .CK(clk_80mhz), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_634[7]), .CK(clk_80mhz), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_634[8]), .CK(clk_80mhz), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_634[9]), .CK(clk_80mhz), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_634[10]), .CK(clk_80mhz), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_634[11]), .CK(clk_80mhz), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_634[12]), .CK(clk_80mhz), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_634[13]), .CK(clk_80mhz), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_634[14]), .CK(clk_80mhz), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_634[15]), .CK(clk_80mhz), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_634[16]), .CK(clk_80mhz), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_634[17]), .CK(clk_80mhz), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_634[18]), .CK(clk_80mhz), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_634[19]), .CK(clk_80mhz), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_634[20]), .CK(clk_80mhz), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_634[21]), .CK(clk_80mhz), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_634[22]), .CK(clk_80mhz), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_634[23]), .CK(clk_80mhz), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_634[24]), .CK(clk_80mhz), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_634[25]), .CK(clk_80mhz), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_634[26]), .CK(clk_80mhz), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_634[27]), .CK(clk_80mhz), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_634[28]), .CK(clk_80mhz), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_634[29]), .CK(clk_80mhz), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_634[30]), .CK(clk_80mhz), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_634[31]), .CK(clk_80mhz), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_634[32]), .CK(clk_80mhz), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_634[33]), .CK(clk_80mhz), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_634[34]), .CK(clk_80mhz), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_634[35]), .CK(clk_80mhz), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_634[36]), .CK(clk_80mhz), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_634[37]), .CK(clk_80mhz), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_634[38]), .CK(clk_80mhz), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_634[39]), .CK(clk_80mhz), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_634[40]), .CK(clk_80mhz), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_634[41]), .CK(clk_80mhz), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_634[42]), .CK(clk_80mhz), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_634[43]), .CK(clk_80mhz), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_634[44]), .CK(clk_80mhz), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_634[45]), .CK(clk_80mhz), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_634[46]), .CK(clk_80mhz), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_634[47]), .CK(clk_80mhz), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_634[48]), .CK(clk_80mhz), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_634[49]), .CK(clk_80mhz), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_634[50]), .CK(clk_80mhz), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_634[51]), .CK(clk_80mhz), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_634[52]), .CK(clk_80mhz), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_634[53]), .CK(clk_80mhz), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_634[54]), .CK(clk_80mhz), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_634[55]), .CK(clk_80mhz), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_634[56]), .CK(clk_80mhz), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_634[57]), .CK(clk_80mhz), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_634[58]), .CK(clk_80mhz), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_634[59]), .CK(clk_80mhz), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_634[60]), .CK(clk_80mhz), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_634[61]), .CK(clk_80mhz), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_634[62]), .CK(clk_80mhz), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_634[63]), .CK(clk_80mhz), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_634[64]), .CK(clk_80mhz), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_634[65]), .CK(clk_80mhz), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_634[66]), .CK(clk_80mhz), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_634[67]), .CK(clk_80mhz), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_634[68]), .CK(clk_80mhz), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_634[69]), .CK(clk_80mhz), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_634[70]), .CK(clk_80mhz), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_634[71]), .CK(clk_80mhz), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_706[1]), .CK(clk_80mhz), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_706[2]), .CK(clk_80mhz), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_706[3]), .CK(clk_80mhz), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_706[4]), .CK(clk_80mhz), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_706[5]), .CK(clk_80mhz), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_706[6]), .CK(clk_80mhz), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_706[7]), .CK(clk_80mhz), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_706[8]), .CK(clk_80mhz), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_706[9]), .CK(clk_80mhz), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_706[10]), .CK(clk_80mhz), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_706[11]), .CK(clk_80mhz), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_706[12]), .CK(clk_80mhz), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_706[13]), .CK(clk_80mhz), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_706[14]), .CK(clk_80mhz), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_706[15]), .CK(clk_80mhz), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_706[16]), .CK(clk_80mhz), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_706[17]), .CK(clk_80mhz), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_706[18]), .CK(clk_80mhz), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_706[19]), .CK(clk_80mhz), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_706[20]), .CK(clk_80mhz), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_706[21]), .CK(clk_80mhz), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_706[22]), .CK(clk_80mhz), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_706[23]), .CK(clk_80mhz), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_706[24]), .CK(clk_80mhz), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_706[25]), .CK(clk_80mhz), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_706[26]), .CK(clk_80mhz), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_706[27]), .CK(clk_80mhz), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_706[28]), .CK(clk_80mhz), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_706[29]), .CK(clk_80mhz), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_706[30]), .CK(clk_80mhz), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_706[31]), .CK(clk_80mhz), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_706[32]), .CK(clk_80mhz), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_706[33]), .CK(clk_80mhz), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_706[34]), .CK(clk_80mhz), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_706[35]), .CK(clk_80mhz), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_706[36]), .CK(clk_80mhz), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_706[37]), .CK(clk_80mhz), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_706[38]), .CK(clk_80mhz), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_706[39]), .CK(clk_80mhz), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_706[40]), .CK(clk_80mhz), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_706[41]), .CK(clk_80mhz), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_706[42]), .CK(clk_80mhz), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_706[43]), .CK(clk_80mhz), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_706[44]), .CK(clk_80mhz), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_706[45]), .CK(clk_80mhz), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_706[46]), .CK(clk_80mhz), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_706[47]), .CK(clk_80mhz), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_706[48]), .CK(clk_80mhz), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_706[49]), .CK(clk_80mhz), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_706[50]), .CK(clk_80mhz), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_706[51]), .CK(clk_80mhz), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_706[52]), .CK(clk_80mhz), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_706[53]), .CK(clk_80mhz), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_706[54]), .CK(clk_80mhz), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_706[55]), .CK(clk_80mhz), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_706[56]), .CK(clk_80mhz), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_706[57]), .CK(clk_80mhz), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_706[58]), .CK(clk_80mhz), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_706[59]), .CK(clk_80mhz), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_706[60]), .CK(clk_80mhz), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_706[61]), .CK(clk_80mhz), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_706[62]), .CK(clk_80mhz), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_706[63]), .CK(clk_80mhz), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_706[64]), .CK(clk_80mhz), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_706[65]), .CK(clk_80mhz), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_706[66]), .CK(clk_80mhz), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_706[67]), .CK(clk_80mhz), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_706[68]), .CK(clk_80mhz), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_706[69]), .CK(clk_80mhz), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_706[70]), .CK(clk_80mhz), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_706[71]), .CK(clk_80mhz), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1459[1]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1459[2]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1459[3]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1459[4]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1459[5]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1459[6]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1459[7]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1459[8]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1459[9]), .SP(clk_80mhz_enable_806), .CK(clk_80mhz), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1459[10]), .SP(clk_80mhz_enable_806), 
            .CK(clk_80mhz), .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1459[11]), .SP(clk_80mhz_enable_806), 
            .CK(clk_80mhz), .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1459[12]), .SP(clk_80mhz_enable_806), 
            .CK(clk_80mhz), .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1459[13]), .SP(clk_80mhz_enable_806), 
            .CK(clk_80mhz), .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1459[14]), .SP(clk_80mhz_enable_806), 
            .CK(clk_80mhz), .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1459[15]), .SP(clk_80mhz_enable_806), 
            .CK(clk_80mhz), .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1459[16]), .SP(clk_80mhz_enable_806), 
            .CK(clk_80mhz), .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1459[17]), .SP(clk_80mhz_enable_806), 
            .CK(clk_80mhz), .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1459[18]), .SP(clk_80mhz_enable_806), 
            .CK(clk_80mhz), .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1459[19]), .SP(clk_80mhz_enable_806), 
            .CK(clk_80mhz), .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1459[20]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1459[21]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1459[22]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1459[23]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1459[24]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1459[25]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1459[26]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1459[27]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1459[28]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1459[29]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1459[30]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1459[31]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1459[32]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1459[33]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1459[34]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1459[35]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1459[36]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1459[37]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1459[38]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1459[39]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1459[40]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1459[41]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1459[42]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1459[43]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1459[44]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1459[45]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1459[46]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1459[47]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1459[48]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1459[49]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1459[50]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1459[51]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1459[52]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1459[53]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1459[54]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1459[55]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1459[56]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1459[57]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1459[58]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1459[59]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1459[60]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1459[61]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1459[62]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1459[63]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1459[64]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1459[65]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1459[66]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1459[67]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1459[68]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1459[69]), .SP(clk_80mhz_enable_856), 
            .CK(clk_80mhz), .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1459[70]), .SP(clk_80mhz_enable_906), 
            .CK(clk_80mhz), .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1459[71]), .SP(clk_80mhz_enable_906), 
            .CK(clk_80mhz), .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(clk_80mhz_enable_906), .CK(clk_80mhz), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1531[1]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1531[2]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1531[3]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1531[4]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1531[5]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1531[6]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1531[7]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1531[8]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1531[9]), .SP(clk_80mhz_enable_956), .CK(clk_80mhz), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1531[10]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1531[11]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1531[12]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1531[13]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1531[14]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1531[15]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1531[16]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1531[17]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1531[18]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1531[19]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1531[20]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1531[21]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1531[22]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1531[23]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1531[24]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1531[25]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1531[26]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1531[27]), .SP(clk_80mhz_enable_956), 
            .CK(clk_80mhz), .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1531[28]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1531[29]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1531[30]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1531[31]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1531[32]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1531[33]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1531[34]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1531[35]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1531[36]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1531[37]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1531[38]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1531[39]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1531[40]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1531[41]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1531[42]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1531[43]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1531[44]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1531[45]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1531[46]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1531[47]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1531[48]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1531[49]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1531[50]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1531[51]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1531[52]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1531[53]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1531[54]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1531[55]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1531[56]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1531[57]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1531[58]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1531[59]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1531[60]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1531[61]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1531[62]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1531[63]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1531[64]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1531[65]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1531[66]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1531[67]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1531[68]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1531[69]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1531[70]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1531[71]), .SP(clk_80mhz_enable_1006), 
            .CK(clk_80mhz), .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(clk_80mhz_enable_1006), .CK(clk_80mhz), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(clk_80mhz_enable_1006), .CK(clk_80mhz), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(clk_80mhz_enable_1006), .CK(clk_80mhz), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(clk_80mhz_enable_1006), .CK(clk_80mhz), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(clk_80mhz_enable_1006), .CK(clk_80mhz), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(clk_80mhz_enable_1006), .CK(clk_80mhz), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(clk_80mhz_enable_1056), .CK(clk_80mhz), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(clk_80mhz_enable_1106), .CK(clk_80mhz), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1603[1]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1603[2]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1603[3]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1603[4]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1603[5]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1603[6]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1603[7]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1603[8]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1603[9]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1603[10]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1603[11]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1603[12]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1603[13]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1603[14]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1603[15]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1603[16]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1603[17]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1603[18]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1603[19]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1603[20]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1603[21]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1603[22]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1603[23]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1603[24]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1603[25]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1603[26]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1603[27]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1603[28]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1603[29]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1603[30]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1603[31]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1603[32]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1603[33]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1603[34]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1603[35]), .SP(clk_80mhz_enable_1106), 
            .CK(clk_80mhz), .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1603[36]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1603[37]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1603[38]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1603[39]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1603[40]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1603[41]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1603[42]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1603[43]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1603[44]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1603[45]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1603[46]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1603[47]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1603[48]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1603[49]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1603[50]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1603[51]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1603[52]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1603[53]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1603[54]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1603[55]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1603[56]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1603[57]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1603[58]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1603[59]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1603[60]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1603[61]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1603[62]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1603[63]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1603[64]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1603[65]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1603[66]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1603[67]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1603[68]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1603[69]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1603[70]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1603[71]), .SP(clk_80mhz_enable_1156), 
            .CK(clk_80mhz), .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(clk_80mhz_enable_1156), .CK(clk_80mhz), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(clk_80mhz_enable_1206), .CK(clk_80mhz), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(clk_80mhz_enable_1256), .CK(clk_80mhz), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(clk_80mhz_enable_1256), .CK(clk_80mhz), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(clk_80mhz_enable_1256), .CK(clk_80mhz), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(clk_80mhz_enable_1256), .CK(clk_80mhz), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(clk_80mhz_enable_1256), .CK(clk_80mhz), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(clk_80mhz_enable_1256), .CK(clk_80mhz), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(clk_80mhz_enable_1256), .CK(clk_80mhz), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1675[1]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1675[2]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1675[3]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1675[4]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1675[5]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1675[6]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1675[7]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1675[8]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1675[9]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1675[10]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1675[11]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1675[12]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1675[13]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1675[14]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1675[15]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1675[16]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1675[17]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1675[18]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1675[19]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1675[20]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1675[21]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1675[22]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1675[23]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1675[24]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1675[25]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1675[26]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1675[27]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1675[28]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1675[29]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1675[30]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1675[31]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1675[32]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1675[33]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1675[34]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1675[35]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1675[36]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1675[37]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1675[38]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1675[39]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1675[40]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1675[41]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1675[42]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1675[43]), .SP(clk_80mhz_enable_1256), 
            .CK(clk_80mhz), .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1675[44]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1675[45]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1675[46]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1675[47]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1675[48]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1675[49]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1675[50]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1675[51]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1675[52]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1675[53]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1675[54]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1675[55]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1675[56]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1675[57]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1675[58]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1675[59]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1675[60]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1675[61]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1675[62]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1675[63]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1675[64]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1675[65]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1675[66]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1675[67]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1675[68]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1675[69]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1675[70]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1675[71]), .SP(clk_80mhz_enable_1306), 
            .CK(clk_80mhz), .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(clk_80mhz_enable_1306), .CK(clk_80mhz), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(clk_80mhz_enable_1356), .CK(clk_80mhz), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1747[57]), .SP(clk_80mhz_enable_1356), 
            .CK(clk_80mhz), .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1747[58]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1747[59]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1747[60]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1747[61]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[61] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1747[62]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[62] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1747[63]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[63] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1747[64]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[64] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1747[65]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[65] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1747[66]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[66] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1747[67]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[67] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1747[68]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[68] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1747[69]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[69] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1747[70]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[70] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1747[71]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[71] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1819[1]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(\d_out_11__N_1819[2] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(\d_out_11__N_1819[3] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(\d_out_11__N_1819[4] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(\d_out_11__N_1819[5] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(\d_out_11__N_1819[6] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(\d_out_11__N_1819[7] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(\d_out_11__N_1819[8] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(\d_out_11__N_1819[9] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(\d_out_11__N_1819[10] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(\d_out_11__N_1819[11] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_418[1]), .CK(clk_80mhz), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_418[2]), .CK(clk_80mhz), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_418[3]), .CK(clk_80mhz), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_418[4]), .CK(clk_80mhz), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_418[5]), .CK(clk_80mhz), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_418[6]), .CK(clk_80mhz), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_418[7]), .CK(clk_80mhz), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_418[8]), .CK(clk_80mhz), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_418[9]), .CK(clk_80mhz), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_418[10]), .CK(clk_80mhz), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_418[11]), .CK(clk_80mhz), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_418[12]), .CK(clk_80mhz), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_418[13]), .CK(clk_80mhz), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_418[14]), .CK(clk_80mhz), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_418[15]), .CK(clk_80mhz), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_418[16]), .CK(clk_80mhz), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_418[17]), .CK(clk_80mhz), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_418[18]), .CK(clk_80mhz), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_418[19]), .CK(clk_80mhz), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_418[20]), .CK(clk_80mhz), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_418[21]), .CK(clk_80mhz), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_418[22]), .CK(clk_80mhz), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_418[23]), .CK(clk_80mhz), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_418[24]), .CK(clk_80mhz), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_418[25]), .CK(clk_80mhz), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_418[26]), .CK(clk_80mhz), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_418[27]), .CK(clk_80mhz), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_418[28]), .CK(clk_80mhz), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_418[29]), .CK(clk_80mhz), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_418[30]), .CK(clk_80mhz), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_418[31]), .CK(clk_80mhz), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_418[32]), .CK(clk_80mhz), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_418[33]), .CK(clk_80mhz), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_418[34]), .CK(clk_80mhz), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_418[35]), .CK(clk_80mhz), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_418[36]), .CK(clk_80mhz), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_418[37]), .CK(clk_80mhz), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_418[38]), .CK(clk_80mhz), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_418[39]), .CK(clk_80mhz), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_418[40]), .CK(clk_80mhz), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_418[41]), .CK(clk_80mhz), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_418[42]), .CK(clk_80mhz), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_418[43]), .CK(clk_80mhz), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_418[44]), .CK(clk_80mhz), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_418[45]), .CK(clk_80mhz), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_418[46]), .CK(clk_80mhz), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_418[47]), .CK(clk_80mhz), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_418[48]), .CK(clk_80mhz), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_418[49]), .CK(clk_80mhz), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_418[50]), .CK(clk_80mhz), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_418[51]), .CK(clk_80mhz), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_418[52]), .CK(clk_80mhz), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_418[53]), .CK(clk_80mhz), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_418[54]), .CK(clk_80mhz), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_418[55]), .CK(clk_80mhz), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_418[56]), .CK(clk_80mhz), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_418[57]), .CK(clk_80mhz), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_418[58]), .CK(clk_80mhz), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_418[59]), .CK(clk_80mhz), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_418[60]), .CK(clk_80mhz), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_418[61]), .CK(clk_80mhz), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_418[62]), .CK(clk_80mhz), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_418[63]), .CK(clk_80mhz), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_418[64]), .CK(clk_80mhz), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_418[65]), .CK(clk_80mhz), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_418[66]), .CK(clk_80mhz), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_418[67]), .CK(clk_80mhz), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_418[68]), .CK(clk_80mhz), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_418[69]), .CK(clk_80mhz), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_418[70]), .CK(clk_80mhz), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_418[71]), .CK(clk_80mhz), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i71.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i63_1_lut (.A(d_d8[62]), .Z(n11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 i6080_else_3_lut (.A(n17325), .B(\CICGain[1] ), .C(\d10[59] ), 
         .Z(n17857)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6080_else_3_lut.init = 16'he2e2;
    LUT4 i3135_2_lut_3_lut (.A(n17191), .B(n16826), .C(n87_adj_228[11]), 
         .Z(count_15__N_1442[11])) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(74[22:52])
    defparam i3135_2_lut_3_lut.init = 16'hf1f1;
    LUT4 i3090_2_lut_3_lut (.A(n17191), .B(n16826), .C(n87_adj_228[0]), 
         .Z(count_15__N_1442[0])) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(74[22:52])
    defparam i3090_2_lut_3_lut.init = 16'hf1f1;
    LUT4 sub_28_inv_0_i64_1_lut (.A(d_d8[63]), .Z(n10_adj_117)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i61_1_lut (.A(d_d8[60]), .Z(n13_adj_118)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i62_1_lut (.A(d_d8[61]), .Z(n12_adj_119)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i59_1_lut (.A(d_d8[58]), .Z(n15_adj_120)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i60_1_lut (.A(d_d8[59]), .Z(n14_adj_121)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i57_1_lut (.A(d_d8[56]), .Z(n17_adj_122)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i58_1_lut (.A(d_d8[57]), .Z(n16_adj_123)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i55_1_lut (.A(d_d8[54]), .Z(n19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i56_1_lut (.A(d_d8[55]), .Z(n18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i53_1_lut (.A(d_d8[52]), .Z(n21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i54_1_lut (.A(d_d8[53]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i51_1_lut (.A(d_d8[50]), .Z(n23_adj_124)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i52_1_lut (.A(d_d8[51]), .Z(n22_adj_125)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i49_1_lut (.A(d_d8[48]), .Z(n25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i50_1_lut (.A(d_d8[49]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 i6052_then_3_lut (.A(\CICGain[1] ), .B(\d10[59] ), .C(d10[57]), 
         .Z(n17876)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6052_then_3_lut.init = 16'he4e4;
    LUT4 sub_28_inv_0_i47_1_lut (.A(d_d8[46]), .Z(n27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i48_1_lut (.A(d_d8[47]), .Z(n26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i43_1_lut (.A(d_d6[42]), .Z(n31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i44_1_lut (.A(d_d6[43]), .Z(n30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i45_1_lut (.A(d_d8[44]), .Z(n29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i46_1_lut (.A(d_d8[45]), .Z(n28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 i6052_else_3_lut (.A(n17302), .B(\CICGain[1] ), .C(d10[58]), 
         .Z(n17875)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6052_else_3_lut.init = 16'he2e2;
    LUT4 sub_26_inv_0_i41_1_lut (.A(d_d6[40]), .Z(n33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i43_1_lut (.A(d_d8[42]), .Z(n31_adj_126)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i42_1_lut (.A(d_d6[41]), .Z(n32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i44_1_lut (.A(d_d8[43]), .Z(n30_adj_127)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i41_1_lut (.A(d_d8[40]), .Z(n33_adj_128)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i55_1_lut (.A(d_d6[54]), .Z(n19_adj_129)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i42_1_lut (.A(d_d8[41]), .Z(n32_adj_130)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i39_1_lut (.A(d_d8[38]), .Z(n35_adj_131)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i39_1_lut (.A(d_d6[38]), .Z(n35_adj_132)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i40_1_lut (.A(d_d6[39]), .Z(n34_adj_133)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i56_1_lut (.A(d_d6[55]), .Z(n18_adj_134)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i40_1_lut (.A(d_d8[39]), .Z(n34_adj_135)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i37_1_lut (.A(d_d8[36]), .Z(n37_adj_136)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i38_1_lut (.A(d_d8[37]), .Z(n36_adj_137)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i71_1_lut (.A(d_d_tmp[70]), .Z(n3_adj_138)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i72_1_lut (.A(d_d_tmp[71]), .Z(n2_adj_139)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i69_1_lut (.A(d_d_tmp[68]), .Z(n5_adj_140)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i37_1_lut (.A(d_d6[36]), .Z(n37_adj_141)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i38_1_lut (.A(d_d6[37]), .Z(n36_adj_142)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i70_1_lut (.A(d_d_tmp[69]), .Z(n4_adj_143)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i67_1_lut (.A(d_d_tmp[66]), .Z(n7_adj_144)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i68_1_lut (.A(d_d_tmp[67]), .Z(n6_adj_145)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i65_1_lut (.A(d_d_tmp[64]), .Z(n9_adj_146)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i66_1_lut (.A(d_d_tmp[65]), .Z(n8_adj_147)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i63_1_lut (.A(d_d_tmp[62]), .Z(n11_adj_148)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i64_1_lut (.A(d_d_tmp[63]), .Z(n10_adj_149)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i61_1_lut (.A(d_d_tmp[60]), .Z(n13_adj_150)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i62_1_lut (.A(d_d_tmp[61]), .Z(n12_adj_151)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i59_1_lut (.A(d_d_tmp[58]), .Z(n15_adj_152)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i60_1_lut (.A(d_d_tmp[59]), .Z(n14_adj_153)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i57_1_lut (.A(d_d_tmp[56]), .Z(n17_adj_154)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i58_1_lut (.A(d_d_tmp[57]), .Z(n16_adj_155)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i55_1_lut (.A(d_d_tmp[54]), .Z(n19_adj_156)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i56_1_lut (.A(d_d_tmp[55]), .Z(n18_adj_157)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i53_1_lut (.A(d_d_tmp[52]), .Z(n21_adj_158)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i54_1_lut (.A(d_d_tmp[53]), .Z(n20_adj_159)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i51_1_lut (.A(d_d_tmp[50]), .Z(n23_adj_160)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i52_1_lut (.A(d_d_tmp[51]), .Z(n22_adj_161)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i49_1_lut (.A(d_d_tmp[48]), .Z(n25_adj_162)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i50_1_lut (.A(d_d_tmp[49]), .Z(n24_adj_163)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i47_1_lut (.A(d_d_tmp[46]), .Z(n27_adj_164)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i48_1_lut (.A(d_d_tmp[47]), .Z(n26_adj_165)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i45_1_lut (.A(d_d_tmp[44]), .Z(n29_adj_166)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i46_1_lut (.A(d_d_tmp[45]), .Z(n28_adj_167)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i46_1_lut.init = 16'h5555;
    FD1S3IX count__i2 (.D(n87_adj_228[2]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n87_adj_228[3]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n87_adj_228[4]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n87_adj_228[5]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n87_adj_228[6]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n87_adj_228[7]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n87_adj_228[8]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n87_adj_228[9]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n87_adj_228[10]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1442[11]), .CK(clk_80mhz), .CD(count_15__N_1458), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n87_adj_228[12]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n87_adj_228[13]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n87_adj_228[14]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n87_adj_228[15]), .CK(clk_80mhz), .CD(n12783), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i15.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i43_1_lut (.A(d_d_tmp[42]), .Z(n31_adj_168)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i44_1_lut (.A(d_d_tmp[43]), .Z(n30_adj_169)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i41_1_lut (.A(d_d_tmp[40]), .Z(n33_adj_170)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i41_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_245 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_806)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_245.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(count[14]), .B(count[13]), .Z(n17193)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 sub_26_inv_0_i69_1_lut (.A(d_d6[68]), .Z(n5_adj_171)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i70_1_lut (.A(d_d6[69]), .Z(n4_adj_172)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i67_1_lut (.A(d_d6[66]), .Z(n7_adj_173)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i68_1_lut (.A(d_d6[67]), .Z(n6_adj_174)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i71_1_lut (.A(d_d6[70]), .Z(n3_adj_175)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i72_1_lut (.A(d_d6[71]), .Z(n2_adj_176)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i71_1_lut (.A(d_d7[70]), .Z(n3_adj_177)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i72_1_lut (.A(d_d7[71]), .Z(n2_adj_178)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i61_1_lut (.A(d_d7[60]), .Z(n13_adj_179)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i62_1_lut (.A(d_d7[61]), .Z(n12_adj_180)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i59_1_lut (.A(d_d7[58]), .Z(n15_adj_181)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i60_1_lut (.A(d_d7[59]), .Z(n14_adj_182)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i42_1_lut (.A(d_d_tmp[41]), .Z(n32_adj_183)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i39_1_lut (.A(d_d_tmp[38]), .Z(n35_adj_184)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i40_1_lut (.A(d_d_tmp[39]), .Z(n34_adj_185)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 mux_1200_i2_3_lut (.A(n118), .B(n120), .C(cout), .Z(d10_71__N_1747[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1200_i3_3_lut (.A(n115), .B(n117), .C(cout), .Z(d10_71__N_1747[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1200_i4_3_lut (.A(n112), .B(n114), .C(cout), .Z(d10_71__N_1747[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1200_i5_3_lut (.A(n109), .B(n111), .C(cout), .Z(d10_71__N_1747[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1200_i6_3_lut (.A(n106), .B(n108), .C(cout), .Z(d10_71__N_1747[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i6_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i57_1_lut (.A(d_d7[56]), .Z(n17_adj_186)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 mux_1200_i7_3_lut (.A(n103), .B(n105), .C(cout), .Z(d10_71__N_1747[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1200_i8_3_lut (.A(n100), .B(n102), .C(cout), .Z(d10_71__N_1747[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1200_i9_3_lut (.A(n97), .B(n99), .C(cout), .Z(d10_71__N_1747[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1200_i10_3_lut (.A(n94), .B(n96), .C(cout), .Z(d10_71__N_1747[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i10_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i69_1_lut (.A(d_d7[68]), .Z(n5_adj_187)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 mux_1200_i11_3_lut (.A(n91), .B(n93), .C(cout), .Z(d10_71__N_1747[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i11_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i58_1_lut (.A(d_d7[57]), .Z(n16_adj_188)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i55_1_lut (.A(d_d7[54]), .Z(n19_adj_189)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i56_1_lut (.A(d_d7[55]), .Z(n18_adj_190)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 mux_1200_i12_3_lut (.A(n88), .B(n90), .C(cout), .Z(d10_71__N_1747[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i12_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i53_1_lut (.A(d_d7[52]), .Z(n21_adj_191)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i54_1_lut (.A(d_d7[53]), .Z(n20_adj_192)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i51_1_lut (.A(d_d7[50]), .Z(n23_adj_193)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i52_1_lut (.A(d_d7[51]), .Z(n22_adj_194)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i49_1_lut (.A(d_d7[48]), .Z(n25_adj_195)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i50_1_lut (.A(d_d7[49]), .Z(n24_adj_196)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i47_1_lut (.A(d_d7[46]), .Z(n27_adj_197)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i48_1_lut (.A(d_d7[47]), .Z(n26_adj_198)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i48_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_244 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_756)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_244.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i49_1_lut (.A(d_d6[48]), .Z(n25_adj_199)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i70_1_lut (.A(d_d7[69]), .Z(n4_adj_200)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i67_1_lut (.A(d_d7[66]), .Z(n7_adj_201)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i45_1_lut (.A(d_d7[44]), .Z(n29_adj_202)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i53_1_lut (.A(d_d6[52]), .Z(n21_adj_203)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i46_1_lut (.A(d_d7[45]), .Z(n28_adj_204)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i61_rep_33_3_lut (.A(\d10[60] ), .B(\d10[61] ), 
         .C(\CICGain[0] ), .Z(n17302)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i61_rep_33_3_lut.init = 16'hcaca;
    LUT4 mux_1200_i13_3_lut (.A(n85), .B(n87), .C(cout), .Z(d10_71__N_1747[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1200_i14_3_lut (.A(n82), .B(n84), .C(cout), .Z(d10_71__N_1747[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i14_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i54_1_lut (.A(d_d6[53]), .Z(n20_adj_205)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i43_1_lut (.A(d_d7[42]), .Z(n31_adj_206)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i68_1_lut (.A(d_d7[67]), .Z(n6_adj_207)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 i5956_2_lut (.A(n17268), .B(n16826), .Z(count_15__N_1458)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(69[13:41])
    defparam i5956_2_lut.init = 16'h2222;
    LUT4 sub_27_inv_0_i44_1_lut (.A(d_d7[43]), .Z(n30_adj_208)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 i5881_4_lut (.A(n17225), .B(n17262), .C(n17219), .D(count[4]), 
         .Z(n17268)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5881_4_lut.init = 16'h8000;
    LUT4 sub_26_inv_0_i47_1_lut (.A(d_d6[46]), .Z(n27_adj_209)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i48_1_lut (.A(d_d6[47]), .Z(n26_adj_210)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i45_1_lut (.A(d_d6[44]), .Z(n29_adj_211)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i46_1_lut (.A(d_d6[45]), .Z(n28_adj_212)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 mux_1200_i15_3_lut (.A(n79), .B(n81_adj_213), .C(cout), .Z(d10_71__N_1747[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i15_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i65_1_lut (.A(d_d7[64]), .Z(n9_adj_214)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 i1_4_lut (.A(count[10]), .B(count[0]), .C(count[7]), .D(count[5]), 
         .Z(n17225)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'h8000;
    LUT4 sub_26_inv_0_i65_1_lut (.A(d_d6[64]), .Z(n9_adj_215)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i66_1_lut (.A(d_d6[65]), .Z(n8_adj_216)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 mux_1200_i16_3_lut (.A(n76), .B(n78_adj_217), .C(cout), .Z(d10_71__N_1747[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1200_i16_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i42_1_lut (.A(d_d7[41]), .Z(n32_adj_218)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 i5875_4_lut (.A(count[1]), .B(count[2]), .C(count[8]), .D(count[3]), 
         .Z(n17262)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5875_4_lut.init = 16'h8000;
    LUT4 sub_27_inv_0_i41_1_lut (.A(d_d7[40]), .Z(n33_adj_219)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i62_rep_56_3_lut (.A(\d10[61] ), .B(\d10[62] ), 
         .C(\CICGain[0] ), .Z(n17325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i62_rep_56_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i63_3_lut (.A(\d10[62] ), .B(\d10[63] ), .C(\CICGain[0] ), 
         .Z(n63_adj_220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_50 (.A(count[6]), .B(count[9]), .Z(n17219)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_50.init = 16'h8888;
    LUT4 i1_4_lut_adj_51 (.A(count[12]), .B(count[11]), .C(n17193), .D(count[15]), 
         .Z(n16826)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_51.init = 16'hfffb;
    LUT4 sub_26_inv_0_i63_1_lut (.A(d_d6[62]), .Z(n11_adj_221)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i63_1_lut.init = 16'h5555;
    PFUMX i6120 (.BLUT(n17875), .ALUT(n17876), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[0]));
    LUT4 shift_right_31_i64_rep_18_3_lut (.A(\d10[63] ), .B(\d10[64] ), 
         .C(\CICGain[0] ), .Z(n17288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i64_rep_18_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i65_3_lut (.A(\d10[64] ), .B(\d10[65] ), .C(\CICGain[0] ), 
         .Z(n65)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i66_1_lut (.A(d_d7[65]), .Z(n8_adj_222)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i66_3_lut (.A(\d10[65] ), .B(\d10[66] ), .C(\CICGain[0] ), 
         .Z(n66_adj_223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i63_1_lut (.A(d_d7[62]), .Z(n11_adj_224)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i37_1_lut (.A(d_d_tmp[36]), .Z(n37_adj_225)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i38_1_lut (.A(d_d_tmp[37]), .Z(n36_adj_226)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i50_1_lut (.A(d_d6[49]), .Z(n24_adj_227)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i50_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_256 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_1356)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_256.GSR = "ENABLED";
    LUT4 i6037_3_lut (.A(n16826), .B(n17191), .C(n17268), .Z(n12783)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam i6037_3_lut.init = 16'h5151;
    FD1S3AX v_comb_66_rep_255 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_1306)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_255.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_52 (.A(n17189), .B(count[10]), .C(n17181), .D(count[7]), 
         .Z(n17191)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(74[22:52])
    defparam i1_4_lut_adj_52.init = 16'hfffe;
    FD1S3AX v_comb_66_rep_254 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_1256)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_254.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_53 (.A(count[8]), .B(n17185), .C(count[1]), .D(count[9]), 
         .Z(n17189)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(74[22:52])
    defparam i1_4_lut_adj_53.init = 16'hfffe;
    LUT4 i1_2_lut_adj_54 (.A(count[6]), .B(count[5]), .Z(n17181)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(74[22:52])
    defparam i1_2_lut_adj_54.init = 16'heeee;
    PFUMX i6108 (.BLUT(n17857), .ALUT(n17858), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[1]));
    LUT4 i1_4_lut_adj_55 (.A(count[2]), .B(count[4]), .C(count[0]), .D(count[3]), 
         .Z(n17185)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(74[22:52])
    defparam i1_4_lut_adj_55.init = 16'hfffe;
    FD1S3AX v_comb_66_rep_253 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_1206)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_253.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_252 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_1156)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_252.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_251 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_1106)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_251.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_250 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_1056)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_250.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_249 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_1006)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_249.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_248 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_956)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_248.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_247 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_906)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_247.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_246 (.D(count_15__N_1458), .CK(clk_80mhz), .Q(clk_80mhz_enable_856)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_246.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \CIC(WIDTH=72,DECIMATION_RATIO=4096)_U0 
//

module \CIC(WIDTH=72,DECIMATION_RATIO=4096)_U0  (d_d7, n15, d_tmp, clk_80mhz, 
            d5, d_d_tmp, d2, d2_71__N_490, n13, n12, n14, d3, 
            d3_71__N_562, count, n87_adj_114, d4, d4_71__N_634, d5_71__N_706, 
            d6, d6_71__N_1459, d_d6, CIC1_out_clkSin, d7, d7_71__N_1531, 
            d8, d8_71__N_1603, d_d8, d9, d9_71__N_1675, d_d9, n17, 
            MultDataB, d1, d1_71__N_418, n16, n15_adj_1, n19, n14_adj_2, 
            n17_adj_3, n16_adj_4, n18, n19_adj_5, n21, n20, n18_adj_6, 
            n23, n22, n21_adj_7, n25, n24, n27, n20_adj_8, n23_adj_9, 
            n22_adj_10, n26, n29, n25_adj_11, n28, n24_adj_12, n27_adj_13, 
            n26_adj_14, n31, n29_adj_15, n28_adj_16, n31_adj_17, n30, 
            n30_adj_18, n33, n32, n33_adj_19, n32_adj_20, n35, n34, 
            n35_adj_21, n37, n36_adj_22, n34_adj_23, n37_adj_24, n36_adj_25, 
            \CICGain[1] , \CICGain[0] , \d10[66] , \d10[67] , \d10[69] , 
            \d10[68] , n3, n2, \d10[65] , n5, \d10[70] , n4, \d10[71] , 
            n7, n6, n9, n8, n11, n10, n13_adj_26, n118, n120, 
            cout, n115, n117, n112, n114, n3_adj_27, n109, n111, 
            n2_adj_28, n5_adj_29, n63_adj_30, \d_out_11__N_1819[2] , 
            n4_adj_31, n12_adj_32, n7_adj_33, n6_adj_34, n9_adj_35, 
            n17288, \d_out_11__N_1819[3] , n65, \d_out_11__N_1819[4] , 
            n8_adj_36, n66_adj_37, \d_out_11__N_1819[5] , n11_adj_38, 
            \d_out_11__N_1819[6] , n10_adj_39, n13_adj_40, n12_adj_41, 
            n15_adj_42, n15_adj_43, n14_adj_44, \d_out_11__N_1819[7] , 
            n14_adj_45, n17_adj_46, n106, n108, n16_adj_47, n17_adj_48, 
            n16_adj_49, n19_adj_50, n18_adj_51, n21_adj_52, n20_adj_53, 
            n23_adj_54, n22_adj_55, n25_adj_56, n24_adj_57, n27_adj_58, 
            n26_adj_59, n29_adj_60, n28_adj_61, n31_adj_62, n30_adj_63, 
            n33_adj_64, n32_adj_65, n35_adj_66, n34_adj_67, n37_adj_68, 
            n36_adj_69, n19_adj_70, n18_adj_71, n21_adj_72, n20_adj_73, 
            n23_adj_74, n22_adj_75, n25_adj_76, n24_adj_77, n27_adj_78, 
            n26_adj_79, n29_adj_80, n28_adj_81, n31_adj_82, n30_adj_83, 
            n33_adj_84, n32_adj_85, n35_adj_86, n34_adj_87, n37_adj_88, 
            n36_adj_89, n103, n105, n3_adj_90, n2_adj_91, n100, 
            n102, n97, n99, n5_adj_92, n4_adj_93, n7_adj_94, n6_adj_95, 
            n9_adj_96, n94, n96, n8_adj_97, n91, n93, n11_adj_98, 
            n10_adj_99, n13_adj_100, n12_adj_101, n88, n90, n85, 
            n87, n82, n84, n79, n81_adj_102, n76, n78_adj_103, 
            \d10[63] , \d10[64] , \d10[62] , n17325, \d10[60] , \d10[61] , 
            n17302, \d10[59] , \d_out_11__N_1819[10] , \d_out_11__N_1819[11] , 
            \d_out_11__N_1819[8] , \d_out_11__N_1819[9] , n3_adj_104, 
            n2_adj_105, n5_adj_106, n4_adj_107, n7_adj_108, n6_adj_109, 
            n9_adj_110, n8_adj_111, n11_adj_112, n10_adj_113) /* synthesis syn_module_defined=1 */ ;
    output [71:0]d_d7;
    output n15;
    output [71:0]d_tmp;
    input clk_80mhz;
    output [71:0]d5;
    output [71:0]d_d_tmp;
    output [71:0]d2;
    input [71:0]d2_71__N_490;
    output n13;
    output n12;
    output n14;
    output [71:0]d3;
    input [71:0]d3_71__N_562;
    output [15:0]count;
    input [15:0]n87_adj_114;
    output [71:0]d4;
    input [71:0]d4_71__N_634;
    input [71:0]d5_71__N_706;
    output [71:0]d6;
    input [71:0]d6_71__N_1459;
    output [71:0]d_d6;
    output CIC1_out_clkSin;
    output [71:0]d7;
    input [71:0]d7_71__N_1531;
    output [71:0]d8;
    input [71:0]d8_71__N_1603;
    output [71:0]d_d8;
    output [71:0]d9;
    input [71:0]d9_71__N_1675;
    output [71:0]d_d9;
    output n17;
    output [11:0]MultDataB;
    output [71:0]d1;
    input [71:0]d1_71__N_418;
    output n16;
    output n15_adj_1;
    output n19;
    output n14_adj_2;
    output n17_adj_3;
    output n16_adj_4;
    output n18;
    output n19_adj_5;
    output n21;
    output n20;
    output n18_adj_6;
    output n23;
    output n22;
    output n21_adj_7;
    output n25;
    output n24;
    output n27;
    output n20_adj_8;
    output n23_adj_9;
    output n22_adj_10;
    output n26;
    output n29;
    output n25_adj_11;
    output n28;
    output n24_adj_12;
    output n27_adj_13;
    output n26_adj_14;
    output n31;
    output n29_adj_15;
    output n28_adj_16;
    output n31_adj_17;
    output n30;
    output n30_adj_18;
    output n33;
    output n32;
    output n33_adj_19;
    output n32_adj_20;
    output n35;
    output n34;
    output n35_adj_21;
    output n37;
    output n36_adj_22;
    output n34_adj_23;
    output n37_adj_24;
    output n36_adj_25;
    input \CICGain[1] ;
    input \CICGain[0] ;
    input \d10[66] ;
    input \d10[67] ;
    input \d10[69] ;
    input \d10[68] ;
    output n3;
    output n2;
    input \d10[65] ;
    output n5;
    input \d10[70] ;
    output n4;
    input \d10[71] ;
    output n7;
    output n6;
    output n9;
    output n8;
    output n11;
    output n10;
    output n13_adj_26;
    input n118;
    input n120;
    input cout;
    input n115;
    input n117;
    input n112;
    input n114;
    output n3_adj_27;
    input n109;
    input n111;
    output n2_adj_28;
    output n5_adj_29;
    input n63_adj_30;
    output \d_out_11__N_1819[2] ;
    output n4_adj_31;
    output n12_adj_32;
    output n7_adj_33;
    output n6_adj_34;
    output n9_adj_35;
    input n17288;
    output \d_out_11__N_1819[3] ;
    input n65;
    output \d_out_11__N_1819[4] ;
    output n8_adj_36;
    input n66_adj_37;
    output \d_out_11__N_1819[5] ;
    output n11_adj_38;
    output \d_out_11__N_1819[6] ;
    output n10_adj_39;
    output n13_adj_40;
    output n12_adj_41;
    output n15_adj_42;
    output n15_adj_43;
    output n14_adj_44;
    output \d_out_11__N_1819[7] ;
    output n14_adj_45;
    output n17_adj_46;
    input n106;
    input n108;
    output n16_adj_47;
    output n17_adj_48;
    output n16_adj_49;
    output n19_adj_50;
    output n18_adj_51;
    output n21_adj_52;
    output n20_adj_53;
    output n23_adj_54;
    output n22_adj_55;
    output n25_adj_56;
    output n24_adj_57;
    output n27_adj_58;
    output n26_adj_59;
    output n29_adj_60;
    output n28_adj_61;
    output n31_adj_62;
    output n30_adj_63;
    output n33_adj_64;
    output n32_adj_65;
    output n35_adj_66;
    output n34_adj_67;
    output n37_adj_68;
    output n36_adj_69;
    output n19_adj_70;
    output n18_adj_71;
    output n21_adj_72;
    output n20_adj_73;
    output n23_adj_74;
    output n22_adj_75;
    output n25_adj_76;
    output n24_adj_77;
    output n27_adj_78;
    output n26_adj_79;
    output n29_adj_80;
    output n28_adj_81;
    output n31_adj_82;
    output n30_adj_83;
    output n33_adj_84;
    output n32_adj_85;
    output n35_adj_86;
    output n34_adj_87;
    output n37_adj_88;
    output n36_adj_89;
    input n103;
    input n105;
    output n3_adj_90;
    output n2_adj_91;
    input n100;
    input n102;
    input n97;
    input n99;
    output n5_adj_92;
    output n4_adj_93;
    output n7_adj_94;
    output n6_adj_95;
    output n9_adj_96;
    input n94;
    input n96;
    output n8_adj_97;
    input n91;
    input n93;
    output n11_adj_98;
    output n10_adj_99;
    output n13_adj_100;
    output n12_adj_101;
    input n88;
    input n90;
    input n85;
    input n87;
    input n82;
    input n84;
    input n79;
    input n81_adj_102;
    input n76;
    input n78_adj_103;
    input \d10[63] ;
    input \d10[64] ;
    input \d10[62] ;
    input n17325;
    input \d10[60] ;
    input \d10[61] ;
    input n17302;
    input \d10[59] ;
    output \d_out_11__N_1819[10] ;
    output \d_out_11__N_1819[11] ;
    output \d_out_11__N_1819[8] ;
    output \d_out_11__N_1819[9] ;
    output n3_adj_104;
    output n2_adj_105;
    output n5_adj_106;
    output n4_adj_107;
    output n7_adj_108;
    output n6_adj_109;
    output n9_adj_110;
    output n8_adj_111;
    output n11_adj_112;
    output n10_adj_113;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(61[23:32])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(74[23:38])
    
    wire clk_80mhz_enable_134, clk_80mhz_enable_70, n12717, d_clk_tmp, 
        n12691, v_comb, clk_80mhz_enable_11;
    wire [71:0]d_out_11__N_1819;
    wire [15:0]count_15__N_1442;
    
    wire clk_80mhz_enable_155, d_clk_tmp_N_1831;
    wire [71:0]d10;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(54[68:71])
    
    wire n17840, n61, n17839, n16823, n17266, n17231, n17260, 
        n17227, n17846, n17845, n17849, n17848, n17852, n17851, 
        n17855, n17854, clk_80mhz_enable_205, clk_80mhz_enable_255, 
        clk_80mhz_enable_305, clk_80mhz_enable_355, clk_80mhz_enable_405, 
        clk_80mhz_enable_455, clk_80mhz_enable_505, clk_80mhz_enable_555, 
        clk_80mhz_enable_605, clk_80mhz_enable_655, clk_80mhz_enable_705;
    wire [71:0]d10_71__N_1747;
    
    wire clk_80mhz_enable_706, clk_80mhz_enable_707, clk_80mhz_enable_708, 
        clk_80mhz_enable_709, clk_80mhz_enable_710, clk_80mhz_enable_711, 
        clk_80mhz_enable_712, clk_80mhz_enable_713, clk_80mhz_enable_714, 
        clk_80mhz_enable_715, clk_80mhz_enable_716, n17861, n17314, 
        n17860, n17864, n17863, n17867, n17866, n17870, n17869, 
        n17873, n17872, n17147, n63_adj_2568, n131, n64, n132, 
        n65_c, n133, n66_adj_2569, n134, n135, n136, n131_adj_2574, 
        n132_adj_2581, n133_adj_2584, n134_adj_2588, n135_adj_2591, 
        n136_adj_2599, n31_adj_2627, n18066, n17163, n17167, n17165;
    
    LUT4 sub_27_inv_0_i59_1_lut (.A(d_d7[58]), .Z(n15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i59_1_lut.init = 16'h5555;
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_490[20]), .CK(clk_80mhz), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i20.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i61_1_lut (.A(d_d_tmp[60]), .Z(n13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i62_1_lut (.A(d_d_tmp[61]), .Z(n12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i60_1_lut (.A(d_d7[59]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i60_1_lut.init = 16'h5555;
    FD1S3AX d2_i0 (.D(d2_71__N_490[0]), .CK(clk_80mhz), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i0.GSR = "ENABLED";
    FD1S3AX d3_i0 (.D(d3_71__N_562[0]), .CK(clk_80mhz), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(n87_adj_114[1]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i1.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_634[0]), .CK(clk_80mhz), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_706[0]), .CK(clk_80mhz), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1459[0]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    FD1S3JX d_clk_tmp_65 (.D(n12691), .CK(clk_80mhz), .PD(clk_80mhz_enable_134), 
            .Q(d_clk_tmp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_clk_tmp_65.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1S3AX d_clk_67 (.D(d_clk_tmp), .CK(clk_80mhz), .Q(CIC1_out_clkSin)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_clk_67.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_490[19]), .CK(clk_80mhz), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_490[18]), .CK(clk_80mhz), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1531[0]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1603[0]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1675[0]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i57_1_lut (.A(d_d7[56]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i57_1_lut.init = 16'h5555;
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1819[0]), .SP(clk_80mhz_enable_11), 
            .CK(clk_80mhz), .Q(MultDataB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_418[0]), .CK(clk_80mhz), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i0.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_490[17]), .CK(clk_80mhz), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_490[16]), .CK(clk_80mhz), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_15__N_1442[0]), .CK(clk_80mhz), .CD(clk_80mhz_enable_134), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i0.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_490[15]), .CK(clk_80mhz), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i15.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i58_1_lut (.A(d_d7[57]), .Z(n16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i58_1_lut.init = 16'h5555;
    FD1S3AX d2_i14 (.D(d2_71__N_490[14]), .CK(clk_80mhz), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i14.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i59_1_lut (.A(d_d_tmp[58]), .Z(n15_adj_1)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i55_1_lut (.A(d_d7[54]), .Z(n19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i55_1_lut.init = 16'h5555;
    FD1S3AX d2_i13 (.D(d2_71__N_490[13]), .CK(clk_80mhz), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i13.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i60_1_lut (.A(d_d_tmp[59]), .Z(n14_adj_2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i57_1_lut (.A(d_d_tmp[56]), .Z(n17_adj_3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i57_1_lut.init = 16'h5555;
    FD1S3AX d2_i12 (.D(d2_71__N_490[12]), .CK(clk_80mhz), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i12.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i58_1_lut (.A(d_d_tmp[57]), .Z(n16_adj_4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i56_1_lut (.A(d_d7[55]), .Z(n18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i55_1_lut (.A(d_d_tmp[54]), .Z(n19_adj_5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i53_1_lut (.A(d_d7[52]), .Z(n21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i54_1_lut (.A(d_d7[53]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i56_1_lut (.A(d_d_tmp[55]), .Z(n18_adj_6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i51_1_lut (.A(d_d7[50]), .Z(n23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i51_1_lut.init = 16'h5555;
    FD1S3AX d2_i11 (.D(d2_71__N_490[11]), .CK(clk_80mhz), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i11.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i52_1_lut (.A(d_d7[51]), .Z(n22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i52_1_lut.init = 16'h5555;
    FD1S3AX d2_i10 (.D(d2_71__N_490[10]), .CK(clk_80mhz), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i10.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i53_1_lut (.A(d_d_tmp[52]), .Z(n21_adj_7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i49_1_lut (.A(d_d7[48]), .Z(n25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i49_1_lut.init = 16'h5555;
    FD1S3AX d2_i9 (.D(d2_71__N_490[9]), .CK(clk_80mhz), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i9.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i50_1_lut (.A(d_d7[49]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i47_1_lut (.A(d_d7[46]), .Z(n27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i54_1_lut (.A(d_d_tmp[53]), .Z(n20_adj_8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i51_1_lut (.A(d_d_tmp[50]), .Z(n23_adj_9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i52_1_lut (.A(d_d_tmp[51]), .Z(n22_adj_10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i48_1_lut (.A(d_d7[47]), .Z(n26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i45_1_lut (.A(d_d7[44]), .Z(n29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i45_1_lut.init = 16'h5555;
    FD1S3AX d2_i8 (.D(d2_71__N_490[8]), .CK(clk_80mhz), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_490[7]), .CK(clk_80mhz), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_490[6]), .CK(clk_80mhz), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i6.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i49_1_lut (.A(d_d_tmp[48]), .Z(n25_adj_11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i49_1_lut.init = 16'h5555;
    FD1S3AX d2_i5 (.D(d2_71__N_490[5]), .CK(clk_80mhz), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_490[4]), .CK(clk_80mhz), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_490[3]), .CK(clk_80mhz), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i2 (.D(d2_71__N_490[2]), .CK(clk_80mhz), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i1 (.D(d2_71__N_490[1]), .CK(clk_80mhz), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i1.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i46_1_lut (.A(d_d7[45]), .Z(n28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i46_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i50_1_lut (.A(d_d_tmp[49]), .Z(n24_adj_12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i47_1_lut (.A(d_d_tmp[46]), .Z(n27_adj_13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i48_1_lut (.A(d_d_tmp[47]), .Z(n26_adj_14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i48_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i43_1_lut (.A(d_d7[42]), .Z(n31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i43_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i45_1_lut (.A(d_d_tmp[44]), .Z(n29_adj_15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i46_1_lut (.A(d_d_tmp[45]), .Z(n28_adj_16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i43_1_lut (.A(d_d_tmp[42]), .Z(n31_adj_17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i43_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i44_1_lut (.A(d_d_tmp[43]), .Z(n30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i44_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i44_1_lut (.A(d_d7[43]), .Z(n30_adj_18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i44_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(clk_80mhz_enable_70), .CK(clk_80mhz), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i41_1_lut (.A(d_d7[40]), .Z(n33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i41_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i42_1_lut (.A(d_d7[41]), .Z(n32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i41_1_lut (.A(d_d_tmp[40]), .Z(n33_adj_19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i41_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i42_1_lut (.A(d_d_tmp[41]), .Z(n32_adj_20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i42_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i39_1_lut (.A(d_d_tmp[38]), .Z(n35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i39_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i40_1_lut (.A(d_d_tmp[39]), .Z(n34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i39_1_lut (.A(d_d7[38]), .Z(n35_adj_21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i39_1_lut.init = 16'h5555;
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i37_1_lut (.A(d_d_tmp[36]), .Z(n37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i37_1_lut.init = 16'h5555;
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i38_1_lut (.A(d_d_tmp[37]), .Z(n36_adj_22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i38_1_lut.init = 16'h5555;
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i40_1_lut (.A(d_d7[39]), .Z(n34_adj_23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i40_1_lut.init = 16'h5555;
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i37_1_lut (.A(d_d7[36]), .Z(n37_adj_24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i37_1_lut.init = 16'h5555;
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i38_1_lut (.A(d_d7[37]), .Z(n36_adj_25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i38_1_lut.init = 16'h5555;
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    LUT4 i6057_then_3_lut (.A(\CICGain[1] ), .B(d10[59]), .C(d10[57]), 
         .Z(n17840)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6057_then_3_lut.init = 16'he4e4;
    LUT4 i6057_else_3_lut (.A(n61), .B(\CICGain[1] ), .C(d10[58]), .Z(n17839)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6057_else_3_lut.init = 16'he2e2;
    FD1S3AX d2_i21 (.D(d2_71__N_490[21]), .CK(clk_80mhz), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i21.GSR = "ENABLED";
    LUT4 i5959_4_lut (.A(n16823), .B(n17266), .C(n17231), .D(count[7]), 
         .Z(d_clk_tmp_N_1831)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(69[13:41])
    defparam i5959_4_lut.init = 16'h4000;
    LUT4 i5879_4_lut (.A(count[0]), .B(n17260), .C(n17227), .D(count[5]), 
         .Z(n17266)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5879_4_lut.init = 16'h8000;
    LUT4 shift_right_31_i210_3_lut_4_lut_then_3_lut (.A(\CICGain[0] ), .B(\d10[66] ), 
         .C(\d10[67] ), .Z(n17846)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 i1_2_lut (.A(count[10]), .B(count[9]), .Z(n17231)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 shift_right_31_i210_3_lut_4_lut_else_3_lut (.A(\CICGain[0] ), .B(\d10[69] ), 
         .C(\d10[68] ), .Z(n17845)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_else_3_lut.init = 16'he4e4;
    LUT4 sub_26_inv_0_i71_1_lut (.A(d_d6[70]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i72_1_lut (.A(d_d6[71]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i209_3_lut_4_lut_then_3_lut (.A(\CICGain[0] ), .B(\d10[65] ), 
         .C(\d10[66] ), .Z(n17849)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam shift_right_31_i209_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 shift_right_31_i209_3_lut_4_lut_else_3_lut (.A(\CICGain[0] ), .B(\d10[68] ), 
         .C(\d10[67] ), .Z(n17848)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam shift_right_31_i209_3_lut_4_lut_else_3_lut.init = 16'he4e4;
    LUT4 shift_right_31_i210_3_lut_4_lut_then_3_lut_adj_25 (.A(\CICGain[0] ), 
         .B(d10[66]), .C(d10[67]), .Z(n17852)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_then_3_lut_adj_25.init = 16'hd8d8;
    LUT4 shift_right_31_i210_3_lut_4_lut_else_3_lut_adj_26 (.A(\CICGain[0] ), 
         .B(d10[69]), .C(d10[68]), .Z(n17851)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_else_3_lut_adj_26.init = 16'he4e4;
    LUT4 shift_right_31_i209_3_lut_4_lut_then_3_lut_adj_27 (.A(\CICGain[0] ), 
         .B(d10[65]), .C(d10[66]), .Z(n17855)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam shift_right_31_i209_3_lut_4_lut_then_3_lut_adj_27.init = 16'hd8d8;
    LUT4 shift_right_31_i209_3_lut_4_lut_else_3_lut_adj_28 (.A(\CICGain[0] ), 
         .B(d10[68]), .C(d10[67]), .Z(n17854)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam shift_right_31_i209_3_lut_4_lut_else_3_lut_adj_28.init = 16'he4e4;
    FD1S3AX d2_i22 (.D(d2_71__N_490[22]), .CK(clk_80mhz), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_490[23]), .CK(clk_80mhz), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_490[24]), .CK(clk_80mhz), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_490[25]), .CK(clk_80mhz), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_490[26]), .CK(clk_80mhz), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_490[27]), .CK(clk_80mhz), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_490[28]), .CK(clk_80mhz), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_490[29]), .CK(clk_80mhz), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_490[30]), .CK(clk_80mhz), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_490[31]), .CK(clk_80mhz), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_490[32]), .CK(clk_80mhz), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_490[33]), .CK(clk_80mhz), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_490[34]), .CK(clk_80mhz), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_490[35]), .CK(clk_80mhz), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_490[36]), .CK(clk_80mhz), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_490[37]), .CK(clk_80mhz), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_490[38]), .CK(clk_80mhz), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_490[39]), .CK(clk_80mhz), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_490[40]), .CK(clk_80mhz), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_490[41]), .CK(clk_80mhz), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_490[42]), .CK(clk_80mhz), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_490[43]), .CK(clk_80mhz), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_490[44]), .CK(clk_80mhz), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_490[45]), .CK(clk_80mhz), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_490[46]), .CK(clk_80mhz), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_490[47]), .CK(clk_80mhz), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_490[48]), .CK(clk_80mhz), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_490[49]), .CK(clk_80mhz), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_490[50]), .CK(clk_80mhz), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_490[51]), .CK(clk_80mhz), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_490[52]), .CK(clk_80mhz), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_490[53]), .CK(clk_80mhz), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_490[54]), .CK(clk_80mhz), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_490[55]), .CK(clk_80mhz), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_490[56]), .CK(clk_80mhz), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_490[57]), .CK(clk_80mhz), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_490[58]), .CK(clk_80mhz), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_490[59]), .CK(clk_80mhz), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_490[60]), .CK(clk_80mhz), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_490[61]), .CK(clk_80mhz), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_490[62]), .CK(clk_80mhz), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_490[63]), .CK(clk_80mhz), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_490[64]), .CK(clk_80mhz), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_490[65]), .CK(clk_80mhz), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_490[66]), .CK(clk_80mhz), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_490[67]), .CK(clk_80mhz), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_490[68]), .CK(clk_80mhz), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_490[69]), .CK(clk_80mhz), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_490[70]), .CK(clk_80mhz), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_490[71]), .CK(clk_80mhz), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_562[1]), .CK(clk_80mhz), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_562[2]), .CK(clk_80mhz), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_562[3]), .CK(clk_80mhz), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_562[4]), .CK(clk_80mhz), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_562[5]), .CK(clk_80mhz), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_562[6]), .CK(clk_80mhz), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_562[7]), .CK(clk_80mhz), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_562[8]), .CK(clk_80mhz), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_562[9]), .CK(clk_80mhz), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_562[10]), .CK(clk_80mhz), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_562[11]), .CK(clk_80mhz), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_562[12]), .CK(clk_80mhz), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_562[13]), .CK(clk_80mhz), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_562[14]), .CK(clk_80mhz), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_562[15]), .CK(clk_80mhz), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_562[16]), .CK(clk_80mhz), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_562[17]), .CK(clk_80mhz), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_562[18]), .CK(clk_80mhz), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_562[19]), .CK(clk_80mhz), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_562[20]), .CK(clk_80mhz), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_562[21]), .CK(clk_80mhz), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_562[22]), .CK(clk_80mhz), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_562[23]), .CK(clk_80mhz), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_562[24]), .CK(clk_80mhz), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_562[25]), .CK(clk_80mhz), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_562[26]), .CK(clk_80mhz), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_562[27]), .CK(clk_80mhz), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_562[28]), .CK(clk_80mhz), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_562[29]), .CK(clk_80mhz), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_562[30]), .CK(clk_80mhz), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_562[31]), .CK(clk_80mhz), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_562[32]), .CK(clk_80mhz), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_562[33]), .CK(clk_80mhz), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_562[34]), .CK(clk_80mhz), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_562[35]), .CK(clk_80mhz), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_562[36]), .CK(clk_80mhz), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_562[37]), .CK(clk_80mhz), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_562[38]), .CK(clk_80mhz), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_562[39]), .CK(clk_80mhz), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_562[40]), .CK(clk_80mhz), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_562[41]), .CK(clk_80mhz), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_562[42]), .CK(clk_80mhz), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_562[43]), .CK(clk_80mhz), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_562[44]), .CK(clk_80mhz), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_562[45]), .CK(clk_80mhz), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_562[46]), .CK(clk_80mhz), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_562[47]), .CK(clk_80mhz), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_562[48]), .CK(clk_80mhz), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_562[49]), .CK(clk_80mhz), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_562[50]), .CK(clk_80mhz), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_562[51]), .CK(clk_80mhz), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_562[52]), .CK(clk_80mhz), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_562[53]), .CK(clk_80mhz), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_562[54]), .CK(clk_80mhz), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_562[55]), .CK(clk_80mhz), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_562[56]), .CK(clk_80mhz), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_562[57]), .CK(clk_80mhz), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_562[58]), .CK(clk_80mhz), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_562[59]), .CK(clk_80mhz), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_562[60]), .CK(clk_80mhz), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_562[61]), .CK(clk_80mhz), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_562[62]), .CK(clk_80mhz), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_562[63]), .CK(clk_80mhz), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_562[64]), .CK(clk_80mhz), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_562[65]), .CK(clk_80mhz), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_562[66]), .CK(clk_80mhz), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_562[67]), .CK(clk_80mhz), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_562[68]), .CK(clk_80mhz), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_562[69]), .CK(clk_80mhz), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_562[70]), .CK(clk_80mhz), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_562[71]), .CK(clk_80mhz), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_634[1]), .CK(clk_80mhz), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_634[2]), .CK(clk_80mhz), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_634[3]), .CK(clk_80mhz), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_634[4]), .CK(clk_80mhz), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_634[5]), .CK(clk_80mhz), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_634[6]), .CK(clk_80mhz), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_634[7]), .CK(clk_80mhz), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_634[8]), .CK(clk_80mhz), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_634[9]), .CK(clk_80mhz), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_634[10]), .CK(clk_80mhz), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_634[11]), .CK(clk_80mhz), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_634[12]), .CK(clk_80mhz), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_634[13]), .CK(clk_80mhz), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_634[14]), .CK(clk_80mhz), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_634[15]), .CK(clk_80mhz), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_634[16]), .CK(clk_80mhz), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_634[17]), .CK(clk_80mhz), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_634[18]), .CK(clk_80mhz), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_634[19]), .CK(clk_80mhz), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_634[20]), .CK(clk_80mhz), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_634[21]), .CK(clk_80mhz), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_634[22]), .CK(clk_80mhz), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_634[23]), .CK(clk_80mhz), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_634[24]), .CK(clk_80mhz), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_634[25]), .CK(clk_80mhz), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_634[26]), .CK(clk_80mhz), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_634[27]), .CK(clk_80mhz), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_634[28]), .CK(clk_80mhz), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_634[29]), .CK(clk_80mhz), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_634[30]), .CK(clk_80mhz), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_634[31]), .CK(clk_80mhz), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_634[32]), .CK(clk_80mhz), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_634[33]), .CK(clk_80mhz), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_634[34]), .CK(clk_80mhz), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_634[35]), .CK(clk_80mhz), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_634[36]), .CK(clk_80mhz), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_634[37]), .CK(clk_80mhz), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_634[38]), .CK(clk_80mhz), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_634[39]), .CK(clk_80mhz), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_634[40]), .CK(clk_80mhz), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_634[41]), .CK(clk_80mhz), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_634[42]), .CK(clk_80mhz), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_634[43]), .CK(clk_80mhz), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_634[44]), .CK(clk_80mhz), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_634[45]), .CK(clk_80mhz), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_634[46]), .CK(clk_80mhz), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_634[47]), .CK(clk_80mhz), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_634[48]), .CK(clk_80mhz), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_634[49]), .CK(clk_80mhz), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_634[50]), .CK(clk_80mhz), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_634[51]), .CK(clk_80mhz), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_634[52]), .CK(clk_80mhz), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_634[53]), .CK(clk_80mhz), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_634[54]), .CK(clk_80mhz), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_634[55]), .CK(clk_80mhz), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_634[56]), .CK(clk_80mhz), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_634[57]), .CK(clk_80mhz), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_634[58]), .CK(clk_80mhz), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_634[59]), .CK(clk_80mhz), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_634[60]), .CK(clk_80mhz), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_634[61]), .CK(clk_80mhz), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_634[62]), .CK(clk_80mhz), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_634[63]), .CK(clk_80mhz), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_634[64]), .CK(clk_80mhz), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_634[65]), .CK(clk_80mhz), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_634[66]), .CK(clk_80mhz), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_634[67]), .CK(clk_80mhz), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_634[68]), .CK(clk_80mhz), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_634[69]), .CK(clk_80mhz), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_634[70]), .CK(clk_80mhz), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_634[71]), .CK(clk_80mhz), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_706[1]), .CK(clk_80mhz), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_706[2]), .CK(clk_80mhz), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_706[3]), .CK(clk_80mhz), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_706[4]), .CK(clk_80mhz), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_706[5]), .CK(clk_80mhz), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_706[6]), .CK(clk_80mhz), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_706[7]), .CK(clk_80mhz), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_706[8]), .CK(clk_80mhz), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_706[9]), .CK(clk_80mhz), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_706[10]), .CK(clk_80mhz), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_706[11]), .CK(clk_80mhz), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_706[12]), .CK(clk_80mhz), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_706[13]), .CK(clk_80mhz), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_706[14]), .CK(clk_80mhz), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_706[15]), .CK(clk_80mhz), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_706[16]), .CK(clk_80mhz), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_706[17]), .CK(clk_80mhz), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_706[18]), .CK(clk_80mhz), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_706[19]), .CK(clk_80mhz), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_706[20]), .CK(clk_80mhz), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_706[21]), .CK(clk_80mhz), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_706[22]), .CK(clk_80mhz), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_706[23]), .CK(clk_80mhz), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_706[24]), .CK(clk_80mhz), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_706[25]), .CK(clk_80mhz), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_706[26]), .CK(clk_80mhz), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_706[27]), .CK(clk_80mhz), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_706[28]), .CK(clk_80mhz), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_706[29]), .CK(clk_80mhz), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_706[30]), .CK(clk_80mhz), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_706[31]), .CK(clk_80mhz), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_706[32]), .CK(clk_80mhz), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_706[33]), .CK(clk_80mhz), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_706[34]), .CK(clk_80mhz), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_706[35]), .CK(clk_80mhz), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_706[36]), .CK(clk_80mhz), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_706[37]), .CK(clk_80mhz), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_706[38]), .CK(clk_80mhz), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_706[39]), .CK(clk_80mhz), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_706[40]), .CK(clk_80mhz), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_706[41]), .CK(clk_80mhz), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_706[42]), .CK(clk_80mhz), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_706[43]), .CK(clk_80mhz), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_706[44]), .CK(clk_80mhz), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_706[45]), .CK(clk_80mhz), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_706[46]), .CK(clk_80mhz), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_706[47]), .CK(clk_80mhz), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_706[48]), .CK(clk_80mhz), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_706[49]), .CK(clk_80mhz), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_706[50]), .CK(clk_80mhz), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_706[51]), .CK(clk_80mhz), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_706[52]), .CK(clk_80mhz), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_706[53]), .CK(clk_80mhz), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_706[54]), .CK(clk_80mhz), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_706[55]), .CK(clk_80mhz), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_706[56]), .CK(clk_80mhz), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_706[57]), .CK(clk_80mhz), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_706[58]), .CK(clk_80mhz), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_706[59]), .CK(clk_80mhz), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_706[60]), .CK(clk_80mhz), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_706[61]), .CK(clk_80mhz), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_706[62]), .CK(clk_80mhz), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_706[63]), .CK(clk_80mhz), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_706[64]), .CK(clk_80mhz), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_706[65]), .CK(clk_80mhz), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_706[66]), .CK(clk_80mhz), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_706[67]), .CK(clk_80mhz), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_706[68]), .CK(clk_80mhz), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_706[69]), .CK(clk_80mhz), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_706[70]), .CK(clk_80mhz), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_706[71]), .CK(clk_80mhz), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1459[1]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1459[2]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1459[3]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1459[4]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1459[5]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1459[6]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1459[7]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1459[8]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1459[9]), .SP(clk_80mhz_enable_155), .CK(clk_80mhz), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1459[10]), .SP(clk_80mhz_enable_155), 
            .CK(clk_80mhz), .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1459[11]), .SP(clk_80mhz_enable_155), 
            .CK(clk_80mhz), .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1459[12]), .SP(clk_80mhz_enable_155), 
            .CK(clk_80mhz), .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1459[13]), .SP(clk_80mhz_enable_155), 
            .CK(clk_80mhz), .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1459[14]), .SP(clk_80mhz_enable_155), 
            .CK(clk_80mhz), .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1459[15]), .SP(clk_80mhz_enable_155), 
            .CK(clk_80mhz), .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1459[16]), .SP(clk_80mhz_enable_155), 
            .CK(clk_80mhz), .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1459[17]), .SP(clk_80mhz_enable_155), 
            .CK(clk_80mhz), .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1459[18]), .SP(clk_80mhz_enable_155), 
            .CK(clk_80mhz), .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1459[19]), .SP(clk_80mhz_enable_155), 
            .CK(clk_80mhz), .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1459[20]), .SP(clk_80mhz_enable_155), 
            .CK(clk_80mhz), .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1459[21]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1459[22]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1459[23]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1459[24]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1459[25]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1459[26]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1459[27]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1459[28]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1459[29]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1459[30]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1459[31]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1459[32]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1459[33]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1459[34]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1459[35]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1459[36]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1459[37]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1459[38]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1459[39]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1459[40]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1459[41]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1459[42]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1459[43]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1459[44]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1459[45]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1459[46]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1459[47]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1459[48]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1459[49]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1459[50]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1459[51]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1459[52]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1459[53]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1459[54]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1459[55]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1459[56]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1459[57]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1459[58]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1459[59]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1459[60]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1459[61]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1459[62]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1459[63]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1459[64]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1459[65]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1459[66]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1459[67]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1459[68]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1459[69]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1459[70]), .SP(clk_80mhz_enable_205), 
            .CK(clk_80mhz), .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1459[71]), .SP(clk_80mhz_enable_255), 
            .CK(clk_80mhz), .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(clk_80mhz_enable_255), .CK(clk_80mhz), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1531[1]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1531[2]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1531[3]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1531[4]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1531[5]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1531[6]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1531[7]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1531[8]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1531[9]), .SP(clk_80mhz_enable_305), .CK(clk_80mhz), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1531[10]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1531[11]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1531[12]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1531[13]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1531[14]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1531[15]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1531[16]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1531[17]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1531[18]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1531[19]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1531[20]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1531[21]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1531[22]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1531[23]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1531[24]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1531[25]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1531[26]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1531[27]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1531[28]), .SP(clk_80mhz_enable_305), 
            .CK(clk_80mhz), .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1531[29]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1531[30]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1531[31]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1531[32]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1531[33]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1531[34]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1531[35]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1531[36]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1531[37]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1531[38]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1531[39]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1531[40]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1531[41]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1531[42]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1531[43]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1531[44]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1531[45]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1531[46]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1531[47]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1531[48]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1531[49]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1531[50]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1531[51]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1531[52]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1531[53]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1531[54]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1531[55]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1531[56]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1531[57]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1531[58]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1531[59]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1531[60]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1531[61]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1531[62]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1531[63]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1531[64]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1531[65]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1531[66]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1531[67]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1531[68]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1531[69]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1531[70]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1531[71]), .SP(clk_80mhz_enable_355), 
            .CK(clk_80mhz), .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(clk_80mhz_enable_355), .CK(clk_80mhz), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(clk_80mhz_enable_355), .CK(clk_80mhz), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(clk_80mhz_enable_355), .CK(clk_80mhz), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(clk_80mhz_enable_355), .CK(clk_80mhz), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(clk_80mhz_enable_355), .CK(clk_80mhz), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(clk_80mhz_enable_355), .CK(clk_80mhz), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(clk_80mhz_enable_355), .CK(clk_80mhz), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(clk_80mhz_enable_405), .CK(clk_80mhz), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1603[1]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1603[2]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1603[3]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1603[4]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1603[5]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1603[6]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1603[7]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1603[8]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1603[9]), .SP(clk_80mhz_enable_455), .CK(clk_80mhz), 
            .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1603[10]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1603[11]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1603[12]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1603[13]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1603[14]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1603[15]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1603[16]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1603[17]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1603[18]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1603[19]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1603[20]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1603[21]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1603[22]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1603[23]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1603[24]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1603[25]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1603[26]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1603[27]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1603[28]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1603[29]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1603[30]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1603[31]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1603[32]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1603[33]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1603[34]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1603[35]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1603[36]), .SP(clk_80mhz_enable_455), 
            .CK(clk_80mhz), .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1603[37]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1603[38]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1603[39]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1603[40]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1603[41]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1603[42]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1603[43]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1603[44]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1603[45]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1603[46]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1603[47]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1603[48]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1603[49]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1603[50]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1603[51]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1603[52]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1603[53]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1603[54]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1603[55]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1603[56]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1603[57]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1603[58]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1603[59]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1603[60]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1603[61]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1603[62]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1603[63]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1603[64]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1603[65]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1603[66]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1603[67]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1603[68]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1603[69]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1603[70]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1603[71]), .SP(clk_80mhz_enable_505), 
            .CK(clk_80mhz), .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(clk_80mhz_enable_505), .CK(clk_80mhz), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(clk_80mhz_enable_555), .CK(clk_80mhz), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1675[1]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1675[2]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1675[3]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1675[4]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1675[5]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1675[6]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1675[7]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1675[8]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1675[9]), .SP(clk_80mhz_enable_605), .CK(clk_80mhz), 
            .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1675[10]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1675[11]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1675[12]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1675[13]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1675[14]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1675[15]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1675[16]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1675[17]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1675[18]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1675[19]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1675[20]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1675[21]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1675[22]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1675[23]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1675[24]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1675[25]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1675[26]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1675[27]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1675[28]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1675[29]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1675[30]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1675[31]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1675[32]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1675[33]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1675[34]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1675[35]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1675[36]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1675[37]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1675[38]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1675[39]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1675[40]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1675[41]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1675[42]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1675[43]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1675[44]), .SP(clk_80mhz_enable_605), 
            .CK(clk_80mhz), .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1675[45]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1675[46]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1675[47]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1675[48]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1675[49]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1675[50]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1675[51]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1675[52]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1675[53]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1675[54]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1675[55]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1675[56]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1675[57]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1675[58]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1675[59]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1675[60]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1675[61]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1675[62]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1675[63]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1675[64]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1675[65]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1675[66]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1675[67]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1675[68]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1675[69]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1675[70]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1675[71]), .SP(clk_80mhz_enable_655), 
            .CK(clk_80mhz), .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(clk_80mhz_enable_655), .CK(clk_80mhz), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(clk_80mhz_enable_705), .CK(clk_80mhz), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1747[57]), .SP(clk_80mhz_enable_705), 
            .CK(clk_80mhz), .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1747[58]), .SP(clk_80mhz_enable_705), 
            .CK(clk_80mhz), .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1747[59]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1747[60]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1747[61]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1747[62]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1747[63]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1747[64]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1747[65]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1747[66]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1747[67]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1747[68]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1747[69]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1747[70]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1747[71]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1819[1]), .SP(clk_80mhz_enable_706), 
            .CK(clk_80mhz), .Q(MultDataB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(d_out_11__N_1819[2]), .SP(clk_80mhz_enable_707), 
            .CK(clk_80mhz), .Q(MultDataB[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(d_out_11__N_1819[3]), .SP(clk_80mhz_enable_708), 
            .CK(clk_80mhz), .Q(MultDataB[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(d_out_11__N_1819[4]), .SP(clk_80mhz_enable_709), 
            .CK(clk_80mhz), .Q(MultDataB[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(d_out_11__N_1819[5]), .SP(clk_80mhz_enable_710), 
            .CK(clk_80mhz), .Q(MultDataB[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(d_out_11__N_1819[6]), .SP(clk_80mhz_enable_711), 
            .CK(clk_80mhz), .Q(MultDataB[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(d_out_11__N_1819[7]), .SP(clk_80mhz_enable_712), 
            .CK(clk_80mhz), .Q(MultDataB[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(d_out_11__N_1819[8]), .SP(clk_80mhz_enable_713), 
            .CK(clk_80mhz), .Q(MultDataB[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(d_out_11__N_1819[9]), .SP(clk_80mhz_enable_714), 
            .CK(clk_80mhz), .Q(MultDataB[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(d_out_11__N_1819[10]), .SP(clk_80mhz_enable_715), 
            .CK(clk_80mhz), .Q(MultDataB[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(d_out_11__N_1819[11]), .SP(clk_80mhz_enable_716), 
            .CK(clk_80mhz), .Q(MultDataB[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_418[1]), .CK(clk_80mhz), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_418[2]), .CK(clk_80mhz), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_418[3]), .CK(clk_80mhz), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_418[4]), .CK(clk_80mhz), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_418[5]), .CK(clk_80mhz), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_418[6]), .CK(clk_80mhz), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_418[7]), .CK(clk_80mhz), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_418[8]), .CK(clk_80mhz), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_418[9]), .CK(clk_80mhz), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_418[10]), .CK(clk_80mhz), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_418[11]), .CK(clk_80mhz), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_418[12]), .CK(clk_80mhz), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_418[13]), .CK(clk_80mhz), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_418[14]), .CK(clk_80mhz), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_418[15]), .CK(clk_80mhz), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_418[16]), .CK(clk_80mhz), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_418[17]), .CK(clk_80mhz), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_418[18]), .CK(clk_80mhz), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_418[19]), .CK(clk_80mhz), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_418[20]), .CK(clk_80mhz), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_418[21]), .CK(clk_80mhz), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_418[22]), .CK(clk_80mhz), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_418[23]), .CK(clk_80mhz), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_418[24]), .CK(clk_80mhz), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_418[25]), .CK(clk_80mhz), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_418[26]), .CK(clk_80mhz), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_418[27]), .CK(clk_80mhz), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_418[28]), .CK(clk_80mhz), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_418[29]), .CK(clk_80mhz), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_418[30]), .CK(clk_80mhz), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_418[31]), .CK(clk_80mhz), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_418[32]), .CK(clk_80mhz), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_418[33]), .CK(clk_80mhz), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_418[34]), .CK(clk_80mhz), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_418[35]), .CK(clk_80mhz), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_418[36]), .CK(clk_80mhz), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_418[37]), .CK(clk_80mhz), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_418[38]), .CK(clk_80mhz), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_418[39]), .CK(clk_80mhz), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_418[40]), .CK(clk_80mhz), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_418[41]), .CK(clk_80mhz), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_418[42]), .CK(clk_80mhz), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_418[43]), .CK(clk_80mhz), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_418[44]), .CK(clk_80mhz), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_418[45]), .CK(clk_80mhz), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_418[46]), .CK(clk_80mhz), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_418[47]), .CK(clk_80mhz), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_418[48]), .CK(clk_80mhz), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_418[49]), .CK(clk_80mhz), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_418[50]), .CK(clk_80mhz), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_418[51]), .CK(clk_80mhz), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_418[52]), .CK(clk_80mhz), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_418[53]), .CK(clk_80mhz), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_418[54]), .CK(clk_80mhz), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_418[55]), .CK(clk_80mhz), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_418[56]), .CK(clk_80mhz), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_418[57]), .CK(clk_80mhz), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_418[58]), .CK(clk_80mhz), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_418[59]), .CK(clk_80mhz), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_418[60]), .CK(clk_80mhz), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_418[61]), .CK(clk_80mhz), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_418[62]), .CK(clk_80mhz), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_418[63]), .CK(clk_80mhz), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_418[64]), .CK(clk_80mhz), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_418[65]), .CK(clk_80mhz), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_418[66]), .CK(clk_80mhz), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_418[67]), .CK(clk_80mhz), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_418[68]), .CK(clk_80mhz), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_418[69]), .CK(clk_80mhz), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_418[70]), .CK(clk_80mhz), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_418[71]), .CK(clk_80mhz), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i71.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(n87_adj_114[2]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n87_adj_114[3]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n87_adj_114[4]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n87_adj_114[5]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n87_adj_114[6]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n87_adj_114[7]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n87_adj_114[8]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n87_adj_114[9]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n87_adj_114[10]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1442[11]), .CK(clk_80mhz), .CD(d_clk_tmp_N_1831), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n87_adj_114[12]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n87_adj_114[13]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n87_adj_114[14]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n87_adj_114[15]), .CK(clk_80mhz), .CD(n12717), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i15.GSR = "ENABLED";
    LUT4 i5873_4_lut (.A(count[2]), .B(count[8]), .C(count[3]), .D(count[1]), 
         .Z(n17260)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i5873_4_lut.init = 16'h8000;
    LUT4 sub_26_inv_0_i69_1_lut (.A(d_d6[68]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 i6077_then_3_lut (.A(\CICGain[1] ), .B(d10[60]), .C(d10[58]), 
         .Z(n17861)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6077_then_3_lut.init = 16'he4e4;
    LUT4 i6077_else_3_lut (.A(n17314), .B(\CICGain[1] ), .C(d10[59]), 
         .Z(n17860)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6077_else_3_lut.init = 16'he2e2;
    LUT4 shift_right_31_i212_3_lut_4_lut_then_3_lut (.A(\CICGain[1] ), .B(\d10[68] ), 
         .C(\d10[70] ), .Z(n17864)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i212_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 sub_26_inv_0_i70_1_lut (.A(d_d6[69]), .Z(n4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i212_3_lut_4_lut_else_3_lut (.A(\d10[71] ), .B(\CICGain[1] ), 
         .C(\d10[69] ), .Z(n17863)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i212_3_lut_4_lut_else_3_lut.init = 16'he2e2;
    LUT4 i11_3_lut_4_lut_then_3_lut (.A(\CICGain[1] ), .B(\d10[67] ), .C(\d10[69] ), 
         .Z(n17867)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam i11_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 sub_26_inv_0_i67_1_lut (.A(d_d6[66]), .Z(n7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i68_1_lut (.A(d_d6[67]), .Z(n6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 i11_3_lut_4_lut_else_3_lut (.A(\d10[70] ), .B(\CICGain[1] ), .C(\d10[68] ), 
         .Z(n17866)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam i11_3_lut_4_lut_else_3_lut.init = 16'he2e2;
    LUT4 shift_right_31_i212_3_lut_4_lut_then_3_lut_adj_29 (.A(\CICGain[1] ), 
         .B(d10[68]), .C(d10[70]), .Z(n17870)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i212_3_lut_4_lut_then_3_lut_adj_29.init = 16'hd8d8;
    LUT4 i1_2_lut_adj_30 (.A(count[6]), .B(count[4]), .Z(n17227)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_30.init = 16'h8888;
    LUT4 shift_right_31_i212_3_lut_4_lut_else_3_lut_adj_31 (.A(d10[71]), .B(\CICGain[1] ), 
         .C(d10[69]), .Z(n17869)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i212_3_lut_4_lut_else_3_lut_adj_31.init = 16'he2e2;
    LUT4 sub_26_inv_0_i65_1_lut (.A(d_d6[64]), .Z(n9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i66_1_lut (.A(d_d6[65]), .Z(n8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 i11_3_lut_4_lut_then_3_lut_adj_32 (.A(\CICGain[1] ), .B(d10[67]), 
         .C(d10[69]), .Z(n17873)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam i11_3_lut_4_lut_then_3_lut_adj_32.init = 16'hd8d8;
    LUT4 i11_3_lut_4_lut_else_3_lut_adj_33 (.A(d10[70]), .B(\CICGain[1] ), 
         .C(d10[68]), .Z(n17872)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam i11_3_lut_4_lut_else_3_lut_adj_33.init = 16'he2e2;
    LUT4 i1_4_lut (.A(count[12]), .B(count[11]), .C(n17147), .D(count[15]), 
         .Z(n16823)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 sub_26_inv_0_i63_1_lut (.A(d_d6[62]), .Z(n11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i64_1_lut (.A(d_d6[63]), .Z(n10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i61_1_lut (.A(d_d6[60]), .Z(n13_adj_26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i203_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_adj_2568), .D(n131), .Z(d_out_11__N_1819[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i204_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(n132), .Z(d_out_11__N_1819[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_2_lut_adj_34 (.A(count[14]), .B(count[13]), .Z(n17147)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_34.init = 16'heeee;
    LUT4 shift_right_31_i205_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65_c), .D(n133), .Z(d_out_11__N_1819[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i206_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_adj_2569), .D(n134), .Z(d_out_11__N_1819[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i207_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(d10[66]), .D(n135), .Z(d_out_11__N_1819[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i208_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(d10[67]), .D(n136), .Z(d_out_11__N_1819[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1201_i2_3_lut (.A(n118), .B(n120), .C(cout), .Z(d10_71__N_1747[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1201_i3_3_lut (.A(n115), .B(n117), .C(cout), .Z(d10_71__N_1747[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1201_i4_3_lut (.A(n112), .B(n114), .C(cout), .Z(d10_71__N_1747[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i4_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i71_1_lut (.A(d_d8[70]), .Z(n3_adj_27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 mux_1201_i5_3_lut (.A(n109), .B(n111), .C(cout), .Z(d10_71__N_1747[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i5_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i72_1_lut (.A(d_d8[71]), .Z(n2_adj_28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i69_1_lut (.A(d_d8[68]), .Z(n5_adj_29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i203_3_lut_4_lut_adj_35 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_adj_30), .D(n131_adj_2574), .Z(\d_out_11__N_1819[2] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut_adj_35.init = 16'hfe10;
    LUT4 sub_28_inv_0_i70_1_lut (.A(d_d8[69]), .Z(n4_adj_31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i62_1_lut (.A(d_d6[61]), .Z(n12_adj_32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i67_1_lut (.A(d_d8[66]), .Z(n7_adj_33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i68_1_lut (.A(d_d8[67]), .Z(n6_adj_34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i65_1_lut (.A(d_d8[64]), .Z(n9_adj_35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i204_3_lut_4_lut_adj_36 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17288), .D(n132_adj_2581), .Z(\d_out_11__N_1819[3] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut_adj_36.init = 16'hfe10;
    LUT4 shift_right_31_i205_3_lut_4_lut_adj_37 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(n133_adj_2584), .Z(\d_out_11__N_1819[4] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut_adj_37.init = 16'hfe10;
    LUT4 sub_28_inv_0_i66_1_lut (.A(d_d8[65]), .Z(n8_adj_36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i206_3_lut_4_lut_adj_38 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_adj_37), .D(n134_adj_2588), .Z(\d_out_11__N_1819[5] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut_adj_38.init = 16'hfe10;
    LUT4 sub_28_inv_0_i63_1_lut (.A(d_d8[62]), .Z(n11_adj_38)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i207_3_lut_4_lut_adj_39 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(\d10[66] ), .D(n135_adj_2591), .Z(\d_out_11__N_1819[6] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut_adj_39.init = 16'hfe10;
    LUT4 sub_28_inv_0_i64_1_lut (.A(d_d8[63]), .Z(n10_adj_39)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i61_1_lut (.A(d_d8[60]), .Z(n13_adj_40)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i62_1_lut (.A(d_d8[61]), .Z(n12_adj_41)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i59_1_lut (.A(d_d6[58]), .Z(n15_adj_42)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i59_1_lut (.A(d_d8[58]), .Z(n15_adj_43)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i60_1_lut (.A(d_d6[59]), .Z(n14_adj_44)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i208_3_lut_4_lut_adj_40 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(\d10[67] ), .D(n136_adj_2599), .Z(\d_out_11__N_1819[7] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut_adj_40.init = 16'hfe10;
    LUT4 sub_28_inv_0_i60_1_lut (.A(d_d8[59]), .Z(n14_adj_45)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i57_1_lut (.A(d_d8[56]), .Z(n17_adj_46)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 mux_1201_i6_3_lut (.A(n106), .B(n108), .C(cout), .Z(d10_71__N_1747[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i6_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i58_1_lut (.A(d_d8[57]), .Z(n16_adj_47)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i57_1_lut (.A(d_d6[56]), .Z(n17_adj_48)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i58_1_lut (.A(d_d6[57]), .Z(n16_adj_49)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i55_1_lut (.A(d_d6[54]), .Z(n19_adj_50)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i56_1_lut (.A(d_d6[55]), .Z(n18_adj_51)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i53_1_lut (.A(d_d6[52]), .Z(n21_adj_52)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i54_1_lut (.A(d_d6[53]), .Z(n20_adj_53)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i51_1_lut (.A(d_d6[50]), .Z(n23_adj_54)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i52_1_lut (.A(d_d6[51]), .Z(n22_adj_55)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i49_1_lut (.A(d_d6[48]), .Z(n25_adj_56)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i50_1_lut (.A(d_d6[49]), .Z(n24_adj_57)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i47_1_lut (.A(d_d6[46]), .Z(n27_adj_58)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i48_1_lut (.A(d_d6[47]), .Z(n26_adj_59)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i45_1_lut (.A(d_d6[44]), .Z(n29_adj_60)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i46_1_lut (.A(d_d6[45]), .Z(n28_adj_61)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i43_1_lut (.A(d_d6[42]), .Z(n31_adj_62)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i44_1_lut (.A(d_d6[43]), .Z(n30_adj_63)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i41_1_lut (.A(d_d6[40]), .Z(n33_adj_64)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i42_1_lut (.A(d_d6[41]), .Z(n32_adj_65)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i39_1_lut (.A(d_d6[38]), .Z(n35_adj_66)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i40_1_lut (.A(d_d6[39]), .Z(n34_adj_67)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i37_1_lut (.A(d_d6[36]), .Z(n37_adj_68)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i38_1_lut (.A(d_d6[37]), .Z(n36_adj_69)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i55_1_lut (.A(d_d8[54]), .Z(n19_adj_70)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 i5961_2_lut (.A(n31_adj_2627), .B(n18066), .Z(n12717)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam i5961_2_lut.init = 16'hdddd;
    LUT4 i3084_2_lut (.A(n87_adj_114[0]), .B(n31_adj_2627), .Z(count_15__N_1442[0])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(78[18] 81[12])
    defparam i3084_2_lut.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_41 (.A(n17163), .B(n16823), .C(n17167), .D(n17165), 
         .Z(n31_adj_2627)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(74[22:52])
    defparam i1_4_lut_adj_41.init = 16'hfffe;
    LUT4 i1_3_lut (.A(count[8]), .B(count[1]), .C(count[9]), .Z(n17163)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(74[22:52])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_42 (.A(count[10]), .B(count[6]), .C(count[7]), .D(count[5]), 
         .Z(n17167)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(74[22:52])
    defparam i1_4_lut_adj_42.init = 16'hfffe;
    LUT4 i1_4_lut_adj_43 (.A(count[2]), .B(count[4]), .C(count[0]), .D(count[3]), 
         .Z(n17165)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(74[22:52])
    defparam i1_4_lut_adj_43.init = 16'hfffe;
    LUT4 sub_28_inv_0_i56_1_lut (.A(d_d8[55]), .Z(n18_adj_71)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 i2781_2_lut (.A(n31_adj_2627), .B(d_clk_tmp), .Z(n12691)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam i2781_2_lut.init = 16'h8888;
    LUT4 sub_28_inv_0_i53_1_lut (.A(d_d8[52]), .Z(n21_adj_72)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i54_1_lut (.A(d_d8[53]), .Z(n20_adj_73)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i54_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_234 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_305)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_234.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i51_1_lut (.A(d_d8[50]), .Z(n23_adj_74)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i52_1_lut (.A(d_d8[51]), .Z(n22_adj_75)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i49_1_lut (.A(d_d8[48]), .Z(n25_adj_76)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i50_1_lut (.A(d_d8[49]), .Z(n24_adj_77)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 i3100_2_lut (.A(n87_adj_114[11]), .B(n31_adj_2627), .Z(count_15__N_1442[11])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(78[18] 81[12])
    defparam i3100_2_lut.init = 16'hbbbb;
    LUT4 sub_28_inv_0_i47_1_lut (.A(d_d8[46]), .Z(n27_adj_78)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i48_1_lut (.A(d_d8[47]), .Z(n26_adj_79)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i45_1_lut (.A(d_d8[44]), .Z(n29_adj_80)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i46_1_lut (.A(d_d8[45]), .Z(n28_adj_81)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i135_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65_c), .D(d10[63]), .Z(n135)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_28_inv_0_i43_1_lut (.A(d_d8[42]), .Z(n31_adj_82)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i44_1_lut (.A(d_d8[43]), .Z(n30_adj_83)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i41_1_lut (.A(d_d8[40]), .Z(n33_adj_84)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i42_1_lut (.A(d_d8[41]), .Z(n32_adj_85)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i39_1_lut (.A(d_d8[38]), .Z(n35_adj_86)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i40_1_lut (.A(d_d8[39]), .Z(n34_adj_87)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i37_1_lut (.A(d_d8[36]), .Z(n37_adj_88)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i38_1_lut (.A(d_d8[37]), .Z(n36_adj_89)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 mux_1201_i7_3_lut (.A(n103), .B(n105), .C(cout), .Z(d10_71__N_1747[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i7_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i71_1_lut (.A(d_d7[70]), .Z(n3_adj_90)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i72_1_lut (.A(d_d7[71]), .Z(n2_adj_91)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 mux_1201_i8_3_lut (.A(n100), .B(n102), .C(cout), .Z(d10_71__N_1747[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1201_i9_3_lut (.A(n97), .B(n99), .C(cout), .Z(d10_71__N_1747[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i9_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i69_1_lut (.A(d_d7[68]), .Z(n5_adj_92)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i70_1_lut (.A(d_d7[69]), .Z(n4_adj_93)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i70_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_233 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_255)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_233.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i67_1_lut (.A(d_d7[66]), .Z(n7_adj_94)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i68_1_lut (.A(d_d7[67]), .Z(n6_adj_95)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i65_1_lut (.A(d_d7[64]), .Z(n9_adj_96)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 mux_1201_i10_3_lut (.A(n94), .B(n96), .C(cout), .Z(d10_71__N_1747[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i10_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i66_1_lut (.A(d_d7[65]), .Z(n8_adj_97)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 mux_1201_i11_3_lut (.A(n91), .B(n93), .C(cout), .Z(d10_71__N_1747[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i11_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i63_1_lut (.A(d_d7[62]), .Z(n11_adj_98)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i63_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_232 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_205)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_232.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i64_1_lut (.A(d_d7[63]), .Z(n10_adj_99)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i61_1_lut (.A(d_d7[60]), .Z(n13_adj_100)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i62_1_lut (.A(d_d7[61]), .Z(n12_adj_101)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 mux_1201_i12_3_lut (.A(n88), .B(n90), .C(cout), .Z(d10_71__N_1747[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i12_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_231 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_155)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_231.GSR = "ENABLED";
    LUT4 mux_1201_i13_3_lut (.A(n85), .B(n87), .C(cout), .Z(d10_71__N_1747[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i13_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_230 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_70)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_230.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_235 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_355)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_235.GSR = "ENABLED";
    LUT4 shift_right_31_i61_3_lut (.A(d10[60]), .B(d10[61]), .C(\CICGain[0] ), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i61_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_226 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_716)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_226.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_236 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_405)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_236.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_237 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_455)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_237.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_238 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_505)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_238.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_242 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_705)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_242.GSR = "ENABLED";
    LUT4 mux_1201_i14_3_lut (.A(n82), .B(n84), .C(cout), .Z(d10_71__N_1747[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i14_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_241 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_655)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_241.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_240 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_605)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_240.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_225 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_715)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_225.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_224 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_714)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_224.GSR = "ENABLED";
    LUT4 mux_1201_i15_3_lut (.A(n79), .B(n81_adj_102), .C(cout), .Z(d10_71__N_1747[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i15_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_239 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_555)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_239.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_223 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_713)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_223.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_222 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_712)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_222.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_221 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_711)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_221.GSR = "ENABLED";
    LUT4 mux_1201_i16_3_lut (.A(n76), .B(n78_adj_103), .C(cout), .Z(d10_71__N_1747[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1201_i16_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_220 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_710)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_220.GSR = "ENABLED";
    LUT4 shift_right_31_i134_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(d10[62]), .Z(n134)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i133_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_adj_2568), .D(d10[61]), .Z(n133)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut.init = 16'hf960;
    FD1S3AX v_comb_66_rep_219 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_709)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_219.GSR = "ENABLED";
    LUT4 shift_right_31_i132_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17314), .D(d10[60]), .Z(n132)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i135_3_lut_4_lut_adj_44 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(\d10[63] ), .Z(n135_adj_2591)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut_adj_44.init = 16'hf960;
    LUT4 shift_right_31_i136_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_adj_37), .D(\d10[64] ), .Z(n136_adj_2599)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i134_3_lut_4_lut_adj_45 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17288), .D(\d10[62] ), .Z(n134_adj_2588)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut_adj_45.init = 16'hf960;
    FD1S3AX v_comb_66_rep_218 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_708)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_218.GSR = "ENABLED";
    LUT4 shift_right_31_i62_rep_45_3_lut (.A(d10[61]), .B(d10[62]), .C(\CICGain[0] ), 
         .Z(n17314)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i62_rep_45_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i132_3_lut_4_lut_adj_46 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17325), .D(\d10[60] ), .Z(n132_adj_2581)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut_adj_46.init = 16'hf960;
    LUT4 shift_right_31_i133_3_lut_4_lut_adj_47 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_adj_30), .D(\d10[61] ), .Z(n133_adj_2584)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut_adj_47.init = 16'hf960;
    LUT4 shift_right_31_i131_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17302), .D(\d10[59] ), .Z(n131_adj_2574)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut.init = 16'hf960;
    FD1S3AX v_comb_66_rep_217 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_707)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_217.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_216 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_706)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_216.GSR = "ENABLED";
    PFUMX i6118 (.BLUT(n17872), .ALUT(n17873), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[10]));
    LUT4 shift_right_31_i136_3_lut_4_lut_adj_48 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_adj_2569), .D(d10[64]), .Z(n136)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut_adj_48.init = 16'hf960;
    FD1S3AX v_comb_66_rep_215 (.D(clk_80mhz_enable_134), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_11)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_215.GSR = "ENABLED";
    LUT4 shift_right_31_i63_3_lut (.A(d10[62]), .B(d10[63]), .C(\CICGain[0] ), 
         .Z(n63_adj_2568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i131_3_lut_4_lut_adj_49 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n61), .D(d10[59]), .Z(n131)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut_adj_49.init = 16'hf960;
    LUT4 shift_right_31_i64_3_lut (.A(d10[63]), .B(d10[64]), .C(\CICGain[0] ), 
         .Z(n64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i65_3_lut (.A(d10[64]), .B(d10[65]), .C(\CICGain[0] ), 
         .Z(n65_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    LUT4 i5959_4_lut_rep_227 (.A(n16823), .B(n17266), .C(n17231), .D(count[7]), 
         .Z(n18066)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(69[13:41])
    defparam i5959_4_lut_rep_227.init = 16'h4000;
    PFUMX i6116 (.BLUT(n17869), .ALUT(n17870), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[11]));
    LUT4 i5959_4_lut_rep_228 (.A(n16823), .B(n17266), .C(n17231), .D(count[7]), 
         .Z(clk_80mhz_enable_134)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(69[13:41])
    defparam i5959_4_lut_rep_228.init = 16'h4000;
    LUT4 shift_right_31_i66_3_lut (.A(d10[65]), .B(d10[66]), .C(\CICGain[0] ), 
         .Z(n66_adj_2569)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    PFUMX i6114 (.BLUT(n17866), .ALUT(n17867), .C0(\CICGain[0] ), .Z(\d_out_11__N_1819[10] ));
    PFUMX i6112 (.BLUT(n17863), .ALUT(n17864), .C0(\CICGain[0] ), .Z(\d_out_11__N_1819[11] ));
    PFUMX i6110 (.BLUT(n17860), .ALUT(n17861), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[1]));
    PFUMX i6106 (.BLUT(n17854), .ALUT(n17855), .C0(\CICGain[1] ), .Z(d_out_11__N_1819[8]));
    PFUMX i6104 (.BLUT(n17851), .ALUT(n17852), .C0(\CICGain[1] ), .Z(d_out_11__N_1819[9]));
    PFUMX i6102 (.BLUT(n17848), .ALUT(n17849), .C0(\CICGain[1] ), .Z(\d_out_11__N_1819[8] ));
    PFUMX i6100 (.BLUT(n17845), .ALUT(n17846), .C0(\CICGain[1] ), .Z(\d_out_11__N_1819[9] ));
    PFUMX i6096 (.BLUT(n17839), .ALUT(n17840), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[0]));
    LUT4 sub_25_inv_0_i71_1_lut (.A(d_d_tmp[70]), .Z(n3_adj_104)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i72_1_lut (.A(d_d_tmp[71]), .Z(n2_adj_105)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i69_1_lut (.A(d_d_tmp[68]), .Z(n5_adj_106)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i70_1_lut (.A(d_d_tmp[69]), .Z(n4_adj_107)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i67_1_lut (.A(d_d_tmp[66]), .Z(n7_adj_108)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i68_1_lut (.A(d_d_tmp[67]), .Z(n6_adj_109)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i65_1_lut (.A(d_d_tmp[64]), .Z(n9_adj_110)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i66_1_lut (.A(d_d_tmp[65]), .Z(n8_adj_111)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i63_1_lut (.A(d_d_tmp[62]), .Z(n11_adj_112)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i64_1_lut (.A(d_d_tmp[63]), .Z(n10_adj_113)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i64_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module AMDemodulator
//

module AMDemodulator (\DataInReg_11__N_1856[0] , CIC1_out_clkSin, CIC1_outCos, 
            MultResult2, \d_out_d_11__N_1874[17] , d_out_d_11__N_1873, 
            MultDataB, MultResult1, VCC_net, GND_net, \DataInReg_11__N_1856[1] , 
            \DataInReg_11__N_1856[2] , \DataInReg_11__N_1856[3] , \DataInReg_11__N_1856[4] , 
            \DataInReg_11__N_1856[5] , \DataInReg_11__N_1856[6] , \DataInReg_11__N_1856[7] , 
            \DataInReg_11__N_1856[8] , \DemodOut[9] , \ISquare[31] , n213, 
            \d_out_d_11__N_1892[17] , \d_out_d_11__N_1890[17] , \d_out_d_11__N_1888[17] , 
            \d_out_d_11__N_1886[17] , \d_out_d_11__N_1884[17] , \d_out_d_11__N_1882[17] , 
            \d_out_d_11__N_1878[17] , d_out_d_11__N_1877, \d_out_d_11__N_1876[17] , 
            d_out_d_11__N_1875, d_out_d_11__N_1879, \d_out_d_11__N_2383[17] , 
            \d_out_d_11__N_2401[17] , \d_out_d_11__N_1880[17] ) /* synthesis syn_module_defined=1 */ ;
    output \DataInReg_11__N_1856[0] ;
    input CIC1_out_clkSin;
    input [11:0]CIC1_outCos;
    output [23:0]MultResult2;
    input \d_out_d_11__N_1874[17] ;
    output d_out_d_11__N_1873;
    input [11:0]MultDataB;
    output [23:0]MultResult1;
    input VCC_net;
    input GND_net;
    output \DataInReg_11__N_1856[1] ;
    output \DataInReg_11__N_1856[2] ;
    output \DataInReg_11__N_1856[3] ;
    output \DataInReg_11__N_1856[4] ;
    output \DataInReg_11__N_1856[5] ;
    output \DataInReg_11__N_1856[6] ;
    output \DataInReg_11__N_1856[7] ;
    output \DataInReg_11__N_1856[8] ;
    output \DemodOut[9] ;
    input \ISquare[31] ;
    output n213;
    input \d_out_d_11__N_1892[17] ;
    input \d_out_d_11__N_1890[17] ;
    input \d_out_d_11__N_1888[17] ;
    input \d_out_d_11__N_1886[17] ;
    input \d_out_d_11__N_1884[17] ;
    input \d_out_d_11__N_1882[17] ;
    input \d_out_d_11__N_1878[17] ;
    output d_out_d_11__N_1877;
    input \d_out_d_11__N_1876[17] ;
    output d_out_d_11__N_1875;
    output d_out_d_11__N_1879;
    input \d_out_d_11__N_2383[17] ;
    input \d_out_d_11__N_2401[17] ;
    input \d_out_d_11__N_1880[17] ;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/top.v(74[23:38])
    wire [15:0]d_out_d;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(30[28:35])
    wire [12:0]n27;
    wire [25:0]n83;
    wire [17:0]d_out_d_11__N_1894;
    
    wire d_out_d_11__N_1891, d_out_d_11__N_1889, d_out_d_11__N_1887, d_out_d_11__N_1885, 
        d_out_d_11__N_1883, d_out_d_11__N_1881;
    
    FD1S3AX d_out_i1 (.D(d_out_d[0]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i1.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i1 (.D(CIC1_outCos[0]), .CK(CIC1_out_clkSin), 
            .Q(n27[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i1.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i0 (.D(n83[0]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i0.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i1 (.D(d_out_d_11__N_1894[17]), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i1.GSR = "ENABLED";
    LUT4 d_out_d_11__I_1_1_lut (.A(\d_out_d_11__N_1874[17] ), .Z(d_out_d_11__N_1873)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_1_1_lut.init = 16'h5555;
    MULT18X18D MultResult1_e3 (.A17(MultDataB[11]), .A16(MultDataB[11]), 
            .A15(MultDataB[11]), .A14(MultDataB[11]), .A13(MultDataB[11]), 
            .A12(MultDataB[11]), .A11(MultDataB[11]), .A10(MultDataB[10]), 
            .A9(MultDataB[9]), .A8(MultDataB[8]), .A7(MultDataB[7]), .A6(MultDataB[6]), 
            .A5(MultDataB[5]), .A4(MultDataB[4]), .A3(MultDataB[3]), .A2(MultDataB[2]), 
            .A1(MultDataB[1]), .A0(MultDataB[0]), .B17(MultDataB[11]), 
            .B16(MultDataB[11]), .B15(MultDataB[11]), .B14(MultDataB[11]), 
            .B13(MultDataB[11]), .B12(MultDataB[11]), .B11(MultDataB[11]), 
            .B10(MultDataB[10]), .B9(MultDataB[9]), .B8(MultDataB[8]), 
            .B7(MultDataB[7]), .B6(MultDataB[6]), .B5(MultDataB[5]), .B4(MultDataB[4]), 
            .B3(MultDataB[3]), .B2(MultDataB[2]), .B1(MultDataB[1]), .B0(MultDataB[0]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(CIC1_out_clkSin), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .P23(MultResult1[23]), 
            .P22(MultResult1[22]), .P21(MultResult1[21]), .P20(MultResult1[20]), 
            .P19(MultResult1[19]), .P18(MultResult1[18]), .P17(MultResult1[17]), 
            .P16(MultResult1[16]), .P15(MultResult1[15]), .P14(MultResult1[14]), 
            .P13(MultResult1[13]), .P12(MultResult1[12]), .P11(MultResult1[11]), 
            .P10(MultResult1[10]), .P9(MultResult1[9]), .P8(MultResult1[8]), 
            .P7(MultResult1[7]), .P6(MultResult1[6]), .P5(MultResult1[5]), 
            .P4(MultResult1[4]), .P3(MultResult1[3]), .P2(MultResult1[2]), 
            .P1(MultResult1[1]), .P0(MultResult1[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(86[20:39])
    defparam MultResult1_e3.REG_INPUTA_CLK = "CLK3";
    defparam MultResult1_e3.REG_INPUTA_CE = "CE3";
    defparam MultResult1_e3.REG_INPUTA_RST = "RST3";
    defparam MultResult1_e3.REG_INPUTB_CLK = "CLK3";
    defparam MultResult1_e3.REG_INPUTB_CE = "CE3";
    defparam MultResult1_e3.REG_INPUTB_RST = "RST3";
    defparam MultResult1_e3.REG_INPUTC_CLK = "NONE";
    defparam MultResult1_e3.REG_INPUTC_CE = "CE0";
    defparam MultResult1_e3.REG_INPUTC_RST = "RST0";
    defparam MultResult1_e3.REG_PIPELINE_CLK = "NONE";
    defparam MultResult1_e3.REG_PIPELINE_CE = "CE0";
    defparam MultResult1_e3.REG_PIPELINE_RST = "RST0";
    defparam MultResult1_e3.REG_OUTPUT_CLK = "CLK3";
    defparam MultResult1_e3.REG_OUTPUT_CE = "CE3";
    defparam MultResult1_e3.REG_OUTPUT_RST = "RST3";
    defparam MultResult1_e3.CLK0_DIV = "ENABLED";
    defparam MultResult1_e3.CLK1_DIV = "ENABLED";
    defparam MultResult1_e3.CLK2_DIV = "ENABLED";
    defparam MultResult1_e3.CLK3_DIV = "ENABLED";
    defparam MultResult1_e3.HIGHSPEED_CLK = "NONE";
    defparam MultResult1_e3.GSR = "ENABLED";
    defparam MultResult1_e3.CAS_MATCH_REG = "FALSE";
    defparam MultResult1_e3.SOURCEB_MODE = "B_SHIFT";
    defparam MultResult1_e3.MULT_BYPASS = "DISABLED";
    defparam MultResult1_e3.RESETMODE = "ASYNC";
    MULT18X18D MultResult2_res2_mult_2 (.A17(n27[12]), .A16(n27[12]), .A15(n27[12]), 
            .A14(n27[12]), .A13(n27[12]), .A12(n27[12]), .A11(n27[12]), 
            .A10(n27[10]), .A9(n27[9]), .A8(n27[8]), .A7(n27[7]), .A6(n27[6]), 
            .A5(n27[5]), .A4(n27[4]), .A3(n27[3]), .A2(n27[2]), .A1(n27[1]), 
            .A0(n27[0]), .B17(n27[12]), .B16(n27[12]), .B15(n27[12]), 
            .B14(n27[12]), .B13(n27[12]), .B12(n27[12]), .B11(n27[12]), 
            .B10(n27[10]), .B9(n27[9]), .B8(n27[8]), .B7(n27[7]), .B6(n27[6]), 
            .B5(n27[5]), .B4(n27[4]), .B3(n27[3]), .B2(n27[2]), .B1(n27[1]), 
            .B0(n27[0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .P23(n83[23]), 
            .P22(n83[22]), .P21(n83[21]), .P20(n83[20]), .P19(n83[19]), 
            .P18(n83[18]), .P17(n83[17]), .P16(n83[16]), .P15(n83[15]), 
            .P14(n83[14]), .P13(n83[13]), .P12(n83[12]), .P11(n83[11]), 
            .P10(n83[10]), .P9(n83[9]), .P8(n83[8]), .P7(n83[7]), .P6(n83[6]), 
            .P5(n83[5]), .P4(n83[4]), .P3(n83[3]), .P2(n83[2]), .P1(n83[1]), 
            .P0(n83[0]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_mult_2.REG_INPUTA_CLK = "NONE";
    defparam MultResult2_res2_mult_2.REG_INPUTA_CE = "CE0";
    defparam MultResult2_res2_mult_2.REG_INPUTA_RST = "RST0";
    defparam MultResult2_res2_mult_2.REG_INPUTB_CLK = "NONE";
    defparam MultResult2_res2_mult_2.REG_INPUTB_CE = "CE0";
    defparam MultResult2_res2_mult_2.REG_INPUTB_RST = "RST0";
    defparam MultResult2_res2_mult_2.REG_INPUTC_CLK = "NONE";
    defparam MultResult2_res2_mult_2.REG_INPUTC_CE = "CE0";
    defparam MultResult2_res2_mult_2.REG_INPUTC_RST = "RST0";
    defparam MultResult2_res2_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam MultResult2_res2_mult_2.REG_PIPELINE_CE = "CE0";
    defparam MultResult2_res2_mult_2.REG_PIPELINE_RST = "RST0";
    defparam MultResult2_res2_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam MultResult2_res2_mult_2.REG_OUTPUT_CE = "CE0";
    defparam MultResult2_res2_mult_2.REG_OUTPUT_RST = "RST0";
    defparam MultResult2_res2_mult_2.CLK0_DIV = "ENABLED";
    defparam MultResult2_res2_mult_2.CLK1_DIV = "ENABLED";
    defparam MultResult2_res2_mult_2.CLK2_DIV = "ENABLED";
    defparam MultResult2_res2_mult_2.CLK3_DIV = "ENABLED";
    defparam MultResult2_res2_mult_2.HIGHSPEED_CLK = "NONE";
    defparam MultResult2_res2_mult_2.GSR = "ENABLED";
    defparam MultResult2_res2_mult_2.CAS_MATCH_REG = "FALSE";
    defparam MultResult2_res2_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam MultResult2_res2_mult_2.MULT_BYPASS = "DISABLED";
    defparam MultResult2_res2_mult_2.RESETMODE = "SYNC";
    FD1S3AX d_out_i2 (.D(d_out_d[1]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i2.GSR = "ENABLED";
    FD1S3AX d_out_i3 (.D(d_out_d[2]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i3.GSR = "ENABLED";
    FD1S3AX d_out_i4 (.D(d_out_d[3]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i4.GSR = "ENABLED";
    FD1S3AX d_out_i5 (.D(d_out_d[4]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i5.GSR = "ENABLED";
    FD1S3AX d_out_i6 (.D(d_out_d[5]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i6.GSR = "ENABLED";
    FD1S3AX d_out_i7 (.D(d_out_d[6]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i7.GSR = "ENABLED";
    FD1S3AX d_out_i8 (.D(d_out_d[7]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i8.GSR = "ENABLED";
    FD1S3AX d_out_i9 (.D(d_out_d[8]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i9.GSR = "ENABLED";
    FD1S3AX d_out_i10 (.D(d_out_d[9]), .CK(CIC1_out_clkSin), .Q(\DemodOut[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i10.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i2 (.D(CIC1_outCos[1]), .CK(CIC1_out_clkSin), 
            .Q(n27[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i2.GSR = "ENABLED";
    LUT4 i1297_1_lut (.A(\ISquare[31] ), .Z(n213)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1297_1_lut.init = 16'h5555;
    FD1S3AX MultResult2_res2_e1__i3 (.D(CIC1_outCos[2]), .CK(CIC1_out_clkSin), 
            .Q(n27[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i3.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i4 (.D(CIC1_outCos[3]), .CK(CIC1_out_clkSin), 
            .Q(n27[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i4.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i5 (.D(CIC1_outCos[4]), .CK(CIC1_out_clkSin), 
            .Q(n27[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i5.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i6 (.D(CIC1_outCos[5]), .CK(CIC1_out_clkSin), 
            .Q(n27[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i6.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i7 (.D(CIC1_outCos[6]), .CK(CIC1_out_clkSin), 
            .Q(n27[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i7.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i8 (.D(CIC1_outCos[7]), .CK(CIC1_out_clkSin), 
            .Q(n27[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i8.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i9 (.D(CIC1_outCos[8]), .CK(CIC1_out_clkSin), 
            .Q(n27[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i9.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i10 (.D(CIC1_outCos[9]), .CK(CIC1_out_clkSin), 
            .Q(n27[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i10.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i11 (.D(CIC1_outCos[10]), .CK(CIC1_out_clkSin), 
            .Q(n27[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i11.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i12 (.D(CIC1_outCos[11]), .CK(CIC1_out_clkSin), 
            .Q(n27[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i12.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i1 (.D(n83[1]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i1.GSR = "ENABLED";
    LUT4 d_out_d_11__I_10_1_lut (.A(\d_out_d_11__N_1892[17] ), .Z(d_out_d_11__N_1891)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_10_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_9_1_lut (.A(\d_out_d_11__N_1890[17] ), .Z(d_out_d_11__N_1889)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_9_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_8_1_lut (.A(\d_out_d_11__N_1888[17] ), .Z(d_out_d_11__N_1887)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_8_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_7_1_lut (.A(\d_out_d_11__N_1886[17] ), .Z(d_out_d_11__N_1885)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_7_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_6_1_lut (.A(\d_out_d_11__N_1884[17] ), .Z(d_out_d_11__N_1883)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_6_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_5_1_lut (.A(\d_out_d_11__N_1882[17] ), .Z(d_out_d_11__N_1881)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_5_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_3_1_lut (.A(\d_out_d_11__N_1878[17] ), .Z(d_out_d_11__N_1877)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_3_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_2_1_lut (.A(\d_out_d_11__N_1876[17] ), .Z(d_out_d_11__N_1875)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_2_1_lut.init = 16'h5555;
    FD1S3AX MultResult2_res2_e3_i0_i2 (.D(n83[2]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i2.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i3 (.D(n83[3]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i3.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i4 (.D(n83[4]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i4.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i5 (.D(n83[5]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i5.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i6 (.D(n83[6]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i6.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i7 (.D(n83[7]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i7.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i8 (.D(n83[8]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i8.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i9 (.D(n83[9]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i9.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i10 (.D(n83[10]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i10.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i11 (.D(n83[11]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i11.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i12 (.D(n83[12]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i12.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i13 (.D(n83[13]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i13.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i14 (.D(n83[14]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i14.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i15 (.D(n83[15]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i15.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i16 (.D(n83[16]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i16.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i17 (.D(n83[17]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i17.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i18 (.D(n83[18]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i18.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i19 (.D(n83[19]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i19.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i20 (.D(n83[20]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i20.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i21 (.D(n83[21]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i21.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i22 (.D(n83[22]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i22.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i23 (.D(n83[23]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i23.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i2 (.D(d_out_d_11__N_1891), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[1]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i2.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i3 (.D(d_out_d_11__N_1889), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[2]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i3.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i4 (.D(d_out_d_11__N_1887), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[3]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i4.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i5 (.D(d_out_d_11__N_1885), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[4]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i5.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i6 (.D(d_out_d_11__N_1883), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[5]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i6.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i7 (.D(d_out_d_11__N_1881), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[6]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i7.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i8 (.D(d_out_d_11__N_1879), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[7]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i8.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i9 (.D(d_out_d_11__N_1877), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[8]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i9.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i10 (.D(d_out_d_11__N_1875), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[9]));   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i10.GSR = "ENABLED";
    LUT4 mux_81_i1_3_lut (.A(\d_out_d_11__N_2383[17] ), .B(\d_out_d_11__N_2401[17] ), 
         .C(\d_out_d_11__N_1892[17] ), .Z(d_out_d_11__N_1894[17])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(70[11:28])
    defparam mux_81_i1_3_lut.init = 16'h3535;
    LUT4 d_out_d_11__I_4_1_lut (.A(\d_out_d_11__N_1880[17] ), .Z(d_out_d_11__N_1879)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/4.lattice/Version1/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_4_1_lut.init = 16'h5555;
    
endmodule
