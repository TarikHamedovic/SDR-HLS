
module quarterwave_table #(
    parameter QLUT_DEPTH = 11,
    parameter DATA_WIDTH = 12
)(
    input  logic        [QLUT_DEPTH-3:0] address, // 9-bit address signal for 512 values
    output logic signed [DATA_WIDTH-1:0] value    // 12-bit output signal
);

    always_comb begin
        unique case(address)
            9'd0: value = 12'h3;
            9'd1: value = 12'h9;
            9'd2: value = 12'hF;
            9'd3: value = 12'h15;
            9'd4: value = 12'h1C;
            9'd5: value = 12'h22;
            9'd6: value = 12'h28;
            9'd7: value = 12'h2F;
            9'd8: value = 12'h35;
            9'd9: value = 12'h3B;
            9'd10: value = 12'h41;
            9'd11: value = 12'h48;
            9'd12: value = 12'h4E;
            9'd13: value = 12'h54;
            9'd14: value = 12'h5B;
            9'd15: value = 12'h61;
            9'd16: value = 12'h67;
            9'd17: value = 12'h6D;
            9'd18: value = 12'h74;
            9'd19: value = 12'h7A;
            9'd20: value = 12'h80;
            9'd21: value = 12'h86;
            9'd22: value = 12'h8D;
            9'd23: value = 12'h93;
            9'd24: value = 12'h99;
            9'd25: value = 12'h9F;
            9'd26: value = 12'hA6;
            9'd27: value = 12'hAC;
            9'd28: value = 12'hB2;
            9'd29: value = 12'hB9;
            9'd30: value = 12'hBF;
            9'd31: value = 12'hC5;
            9'd32: value = 12'hCB;
            9'd33: value = 12'hD2;
            9'd34: value = 12'hD8;
            9'd35: value = 12'hDE;
            9'd36: value = 12'hE4;
            9'd37: value = 12'hEA;
            9'd38: value = 12'hF1;
            9'd39: value = 12'hF7;
            9'd40: value = 12'hFD;
            9'd41: value = 12'h103;
            9'd42: value = 12'h10A;
            9'd43: value = 12'h110;
            9'd44: value = 12'h116;
            9'd45: value = 12'h11C;
            9'd46: value = 12'h123;
            9'd47: value = 12'h129;
            9'd48: value = 12'h12F;
            9'd49: value = 12'h135;
            9'd50: value = 12'h13B;
            9'd51: value = 12'h142;
            9'd52: value = 12'h148;
            9'd53: value = 12'h14E;
            9'd54: value = 12'h154;
            9'd55: value = 12'h15A;
            9'd56: value = 12'h161;
            9'd57: value = 12'h167;
            9'd58: value = 12'h16D;
            9'd59: value = 12'h173;
            9'd60: value = 12'h179;
            9'd61: value = 12'h17F;
            9'd62: value = 12'h186;
            9'd63: value = 12'h18C;
            9'd64: value = 12'h192;
            9'd65: value = 12'h198;
            9'd66: value = 12'h19E;
            9'd67: value = 12'h1A4;
            9'd68: value = 12'h1AB;
            9'd69: value = 12'h1B1;
            9'd70: value = 12'h1B7;
            9'd71: value = 12'h1BD;
            9'd72: value = 12'h1C3;
            9'd73: value = 12'h1C9;
            9'd74: value = 12'h1CF;
            9'd75: value = 12'h1D5;
            9'd76: value = 12'h1DC;
            9'd77: value = 12'h1E2;
            9'd78: value = 12'h1E8;
            9'd79: value = 12'h1EE;
            9'd80: value = 12'h1F4;
            9'd81: value = 12'h1FA;
            9'd82: value = 12'h200;
            9'd83: value = 12'h206;
            9'd84: value = 12'h20C;
            9'd85: value = 12'h212;
            9'd86: value = 12'h218;
            9'd87: value = 12'h21E;
            9'd88: value = 12'h224;
            9'd89: value = 12'h22B;
            9'd90: value = 12'h231;
            9'd91: value = 12'h237;
            9'd92: value = 12'h23D;
            9'd93: value = 12'h243;
            9'd94: value = 12'h249;
            9'd95: value = 12'h24F;
            9'd96: value = 12'h255;
            9'd97: value = 12'h25B;
            9'd98: value = 12'h261;
            9'd99: value = 12'h267;
            9'd100: value = 12'h26D;
            9'd101: value = 12'h273;
            9'd102: value = 12'h279;
            9'd103: value = 12'h27F;
            9'd104: value = 12'h285;
            9'd105: value = 12'h28B;
            9'd106: value = 12'h290;
            9'd107: value = 12'h296;
            9'd108: value = 12'h29C;
            9'd109: value = 12'h2A2;
            9'd110: value = 12'h2A8;
            9'd111: value = 12'h2AE;
            9'd112: value = 12'h2B4;
            9'd113: value = 12'h2BA;
            9'd114: value = 12'h2C0;
            9'd115: value = 12'h2C6;
            9'd116: value = 12'h2CC;
            9'd117: value = 12'h2D2;
            9'd118: value = 12'h2D7;
            9'd119: value = 12'h2DD;
            9'd120: value = 12'h2E3;
            9'd121: value = 12'h2E9;
            9'd122: value = 12'h2EF;
            9'd123: value = 12'h2F5;
            9'd124: value = 12'h2FB;
            9'd125: value = 12'h300;
            9'd126: value = 12'h306;
            9'd127: value = 12'h30C;
            9'd128: value = 12'h312;
            9'd129: value = 12'h318;
            9'd130: value = 12'h31D;
            9'd131: value = 12'h323;
            9'd132: value = 12'h329;
            9'd133: value = 12'h32F;
            9'd134: value = 12'h334;
            9'd135: value = 12'h33A;
            9'd136: value = 12'h340;
            9'd137: value = 12'h346;
            9'd138: value = 12'h34B;
            9'd139: value = 12'h351;
            9'd140: value = 12'h357;
            9'd141: value = 12'h35C;
            9'd142: value = 12'h362;
            9'd143: value = 12'h368;
            9'd144: value = 12'h36E;
            9'd145: value = 12'h373;
            9'd146: value = 12'h379;
            9'd147: value = 12'h37F;
            9'd148: value = 12'h384;
            9'd149: value = 12'h38A;
            9'd150: value = 12'h38F;
            9'd151: value = 12'h395;
            9'd152: value = 12'h39B;
            9'd153: value = 12'h3A0;
            9'd154: value = 12'h3A6;
            9'd155: value = 12'h3AB;
            9'd156: value = 12'h3B1;
            9'd157: value = 12'h3B7;
            9'd158: value = 12'h3BC;
            9'd159: value = 12'h3C2;
            9'd160: value = 12'h3C7;
            9'd161: value = 12'h3CD;
            9'd162: value = 12'h3D2;
            9'd163: value = 12'h3D8;
            9'd164: value = 12'h3DD;
            9'd165: value = 12'h3E3;
            9'd166: value = 12'h3E8;
            9'd167: value = 12'h3EE;
            9'd168: value = 12'h3F3;
            9'd169: value = 12'h3F9;
            9'd170: value = 12'h3FE;
            9'd171: value = 12'h404;
            9'd172: value = 12'h409;
            9'd173: value = 12'h40E;
            9'd174: value = 12'h414;
            9'd175: value = 12'h419;
            9'd176: value = 12'h41F;
            9'd177: value = 12'h424;
            9'd178: value = 12'h429;
            9'd179: value = 12'h42F;
            9'd180: value = 12'h434;
            9'd181: value = 12'h439;
            9'd182: value = 12'h43F;
            9'd183: value = 12'h444;
            9'd184: value = 12'h449;
            9'd185: value = 12'h44F;
            9'd186: value = 12'h454;
            9'd187: value = 12'h459;
            9'd188: value = 12'h45E;
            9'd189: value = 12'h464;
            9'd190: value = 12'h469;
            9'd191: value = 12'h46E;
            9'd192: value = 12'h473;
            9'd193: value = 12'h479;
            9'd194: value = 12'h47E;
            9'd195: value = 12'h483;
            9'd196: value = 12'h488;
            9'd197: value = 12'h48D;
            9'd198: value = 12'h492;
            9'd199: value = 12'h498;
            9'd200: value = 12'h49D;
            9'd201: value = 12'h4A2;
            9'd202: value = 12'h4A7;
            9'd203: value = 12'h4AC;
            9'd204: value = 12'h4B1;
            9'd205: value = 12'h4B6;
            9'd206: value = 12'h4BB;
            9'd207: value = 12'h4C0;
            9'd208: value = 12'h4C5;
            9'd209: value = 12'h4CA;
            9'd210: value = 12'h4CF;
            9'd211: value = 12'h4D4;
            9'd212: value = 12'h4D9;
            9'd213: value = 12'h4DE;
            9'd214: value = 12'h4E3;
            9'd215: value = 12'h4E8;
            9'd216: value = 12'h4ED;
            9'd217: value = 12'h4F2;
            9'd218: value = 12'h4F7;
            9'd219: value = 12'h4FC;
            9'd220: value = 12'h501;
            9'd221: value = 12'h506;
            9'd222: value = 12'h50B;
            9'd223: value = 12'h510;
            9'd224: value = 12'h515;
            9'd225: value = 12'h519;
            9'd226: value = 12'h51E;
            9'd227: value = 12'h523;
            9'd228: value = 12'h528;
            9'd229: value = 12'h52D;
            9'd230: value = 12'h531;
            9'd231: value = 12'h536;
            9'd232: value = 12'h53B;
            9'd233: value = 12'h540;
            9'd234: value = 12'h544;
            9'd235: value = 12'h549;
            9'd236: value = 12'h54E;
            9'd237: value = 12'h553;
            9'd238: value = 12'h557;
            9'd239: value = 12'h55C;
            9'd240: value = 12'h561;
            9'd241: value = 12'h565;
            9'd242: value = 12'h56A;
            9'd243: value = 12'h56E;
            9'd244: value = 12'h573;
            9'd245: value = 12'h578;
            9'd246: value = 12'h57C;
            9'd247: value = 12'h581;
            9'd248: value = 12'h585;
            9'd249: value = 12'h58A;
            9'd250: value = 12'h58E;
            9'd251: value = 12'h593;
            9'd252: value = 12'h597;
            9'd253: value = 12'h59C;
            9'd254: value = 12'h5A0;
            9'd255: value = 12'h5A5;
            9'd256: value = 12'h5A9;
            9'd257: value = 12'h5AE;
            9'd258: value = 12'h5B2;
            9'd259: value = 12'h5B6;
            9'd260: value = 12'h5BB;
            9'd261: value = 12'h5BF;
            9'd262: value = 12'h5C4;
            9'd263: value = 12'h5C8;
            9'd264: value = 12'h5CC;
            9'd265: value = 12'h5D1;
            9'd266: value = 12'h5D5;
            9'd267: value = 12'h5D9;
            9'd268: value = 12'h5DD;
            9'd269: value = 12'h5E2;
            9'd270: value = 12'h5E6;
            9'd271: value = 12'h5EA;
            9'd272: value = 12'h5EE;
            9'd273: value = 12'h5F3;
            9'd274: value = 12'h5F7;
            9'd275: value = 12'h5FB;
            9'd276: value = 12'h5FF;
            9'd277: value = 12'h603;
            9'd278: value = 12'h607;
            9'd279: value = 12'h60B;
            9'd280: value = 12'h610;
            9'd281: value = 12'h614;
            9'd282: value = 12'h618;
            9'd283: value = 12'h61C;
            9'd284: value = 12'h620;
            9'd285: value = 12'h624;
            9'd286: value = 12'h628;
            9'd287: value = 12'h62C;
            9'd288: value = 12'h630;
            9'd289: value = 12'h634;
            9'd290: value = 12'h638;
            9'd291: value = 12'h63C;
            9'd292: value = 12'h640;
            9'd293: value = 12'h644;
            9'd294: value = 12'h647;
            9'd295: value = 12'h64B;
            9'd296: value = 12'h64F;
            9'd297: value = 12'h653;
            9'd298: value = 12'h657;
            9'd299: value = 12'h65B;
            9'd300: value = 12'h65E;
            9'd301: value = 12'h662;
            9'd302: value = 12'h666;
            9'd303: value = 12'h66A;
            9'd304: value = 12'h66E;
            9'd305: value = 12'h671;
            9'd306: value = 12'h675;
            9'd307: value = 12'h679;
            9'd308: value = 12'h67C;
            9'd309: value = 12'h680;
            9'd310: value = 12'h684;
            9'd311: value = 12'h687;
            9'd312: value = 12'h68B;
            9'd313: value = 12'h68F;
            9'd314: value = 12'h692;
            9'd315: value = 12'h696;
            9'd316: value = 12'h699;
            9'd317: value = 12'h69D;
            9'd318: value = 12'h6A0;
            9'd319: value = 12'h6A4;
            9'd320: value = 12'h6A7;
            9'd321: value = 12'h6AB;
            9'd322: value = 12'h6AE;
            9'd323: value = 12'h6B2;
            9'd324: value = 12'h6B5;
            9'd325: value = 12'h6B8;
            9'd326: value = 12'h6BC;
            9'd327: value = 12'h6BF;
            9'd328: value = 12'h6C3;
            9'd329: value = 12'h6C6;
            9'd330: value = 12'h6C9;
            9'd331: value = 12'h6CD;
            9'd332: value = 12'h6D0;
            9'd333: value = 12'h6D3;
            9'd334: value = 12'h6D6;
            9'd335: value = 12'h6DA;
            9'd336: value = 12'h6DD;
            9'd337: value = 12'h6E0;
            9'd338: value = 12'h6E3;
            9'd339: value = 12'h6E6;
            9'd340: value = 12'h6EA;
            9'd341: value = 12'h6ED;
            9'd342: value = 12'h6F0;
            9'd343: value = 12'h6F3;
            9'd344: value = 12'h6F6;
            9'd345: value = 12'h6F9;
            9'd346: value = 12'h6FC;
            9'd347: value = 12'h6FF;
            9'd348: value = 12'h702;
            9'd349: value = 12'h705;
            9'd350: value = 12'h708;
            9'd351: value = 12'h70B;
            9'd352: value = 12'h70E;
            9'd353: value = 12'h711;
            9'd354: value = 12'h714;
            9'd355: value = 12'h717;
            9'd356: value = 12'h71A;
            9'd357: value = 12'h71D;
            9'd358: value = 12'h720;
            9'd359: value = 12'h723;
            9'd360: value = 12'h725;
            9'd361: value = 12'h728;
            9'd362: value = 12'h72B;
            9'd363: value = 12'h72E;
            9'd364: value = 12'h730;
            9'd365: value = 12'h733;
            9'd366: value = 12'h736;
            9'd367: value = 12'h739;
            9'd368: value = 12'h73B;
            9'd369: value = 12'h73E;
            9'd370: value = 12'h741;
            9'd371: value = 12'h743;
            9'd372: value = 12'h746;
            9'd373: value = 12'h748;
            9'd374: value = 12'h74B;
            9'd375: value = 12'h74E;
            9'd376: value = 12'h750;
            9'd377: value = 12'h753;
            9'd378: value = 12'h755;
            9'd379: value = 12'h758;
            9'd380: value = 12'h75A;
            9'd381: value = 12'h75D;
            9'd382: value = 12'h75F;
            9'd383: value = 12'h761;
            9'd384: value = 12'h764;
            9'd385: value = 12'h766;
            9'd386: value = 12'h769;
            9'd387: value = 12'h76B;
            9'd388: value = 12'h76D;
            9'd389: value = 12'h770;
            9'd390: value = 12'h772;
            9'd391: value = 12'h774;
            9'd392: value = 12'h776;
            9'd393: value = 12'h779;
            9'd394: value = 12'h77B;
            9'd395: value = 12'h77D;
            9'd396: value = 12'h77F;
            9'd397: value = 12'h781;
            9'd398: value = 12'h784;
            9'd399: value = 12'h786;
            9'd400: value = 12'h788;
            9'd401: value = 12'h78A;
            9'd402: value = 12'h78C;
            9'd403: value = 12'h78E;
            9'd404: value = 12'h790;
            9'd405: value = 12'h792;
            9'd406: value = 12'h794;
            9'd407: value = 12'h796;
            9'd408: value = 12'h798;
            9'd409: value = 12'h79A;
            9'd410: value = 12'h79C;
            9'd411: value = 12'h79E;
            9'd412: value = 12'h7A0;
            9'd413: value = 12'h7A2;
            9'd414: value = 12'h7A4;
            9'd415: value = 12'h7A5;
            9'd416: value = 12'h7A7;
            9'd417: value = 12'h7A9;
            9'd418: value = 12'h7AB;
            9'd419: value = 12'h7AD;
            9'd420: value = 12'h7AE;
            9'd421: value = 12'h7B0;
            9'd422: value = 12'h7B2;
            9'd423: value = 12'h7B4;
            9'd424: value = 12'h7B5;
            9'd425: value = 12'h7B7;
            9'd426: value = 12'h7B8;
            9'd427: value = 12'h7BA;
            9'd428: value = 12'h7BC;
            9'd429: value = 12'h7BD;
            9'd430: value = 12'h7BF;
            9'd431: value = 12'h7C0;
            9'd432: value = 12'h7C2;
            9'd433: value = 12'h7C3;
            9'd434: value = 12'h7C5;
            9'd435: value = 12'h7C6;
            9'd436: value = 12'h7C8;
            9'd437: value = 12'h7C9;
            9'd438: value = 12'h7CB;
            9'd439: value = 12'h7CC;
            9'd440: value = 12'h7CD;
            9'd441: value = 12'h7CF;
            9'd442: value = 12'h7D0;
            9'd443: value = 12'h7D1;
            9'd444: value = 12'h7D3;
            9'd445: value = 12'h7D4;
            9'd446: value = 12'h7D5;
            9'd447: value = 12'h7D7;
            9'd448: value = 12'h7D8;
            9'd449: value = 12'h7D9;
            9'd450: value = 12'h7DA;
            9'd451: value = 12'h7DB;
            9'd452: value = 12'h7DC;
            9'd453: value = 12'h7DE;
            9'd454: value = 12'h7DF;
            9'd455: value = 12'h7E0;
            9'd456: value = 12'h7E1;
            9'd457: value = 12'h7E2;
            9'd458: value = 12'h7E3;
            9'd459: value = 12'h7E4;
            9'd460: value = 12'h7E5;
            9'd461: value = 12'h7E6;
            9'd462: value = 12'h7E7;
            9'd463: value = 12'h7E8;
            9'd464: value = 12'h7E9;
            9'd465: value = 12'h7EA;
            9'd466: value = 12'h7EB;
            9'd467: value = 12'h7EB;
            9'd468: value = 12'h7EC;
            9'd469: value = 12'h7ED;
            9'd470: value = 12'h7EE;
            9'd471: value = 12'h7EF;
            9'd472: value = 12'h7EF;
            9'd473: value = 12'h7F0;
            9'd474: value = 12'h7F1;
            9'd475: value = 12'h7F2;
            9'd476: value = 12'h7F2;
            9'd477: value = 12'h7F3;
            9'd478: value = 12'h7F4;
            9'd479: value = 12'h7F4;
            9'd480: value = 12'h7F5;
            9'd481: value = 12'h7F6;
            9'd482: value = 12'h7F6;
            9'd483: value = 12'h7F7;
            9'd484: value = 12'h7F7;
            9'd485: value = 12'h7F8;
            9'd486: value = 12'h7F8;
            9'd487: value = 12'h7F9;
            9'd488: value = 12'h7F9;
            9'd489: value = 12'h7FA;
            9'd490: value = 12'h7FA;
            9'd491: value = 12'h7FA;
            9'd492: value = 12'h7FB;
            9'd493: value = 12'h7FB;
            9'd494: value = 12'h7FC;
            9'd495: value = 12'h7FC;
            9'd496: value = 12'h7FC;
            9'd497: value = 12'h7FC;
            9'd498: value = 12'h7FD;
            9'd499: value = 12'h7FD;
            9'd500: value = 12'h7FD;
            9'd501: value = 12'h7FD;
            9'd502: value = 12'h7FE;
            9'd503: value = 12'h7FE;
            9'd504: value = 12'h7FE;
            9'd505: value = 12'h7FE;
            9'd506: value = 12'h7FE;
            9'd507: value = 12'h7FE;
            9'd508: value = 12'h7FE;
            9'd509: value = 12'h7FE;
            9'd510: value = 12'h7FE;
            9'd511: value = 12'h7FE;

            default: value = 12'd0;
        endcase
    end

endmodule
