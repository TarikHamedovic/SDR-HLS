
module quarterwave_table #(
    parameter QLUT_DEPTH = 11,
    parameter DATA_WIDTH = 16
)(
    input  logic        [QLUT_DEPTH-3:0] address, // 9-bit address signal for 512 values
    output logic signed [DATA_WIDTH-1:0] value    // 16-bit output signal
);

    always_comb begin
        unique case(address)
            9'd0: value = 16'h32;
            9'd1: value = 16'h96;
            9'd2: value = 16'hFB;
            9'd3: value = 16'h15F;
            9'd4: value = 16'h1C4;
            9'd5: value = 16'h228;
            9'd6: value = 16'h28D;
            9'd7: value = 16'h2F1;
            9'd8: value = 16'h356;
            9'd9: value = 16'h3BA;
            9'd10: value = 16'h41F;
            9'd11: value = 16'h483;
            9'd12: value = 16'h4E8;
            9'd13: value = 16'h54C;
            9'd14: value = 16'h5B1;
            9'd15: value = 16'h615;
            9'd16: value = 16'h67A;
            9'd17: value = 16'h6DE;
            9'd18: value = 16'h742;
            9'd19: value = 16'h7A7;
            9'd20: value = 16'h80B;
            9'd21: value = 16'h86F;
            9'd22: value = 16'h8D4;
            9'd23: value = 16'h938;
            9'd24: value = 16'h99C;
            9'd25: value = 16'hA00;
            9'd26: value = 16'hA65;
            9'd27: value = 16'hAC9;
            9'd28: value = 16'hB2D;
            9'd29: value = 16'hB91;
            9'd30: value = 16'hBF5;
            9'd31: value = 16'hC59;
            9'd32: value = 16'hCBD;
            9'd33: value = 16'hD21;
            9'd34: value = 16'hD85;
            9'd35: value = 16'hDE9;
            9'd36: value = 16'hE4D;
            9'd37: value = 16'hEB1;
            9'd38: value = 16'hF15;
            9'd39: value = 16'hF79;
            9'd40: value = 16'hFDC;
            9'd41: value = 16'h1040;
            9'd42: value = 16'h10A4;
            9'd43: value = 16'h1107;
            9'd44: value = 16'h116B;
            9'd45: value = 16'h11CF;
            9'd46: value = 16'h1232;
            9'd47: value = 16'h1296;
            9'd48: value = 16'h12F9;
            9'd49: value = 16'h135D;
            9'd50: value = 16'h13C0;
            9'd51: value = 16'h1423;
            9'd52: value = 16'h1486;
            9'd53: value = 16'h14EA;
            9'd54: value = 16'h154D;
            9'd55: value = 16'h15B0;
            9'd56: value = 16'h1613;
            9'd57: value = 16'h1676;
            9'd58: value = 16'h16D9;
            9'd59: value = 16'h173C;
            9'd60: value = 16'h179F;
            9'd61: value = 16'h1801;
            9'd62: value = 16'h1864;
            9'd63: value = 16'h18C7;
            9'd64: value = 16'h1929;
            9'd65: value = 16'h198C;
            9'd66: value = 16'h19EE;
            9'd67: value = 16'h1A51;
            9'd68: value = 16'h1AB3;
            9'd69: value = 16'h1B15;
            9'd70: value = 16'h1B78;
            9'd71: value = 16'h1BDA;
            9'd72: value = 16'h1C3C;
            9'd73: value = 16'h1C9E;
            9'd74: value = 16'h1D00;
            9'd75: value = 16'h1D62;
            9'd76: value = 16'h1DC3;
            9'd77: value = 16'h1E25;
            9'd78: value = 16'h1E87;
            9'd79: value = 16'h1EE8;
            9'd80: value = 16'h1F4A;
            9'd81: value = 16'h1FAB;
            9'd82: value = 16'h200D;
            9'd83: value = 16'h206E;
            9'd84: value = 16'h20CF;
            9'd85: value = 16'h2130;
            9'd86: value = 16'h2191;
            9'd87: value = 16'h21F2;
            9'd88: value = 16'h2253;
            9'd89: value = 16'h22B4;
            9'd90: value = 16'h2315;
            9'd91: value = 16'h2375;
            9'd92: value = 16'h23D6;
            9'd93: value = 16'h2436;
            9'd94: value = 16'h2497;
            9'd95: value = 16'h24F7;
            9'd96: value = 16'h2557;
            9'd97: value = 16'h25B7;
            9'd98: value = 16'h2617;
            9'd99: value = 16'h2677;
            9'd100: value = 16'h26D7;
            9'd101: value = 16'h2737;
            9'd102: value = 16'h2797;
            9'd103: value = 16'h27F6;
            9'd104: value = 16'h2856;
            9'd105: value = 16'h28B5;
            9'd106: value = 16'h2914;
            9'd107: value = 16'h2973;
            9'd108: value = 16'h29D2;
            9'd109: value = 16'h2A31;
            9'd110: value = 16'h2A90;
            9'd111: value = 16'h2AEF;
            9'd112: value = 16'h2B4E;
            9'd113: value = 16'h2BAC;
            9'd114: value = 16'h2C0B;
            9'd115: value = 16'h2C69;
            9'd116: value = 16'h2CC7;
            9'd117: value = 16'h2D25;
            9'd118: value = 16'h2D83;
            9'd119: value = 16'h2DE1;
            9'd120: value = 16'h2E3F;
            9'd121: value = 16'h2E9D;
            9'd122: value = 16'h2EFA;
            9'd123: value = 16'h2F58;
            9'd124: value = 16'h2FB5;
            9'd125: value = 16'h3012;
            9'd126: value = 16'h306F;
            9'd127: value = 16'h30CC;
            9'd128: value = 16'h3129;
            9'd129: value = 16'h3186;
            9'd130: value = 16'h31E3;
            9'd131: value = 16'h323F;
            9'd132: value = 16'h329C;
            9'd133: value = 16'h32F8;
            9'd134: value = 16'h3354;
            9'd135: value = 16'h33B0;
            9'd136: value = 16'h340C;
            9'd137: value = 16'h3468;
            9'd138: value = 16'h34C3;
            9'd139: value = 16'h351F;
            9'd140: value = 16'h357A;
            9'd141: value = 16'h35D6;
            9'd142: value = 16'h3631;
            9'd143: value = 16'h368C;
            9'd144: value = 16'h36E7;
            9'd145: value = 16'h3741;
            9'd146: value = 16'h379C;
            9'd147: value = 16'h37F6;
            9'd148: value = 16'h3851;
            9'd149: value = 16'h38AB;
            9'd150: value = 16'h3905;
            9'd151: value = 16'h395F;
            9'd152: value = 16'h39B9;
            9'd153: value = 16'h3A12;
            9'd154: value = 16'h3A6C;
            9'd155: value = 16'h3AC5;
            9'd156: value = 16'h3B1F;
            9'd157: value = 16'h3B78;
            9'd158: value = 16'h3BD1;
            9'd159: value = 16'h3C29;
            9'd160: value = 16'h3C82;
            9'd161: value = 16'h3CDB;
            9'd162: value = 16'h3D33;
            9'd163: value = 16'h3D8B;
            9'd164: value = 16'h3DE3;
            9'd165: value = 16'h3E3B;
            9'd166: value = 16'h3E93;
            9'd167: value = 16'h3EEB;
            9'd168: value = 16'h3F42;
            9'd169: value = 16'h3F99;
            9'd170: value = 16'h3FF0;
            9'd171: value = 16'h4047;
            9'd172: value = 16'h409E;
            9'd173: value = 16'h40F5;
            9'd174: value = 16'h414C;
            9'd175: value = 16'h41A2;
            9'd176: value = 16'h41F8;
            9'd177: value = 16'h424E;
            9'd178: value = 16'h42A4;
            9'd179: value = 16'h42FA;
            9'd180: value = 16'h4350;
            9'd181: value = 16'h43A5;
            9'd182: value = 16'h43FA;
            9'd183: value = 16'h444F;
            9'd184: value = 16'h44A4;
            9'd185: value = 16'h44F9;
            9'd186: value = 16'h454E;
            9'd187: value = 16'h45A2;
            9'd188: value = 16'h45F6;
            9'd189: value = 16'h464A;
            9'd190: value = 16'h469E;
            9'd191: value = 16'h46F2;
            9'd192: value = 16'h4746;
            9'd193: value = 16'h4799;
            9'd194: value = 16'h47EC;
            9'd195: value = 16'h483F;
            9'd196: value = 16'h4892;
            9'd197: value = 16'h48E5;
            9'd198: value = 16'h4938;
            9'd199: value = 16'h498A;
            9'd200: value = 16'h49DC;
            9'd201: value = 16'h4A2E;
            9'd202: value = 16'h4A80;
            9'd203: value = 16'h4AD2;
            9'd204: value = 16'h4B23;
            9'd205: value = 16'h4B74;
            9'd206: value = 16'h4BC5;
            9'd207: value = 16'h4C16;
            9'd208: value = 16'h4C67;
            9'd209: value = 16'h4CB8;
            9'd210: value = 16'h4D08;
            9'd211: value = 16'h4D58;
            9'd212: value = 16'h4DA8;
            9'd213: value = 16'h4DF8;
            9'd214: value = 16'h4E48;
            9'd215: value = 16'h4E97;
            9'd216: value = 16'h4EE6;
            9'd217: value = 16'h4F35;
            9'd218: value = 16'h4F84;
            9'd219: value = 16'h4FD3;
            9'd220: value = 16'h5021;
            9'd221: value = 16'h5070;
            9'd222: value = 16'h50BE;
            9'd223: value = 16'h510C;
            9'd224: value = 16'h5159;
            9'd225: value = 16'h51A7;
            9'd226: value = 16'h51F4;
            9'd227: value = 16'h5241;
            9'd228: value = 16'h528E;
            9'd229: value = 16'h52DB;
            9'd230: value = 16'h5328;
            9'd231: value = 16'h5374;
            9'd232: value = 16'h53C0;
            9'd233: value = 16'h540C;
            9'd234: value = 16'h5458;
            9'd235: value = 16'h54A3;
            9'd236: value = 16'h54EF;
            9'd237: value = 16'h553A;
            9'd238: value = 16'h5585;
            9'd239: value = 16'h55CF;
            9'd240: value = 16'h561A;
            9'd241: value = 16'h5664;
            9'd242: value = 16'h56AE;
            9'd243: value = 16'h56F8;
            9'd244: value = 16'h5742;
            9'd245: value = 16'h578B;
            9'd246: value = 16'h57D4;
            9'd247: value = 16'h581D;
            9'd248: value = 16'h5866;
            9'd249: value = 16'h58AF;
            9'd250: value = 16'h58F7;
            9'd251: value = 16'h593F;
            9'd252: value = 16'h5987;
            9'd253: value = 16'h59CF;
            9'd254: value = 16'h5A16;
            9'd255: value = 16'h5A5E;
            9'd256: value = 16'h5AA5;
            9'd257: value = 16'h5AEC;
            9'd258: value = 16'h5B32;
            9'd259: value = 16'h5B79;
            9'd260: value = 16'h5BBF;
            9'd261: value = 16'h5C05;
            9'd262: value = 16'h5C4B;
            9'd263: value = 16'h5C90;
            9'd264: value = 16'h5CD6;
            9'd265: value = 16'h5D1B;
            9'd266: value = 16'h5D5F;
            9'd267: value = 16'h5DA4;
            9'd268: value = 16'h5DE9;
            9'd269: value = 16'h5E2D;
            9'd270: value = 16'h5E71;
            9'd271: value = 16'h5EB4;
            9'd272: value = 16'h5EF8;
            9'd273: value = 16'h5F3B;
            9'd274: value = 16'h5F7E;
            9'd275: value = 16'h5FC1;
            9'd276: value = 16'h6004;
            9'd277: value = 16'h6046;
            9'd278: value = 16'h6088;
            9'd279: value = 16'h60CA;
            9'd280: value = 16'h610C;
            9'd281: value = 16'h614D;
            9'd282: value = 16'h618E;
            9'd283: value = 16'h61CF;
            9'd284: value = 16'h6210;
            9'd285: value = 16'h6251;
            9'd286: value = 16'h6291;
            9'd287: value = 16'h62D1;
            9'd288: value = 16'h6311;
            9'd289: value = 16'h6350;
            9'd290: value = 16'h638F;
            9'd291: value = 16'h63CE;
            9'd292: value = 16'h640D;
            9'd293: value = 16'h644C;
            9'd294: value = 16'h648A;
            9'd295: value = 16'h64C8;
            9'd296: value = 16'h6506;
            9'd297: value = 16'h6544;
            9'd298: value = 16'h6581;
            9'd299: value = 16'h65BE;
            9'd300: value = 16'h65FB;
            9'd301: value = 16'h6638;
            9'd302: value = 16'h6674;
            9'd303: value = 16'h66B0;
            9'd304: value = 16'h66EC;
            9'd305: value = 16'h6728;
            9'd306: value = 16'h6763;
            9'd307: value = 16'h679E;
            9'd308: value = 16'h67D9;
            9'd309: value = 16'h6814;
            9'd310: value = 16'h684E;
            9'd311: value = 16'h6888;
            9'd312: value = 16'h68C2;
            9'd313: value = 16'h68FC;
            9'd314: value = 16'h6935;
            9'd315: value = 16'h696E;
            9'd316: value = 16'h69A7;
            9'd317: value = 16'h69E0;
            9'd318: value = 16'h6A18;
            9'd319: value = 16'h6A50;
            9'd320: value = 16'h6A88;
            9'd321: value = 16'h6AC0;
            9'd322: value = 16'h6AF7;
            9'd323: value = 16'h6B2E;
            9'd324: value = 16'h6B65;
            9'd325: value = 16'h6B9C;
            9'd326: value = 16'h6BD2;
            9'd327: value = 16'h6C08;
            9'd328: value = 16'h6C3E;
            9'd329: value = 16'h6C73;
            9'd330: value = 16'h6CA8;
            9'd331: value = 16'h6CDD;
            9'd332: value = 16'h6D12;
            9'd333: value = 16'h6D47;
            9'd334: value = 16'h6D7B;
            9'd335: value = 16'h6DAF;
            9'd336: value = 16'h6DE3;
            9'd337: value = 16'h6E16;
            9'd338: value = 16'h6E49;
            9'd339: value = 16'h6E7C;
            9'd340: value = 16'h6EAF;
            9'd341: value = 16'h6EE1;
            9'd342: value = 16'h6F13;
            9'd343: value = 16'h6F45;
            9'd344: value = 16'h6F76;
            9'd345: value = 16'h6FA8;
            9'd346: value = 16'h6FD9;
            9'd347: value = 16'h7009;
            9'd348: value = 16'h703A;
            9'd349: value = 16'h706A;
            9'd350: value = 16'h709A;
            9'd351: value = 16'h70CA;
            9'd352: value = 16'h70F9;
            9'd353: value = 16'h7128;
            9'd354: value = 16'h7157;
            9'd355: value = 16'h7186;
            9'd356: value = 16'h71B4;
            9'd357: value = 16'h71E2;
            9'd358: value = 16'h7210;
            9'd359: value = 16'h723D;
            9'd360: value = 16'h726A;
            9'd361: value = 16'h7297;
            9'd362: value = 16'h72C4;
            9'd363: value = 16'h72F0;
            9'd364: value = 16'h731C;
            9'd365: value = 16'h7348;
            9'd366: value = 16'h7374;
            9'd367: value = 16'h739F;
            9'd368: value = 16'h73CA;
            9'd369: value = 16'h73F5;
            9'd370: value = 16'h741F;
            9'd371: value = 16'h7449;
            9'd372: value = 16'h7473;
            9'd373: value = 16'h749D;
            9'd374: value = 16'h74C6;
            9'd375: value = 16'h74EF;
            9'd376: value = 16'h7518;
            9'd377: value = 16'h7540;
            9'd378: value = 16'h7568;
            9'd379: value = 16'h7590;
            9'd380: value = 16'h75B8;
            9'd381: value = 16'h75DF;
            9'd382: value = 16'h7606;
            9'd383: value = 16'h762D;
            9'd384: value = 16'h7653;
            9'd385: value = 16'h767A;
            9'd386: value = 16'h76A0;
            9'd387: value = 16'h76C5;
            9'd388: value = 16'h76EA;
            9'd389: value = 16'h7710;
            9'd390: value = 16'h7734;
            9'd391: value = 16'h7759;
            9'd392: value = 16'h777D;
            9'd393: value = 16'h77A1;
            9'd394: value = 16'h77C4;
            9'd395: value = 16'h77E8;
            9'd396: value = 16'h780B;
            9'd397: value = 16'h782E;
            9'd398: value = 16'h7850;
            9'd399: value = 16'h7872;
            9'd400: value = 16'h7894;
            9'd401: value = 16'h78B6;
            9'd402: value = 16'h78D7;
            9'd403: value = 16'h78F8;
            9'd404: value = 16'h7919;
            9'd405: value = 16'h7939;
            9'd406: value = 16'h7959;
            9'd407: value = 16'h7979;
            9'd408: value = 16'h7998;
            9'd409: value = 16'h79B8;
            9'd410: value = 16'h79D7;
            9'd411: value = 16'h79F5;
            9'd412: value = 16'h7A14;
            9'd413: value = 16'h7A32;
            9'd414: value = 16'h7A4F;
            9'd415: value = 16'h7A6D;
            9'd416: value = 16'h7A8A;
            9'd417: value = 16'h7AA7;
            9'd418: value = 16'h7AC4;
            9'd419: value = 16'h7AE0;
            9'd420: value = 16'h7AFC;
            9'd421: value = 16'h7B18;
            9'd422: value = 16'h7B33;
            9'd423: value = 16'h7B4E;
            9'd424: value = 16'h7B69;
            9'd425: value = 16'h7B83;
            9'd426: value = 16'h7B9E;
            9'd427: value = 16'h7BB8;
            9'd428: value = 16'h7BD1;
            9'd429: value = 16'h7BEB;
            9'd430: value = 16'h7C04;
            9'd431: value = 16'h7C1C;
            9'd432: value = 16'h7C35;
            9'd433: value = 16'h7C4D;
            9'd434: value = 16'h7C65;
            9'd435: value = 16'h7C7C;
            9'd436: value = 16'h7C93;
            9'd437: value = 16'h7CAA;
            9'd438: value = 16'h7CC1;
            9'd439: value = 16'h7CD7;
            9'd440: value = 16'h7CED;
            9'd441: value = 16'h7D03;
            9'd442: value = 16'h7D18;
            9'd443: value = 16'h7D2E;
            9'd444: value = 16'h7D42;
            9'd445: value = 16'h7D57;
            9'd446: value = 16'h7D6B;
            9'd447: value = 16'h7D7F;
            9'd448: value = 16'h7D93;
            9'd449: value = 16'h7DA6;
            9'd450: value = 16'h7DB9;
            9'd451: value = 16'h7DCC;
            9'd452: value = 16'h7DDE;
            9'd453: value = 16'h7DF0;
            9'd454: value = 16'h7E02;
            9'd455: value = 16'h7E13;
            9'd456: value = 16'h7E25;
            9'd457: value = 16'h7E36;
            9'd458: value = 16'h7E46;
            9'd459: value = 16'h7E56;
            9'd460: value = 16'h7E66;
            9'd461: value = 16'h7E76;
            9'd462: value = 16'h7E85;
            9'd463: value = 16'h7E94;
            9'd464: value = 16'h7EA3;
            9'd465: value = 16'h7EB2;
            9'd466: value = 16'h7EC0;
            9'd467: value = 16'h7ECE;
            9'd468: value = 16'h7EDB;
            9'd469: value = 16'h7EE8;
            9'd470: value = 16'h7EF5;
            9'd471: value = 16'h7F02;
            9'd472: value = 16'h7F0E;
            9'd473: value = 16'h7F1A;
            9'd474: value = 16'h7F26;
            9'd475: value = 16'h7F31;
            9'd476: value = 16'h7F3C;
            9'd477: value = 16'h7F47;
            9'd478: value = 16'h7F52;
            9'd479: value = 16'h7F5C;
            9'd480: value = 16'h7F66;
            9'd481: value = 16'h7F6F;
            9'd482: value = 16'h7F78;
            9'd483: value = 16'h7F81;
            9'd484: value = 16'h7F8A;
            9'd485: value = 16'h7F92;
            9'd486: value = 16'h7F9A;
            9'd487: value = 16'h7FA2;
            9'd488: value = 16'h7FA9;
            9'd489: value = 16'h7FB0;
            9'd490: value = 16'h7FB7;
            9'd491: value = 16'h7FBE;
            9'd492: value = 16'h7FC4;
            9'd493: value = 16'h7FCA;
            9'd494: value = 16'h7FCF;
            9'd495: value = 16'h7FD5;
            9'd496: value = 16'h7FD9;
            9'd497: value = 16'h7FDE;
            9'd498: value = 16'h7FE2;
            9'd499: value = 16'h7FE6;
            9'd500: value = 16'h7FEA;
            9'd501: value = 16'h7FEE;
            9'd502: value = 16'h7FF1;
            9'd503: value = 16'h7FF3;
            9'd504: value = 16'h7FF6;
            9'd505: value = 16'h7FF8;
            9'd506: value = 16'h7FFA;
            9'd507: value = 16'h7FFB;
            9'd508: value = 16'h7FFD;
            9'd509: value = 16'h7FFE;
            9'd510: value = 16'h7FFE;
            9'd511: value = 16'h7FFE;

            default: value = 16'd0;
        endcase
    end

endmodule
