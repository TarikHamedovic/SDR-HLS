// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.13.0.56.2
// Netlist written on Thu May 30 00:34:09 2024
//
// Verilog Description of module top
//

module top (clk_25mhz, i_Rx_Serial, RFIn, o_Tx_Serial, led, XOut, 
            DiffOut, PWMOut, PWMOutP1, PWMOutP2, PWMOutP3, PWMOutP4, 
            PWMOutN1, PWMOutN2, PWMOutN3, PWMOutN4, sinGen, sin_out, 
            CIC_out_clkSin) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(39[8:11])
    input clk_25mhz;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(40[22:31])
    input i_Rx_Serial;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(41[22:33])
    input RFIn;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(42[22:26])
    output o_Tx_Serial;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(43[22:33])
    output [7:0]led;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    output XOut;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(45[22:26])
    output DiffOut;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(46[22:29])
    output PWMOut;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(47[22:28])
    output PWMOutP1;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(48[22:30])
    output PWMOutP2;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(49[22:30])
    output PWMOutP3;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(50[22:30])
    output PWMOutP4;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(51[22:30])
    output PWMOutN1;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(52[22:30])
    output PWMOutN2;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(53[22:30])
    output PWMOutN3;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(54[22:30])
    output PWMOutN4;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(55[22:30])
    output sinGen;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(56[22:28])
    output sin_out;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(57[22:29])
    output CIC_out_clkSin;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(58[22:36])
    
    wire clk_25mhz_c /* synthesis is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(40[22:31])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(61[23:32])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(74[23:38])
    
    wire GND_net, VCC_net, i_Rx_Serial_c, RFIn_c, led_c_7, led_c_6, 
        led_c_5, led_c_4, led_c_3, led_c_2, led_c_1, led_c_0, DiffOut_c, 
        PWMOutP4_c, PWMOutN4_c, sinGen_c, o_Rx_DV, o_Rx_DV1;
    wire [7:0]o_Rx_Byte1;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(67[23:33])
    wire [11:0]MixerOutSin;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(70[23:34])
    wire [11:0]MixerOutCos;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(71[23:34])
    wire [11:0]CIC1_outCos;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(76[23:34])
    wire [63:0]phase_accum;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(78[23:34])
    wire [12:0]LOSine;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(79[23:29])
    wire [12:0]LOCosine;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(80[23:31])
    wire [63:0]phase_inc_carrGen;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(82[23:40])
    wire [63:0]phase_inc_carrGen1;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(83[23:41])
    wire [11:0]DemodOut;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(85[23:31])
    
    wire n24, n25, n26, n27, n28, n29, n30, n31;
    wire [7:0]CICGain;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(86[23:30])
    
    wire n16626, n7, n6, n5, n4, n3, n2, n37, n36, n35, 
        n34, n33, n32, n31_adj_2808, n30_adj_2809, n29_adj_2810, 
        n28_adj_2811, n27_adj_2812, n26_adj_2813, n25_adj_2814, n24_adj_2815, 
        n23, n22, n21, n20, n19, n18, n17, cout, n16625, n16624, 
        n16, n15, n14, n13, n12, n11, n10, n9, n8, n7_adj_2816, 
        n6_adj_2817, n5_adj_2818, n4_adj_2819, n3_adj_2820, n2_adj_2821, 
        n16623, n16388, n16387, n16622, n16621, n2422, n16620, 
        n16619, n16618, n16617, n16616, n16615, n16614, n16613, 
        n16612, n16607, n16606, n16605, n16604, n16603, n16597, 
        n16596, n16595, n16594, n16593, n2393, n16592, n2388, 
        n16586, n16585, n16584, n16583, n16582, n16581, n16580, 
        n16579, n16577, n16576, n16575, n16160;
    wire [63:0]phase_accum_adj_5732;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(26[28:39])
    
    wire n16159, n16156, n16155, n16154;
    wire [11:0]MixerOutSin_11__N_236;
    wire [11:0]MixerOutCos_11__N_250;
    
    wire n2332;
    wire [71:0]d_tmp;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(52[28:33])
    wire [71:0]d_d_tmp;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(52[35:42])
    wire [71:0]d1;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(53[28:30])
    wire [71:0]d2;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(53[32:34])
    wire [71:0]d3;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(53[36:38])
    wire [71:0]d4;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(53[40:42])
    wire [71:0]d5;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(53[44:46])
    wire [71:0]d6;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[28:30])
    wire [71:0]d_d6;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[32:36])
    wire [71:0]d7;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[38:40])
    wire [71:0]d_d7;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[42:46])
    wire [71:0]d8;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[48:50])
    wire [71:0]d_d8;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[52:56])
    wire [71:0]d9;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[58:60])
    wire [71:0]d_d9;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[62:66])
    wire [71:0]d10;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[68:71])
    
    wire n16386;
    wire [15:0]count;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(56[28:33])
    wire [71:0]d1_71__N_418;
    wire [71:0]d2_71__N_490;
    wire [71:0]d3_71__N_562;
    wire [71:0]d4_71__N_634;
    wire [71:0]d5_71__N_706;
    
    wire n16574, n16170, n16573, n16572, n16571, n16565, n16564, 
        n16563, n16562, n16561, n16560, n16559, n16174, n32_adj_2822, 
        n23_adj_2823;
    wire [71:0]d6_71__N_1459;
    wire [71:0]d7_71__N_1531;
    wire [71:0]d8_71__N_1603;
    wire [71:0]d9_71__N_1675;
    
    wire n16385;
    wire [71:0]d_out_11__N_1819;
    
    wire cout_adj_2824, n183, n180, n177, n174, n171, n168, n165, 
        n162, n159, n156, n153, n150, n147, n144, n141, n138, 
        n135, n132, n129, n126, n123, n120, n117, n114, n111, 
        n108, n105, n102, n99, n96, n93, n90, n87, n84, n81, 
        n78, n183_adj_2825, n180_adj_2826, n177_adj_2827, n174_adj_2828, 
        n171_adj_2829, n168_adj_2830, n165_adj_2831, n162_adj_2832, 
        n159_adj_2833, n156_adj_2834, n153_adj_2835, n150_adj_2836, 
        n147_adj_2837, n144_adj_2838, n141_adj_2839, n138_adj_2840, 
        n135_adj_2841, n132_adj_2842, n129_adj_2843, n126_adj_2844, 
        n123_adj_2845, n120_adj_2846, n117_adj_2847, n114_adj_2848, 
        n111_adj_2849, n108_adj_2850, n105_adj_2851, n102_adj_2852, 
        n99_adj_2853, n96_adj_2854, n93_adj_2855, n90_adj_2856, n87_adj_2857, 
        n84_adj_2858, n81_adj_2859, n78_adj_2860;
    wire [71:0]d_tmp_adj_5738;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(52[28:33])
    wire [71:0]d_d_tmp_adj_5739;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(52[35:42])
    wire [71:0]d1_adj_5740;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(53[28:30])
    wire [71:0]d2_adj_5741;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(53[32:34])
    wire [71:0]d3_adj_5742;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(53[36:38])
    wire [71:0]d4_adj_5743;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(53[40:42])
    wire [71:0]d5_adj_5744;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(53[44:46])
    wire [71:0]d6_adj_5745;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[28:30])
    wire [71:0]d_d6_adj_5746;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[32:36])
    wire [71:0]d7_adj_5747;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[38:40])
    wire [71:0]d_d7_adj_5748;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[42:46])
    wire [71:0]d8_adj_5749;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[48:50])
    wire [71:0]d_d8_adj_5750;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[52:56])
    wire [71:0]d9_adj_5751;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[58:60])
    wire [71:0]d_d9_adj_5752;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[62:66])
    wire [71:0]d10_adj_5753;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[68:71])
    wire [15:0]count_adj_5755;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(56[28:33])
    wire [71:0]d1_71__N_418_adj_5756;
    wire [71:0]d2_71__N_490_adj_5757;
    wire [71:0]d3_71__N_562_adj_5758;
    wire [71:0]d4_71__N_634_adj_5759;
    wire [71:0]d5_71__N_706_adj_5760;
    
    wire n16384, n16558, n16557, n16551, n16550, n16549, n16548, 
        n16547, n16546, n16545, n16544, n321, n318, n315, n312, 
        n309, n306, n303, n300, n297, n294, n291, n288, n285, 
        n282, n279, n276, n273, n270, n267;
    wire [71:0]d6_71__N_1459_adj_5772;
    wire [71:0]d7_71__N_1531_adj_5773;
    wire [71:0]d8_71__N_1603_adj_5774;
    wire [71:0]d9_71__N_1675_adj_5775;
    
    wire n16153, n16152, n16151, n16150, n16149, n16148, n16147, 
        n16146, n16145, n16144, n16143, n16142, n16141, n16140, 
        n16139, n16135, n16134, n16133, n16132, n16131, n16130, 
        n16129, n16128, n16127, n16126, n16125, n16124, n16123, 
        n16122;
    wire [71:0]d_out_11__N_1819_adj_5778;
    
    wire n264, n261, n258, n255, n252, n249, n246, n243, n240, 
        n237, n234, n231, n228, n225, n222, n219, n216, n213, 
        n210, n207, n204, n201, n198, n195, n192, n189, n186, 
        n183_adj_4607, n180_adj_4608, n177_adj_4609, n174_adj_4610, 
        n171_adj_4611, n168_adj_4612, n165_adj_4613, n162_adj_4614, 
        n159_adj_4615, n156_adj_4616, n153_adj_4617, n150_adj_4618, 
        n147_adj_4619, n144_adj_4620, n141_adj_4621, n138_adj_4622, 
        n135_adj_4623, n132_adj_4624, cout_adj_4625, n16383, n16248, 
        n16382, n16381, n16247, n16377, n16376, n16250, n16375, 
        n16374, n16373;
    wire [9:0]counter;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(36[12:19])
    wire [11:0]DataInReg;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(39[12:21])
    wire [11:0]DataInReg_11__N_1856;
    
    wire n16121, n16120;
    wire [31:0]ISquare;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(33[28:35])
    
    wire n3_adj_4626, n2_adj_4627, n16372;
    wire [11:0]MultDataB;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(38[28:37])
    wire [23:0]MultResult1;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(39[28:39])
    wire [23:0]MultResult2;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(43[28:39])
    
    wire n21_adj_4628, n20_adj_4629, n19_adj_4630, n18_adj_4631, n17_adj_4632, 
        n16_adj_4633, n15_adj_4634, n16371, n2328, n16370, n16369, 
        n2327, n14_adj_4635, n16246, n2326, n2325, n13_adj_4636, 
        n16368, n16367, n213_adj_4637, n2324, n2323, n12_adj_4638, 
        n2322, n2321, n37_adj_4639, n36_adj_4640, n35_adj_4641, n34_adj_4642, 
        n33_adj_4643, n32_adj_4644, n31_adj_4645, n30_adj_4646, n29_adj_4647, 
        n28_adj_4648, n27_adj_4649, n26_adj_4650, n11_adj_4651, n25_adj_4652, 
        n2320, n24_adj_4653, n23_adj_4654, n22_adj_4655, n21_adj_4656, 
        n20_adj_4657, n19_adj_4658, n18_adj_4659, n17_adj_4660, n16_adj_4661, 
        n15_adj_4662, n14_adj_4663, n13_adj_4664, n12_adj_4665, n11_adj_4666, 
        n10_adj_4667, n9_adj_4668, n8_adj_4669, n7_adj_4670, n6_adj_4671, 
        n5_adj_4672, n4_adj_4673, n3_adj_4674, n2_adj_4675;
    wire [17:0]d_out_d_11__N_1874;
    
    wire d_out_d_11__N_1873, n10_adj_4676, n2318, n2317, n37_adj_4677, 
        n36_adj_4678, n35_adj_4679, n34_adj_4680, n33_adj_4681, n32_adj_4682, 
        n31_adj_4683;
    wire [17:0]d_out_d_11__N_1876;
    
    wire d_out_d_11__N_1875, n9_adj_4684, n30_adj_4685, n29_adj_4686, 
        n28_adj_4687, n27_adj_4688, n26_adj_4689, n25_adj_4690, n24_adj_4691, 
        n23_adj_4692, n22_adj_4693, n21_adj_4694, n20_adj_4695, n19_adj_4696, 
        n18_adj_4697, n17_adj_4698, n16_adj_4699, n15_adj_4700, n14_adj_4701, 
        n13_adj_4702, n2315, n12_adj_4703, n11_adj_4704, n10_adj_4705, 
        n9_adj_4706, n8_adj_4707, n7_adj_4708, n6_adj_4709, n5_adj_4710, 
        n4_adj_4711, n3_adj_4712, n2_adj_4713;
    wire [17:0]d_out_d_11__N_1878;
    
    wire d_out_d_11__N_1877, n8_adj_4714, n2313, n37_adj_4715, n36_adj_4716;
    wire [17:0]d_out_d_11__N_1880;
    
    wire d_out_d_11__N_1879, n7_adj_4717, n35_adj_4718, n2312, n34_adj_4719, 
        n33_adj_4720, n32_adj_4721, n31_adj_4722, n30_adj_4723, n29_adj_4724, 
        n28_adj_4725, n27_adj_4726, n26_adj_4727, n25_adj_4728, n24_adj_4729, 
        n23_adj_4730, n22_adj_4731, n21_adj_4732, n20_adj_4733, n19_adj_4734, 
        n18_adj_4735, n2311, n17_adj_4736, n16_adj_4737, n15_adj_4738, 
        n14_adj_4739, n13_adj_4740, n9_adj_4741, n10_adj_4742, n11_adj_4743, 
        n12_adj_4744, n8_adj_4745;
    wire [17:0]d_out_d_11__N_1882;
    
    wire n6_adj_4746, n37_adj_4747, n5_adj_4748, n4_adj_4749, n3_adj_4750, 
        n2_adj_4751, n36_adj_4752, n35_adj_4753, n34_adj_4754, n33_adj_4755;
    wire [17:0]d_out_d_11__N_1884;
    
    wire cout_adj_4756, n16206, n16175, n16176, n16180, n16181, 
        n16182, n16183, n16184, n16185, n16186, n16187, n3692, 
        n16189, n16190, n16208, n16192, n16193, n16194, n16195, 
        n16196, n16197, n16202, n16203, n3678, n3677;
    wire [17:0]d_out_d_11__N_1886;
    
    wire n16207, n16188, n16209, n16213, n16210, n16211, n16212, 
        n16204, n16214, n16215, n16216, n16217, n16226, n16205, 
        n3660, n16245, n3657, n16224, n16223, n16225, n16169, 
        n16168, n16167, n16119, n16166, n16165;
    wire [17:0]d_out_d_11__N_1888;
    
    wire n16366, n37_adj_4757, n36_adj_4758, n35_adj_4759;
    wire [17:0]d_out_d_11__N_1890;
    
    wire n34_adj_4760, n33_adj_4761, n32_adj_4762, n31_adj_4763, n30_adj_4764, 
        n29_adj_4765, n28_adj_4766, n27_adj_4767, n26_adj_4768, n25_adj_4769, 
        n24_adj_4770, n23_adj_4771, n22_adj_4772, n21_adj_4773, n20_adj_4774, 
        n19_adj_4775, n18_adj_4776, n17_adj_4777, n16_adj_4778, n15_adj_4779, 
        n14_adj_4780, n13_adj_4781, n12_adj_4782, n11_adj_4783, n10_adj_4784, 
        n9_adj_4785, n8_adj_4786, n7_adj_4787, n6_adj_4788, n5_adj_4789, 
        n16244;
    wire [17:0]d_out_d_11__N_1892;
    
    wire n916, n917, n918, n919, n920, n921, n922, n923, n924, 
        n925, n926, n927, n928, n929, n930, n931, n4_adj_4790;
    wire [17:0]d_out_d_11__N_2401;
    
    wire n16365, n16243, n16543;
    wire [17:0]d_out_d_11__N_2383;
    
    wire n16364, r_Rx_Data, n17948;
    wire [7:0]r_Rx_Byte;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(41[17:26])
    
    wire n16363, n16362, n16361, n16360, n2333, n16358, n16357, 
        n16356, n2337, n16118, n16355, n2335, n2336, n16523, n16522, 
        n16521, n17900, n16117, n11_adj_4791, n16116, n16242, n16354, 
        n16353, n16352, n16351, n16350, n2334, n16520, n16519, 
        n16518, n16517, n16516, n16515, n16514, n16513, n16512, 
        n16115, n16114, n16113, n16349, n16348, n16347, n16346, 
        n16511, n16510, n16509, n16508, n16507, n16506, n16112, 
        n16111, n16110, n16109, n16108, n16107, n16106, n16105, 
        n16104, n16103, n16102, n16101, n16100, n16098, n16097, 
        n16096, n16095, n16094, n16093, n2329, n16345, n16092, 
        n16344, n17930, n17929, n63, n64, n65, n66, n16091, 
        n16343, n17946, n131, n132_adj_4792, n133, n134, n135_adj_4793, 
        n136, n17945, n16090, n15227, n16342, n16089, n16341, 
        n16164, n2367, n2366, n16088, n2365, n2364, n2363, n2362, 
        n2361, n2359, n2358, n2357, n2356, n2355, n2354, n2353, 
        n2351, n2348, n2347, n2346, n2558, n16504, n2554, n16503, 
        n12306, n16502, n16163, n12304, n2542, n16162, n16161, 
        n15226, n12302, n16501, n16500, n12300, n16499, n2521, 
        n12298, n16498, n12296, n16497, n2515, n16496, n12292, 
        n16495, n16494, n16493, n16087, n16340, n16339, n16338, 
        n16337, n16336, n16335, n16334, n16333, n16332, n16331, 
        n16330, n16329, n16328, n16327, n16326, n13_adj_4794, n17630, 
        n16492, n16325, n16324, n15225, n16086, n16085, n16323, 
        n17926, n63_adj_4795, n64_adj_4796, n65_adj_4797, n66_adj_4798, 
        n16084, n17943, n131_adj_4799, n132_adj_4800, n133_adj_4801, 
        n134_adj_4802, n135_adj_4803, n136_adj_4804, n16083, n16082, 
        n16081, n16321, n16080, n17942, n16320, n16491, n16490, 
        n16489, n16079, n16078, n16488, n16487, n2430, n2345, 
        n2344, n2343, n2342, n2341, n2340, n2339, n2338, n16077, 
        n15_adj_4805, n14_adj_4806, n13_adj_4807, n12_adj_4808, n11_adj_4809, 
        n10_adj_4810, n9_adj_4811, n8_adj_4812, n7_adj_4813, n6_adj_4814, 
        n5_adj_4815, n4_adj_4816, n3_adj_4817, n2_adj_4818, n16076, 
        n16075, n16074, n16073, n16072, n16071, n16070, n16069, 
        n16068, n16482, n16481, n16480, n16479, n16478, n16477, 
        n2572, n16319, n16476, n2565, n16475, n16474, n16473, 
        n37_adj_4819, n36_adj_4820, n35_adj_4821, n34_adj_4822, n16472, 
        n33_adj_4823, n32_adj_4824, n31_adj_4825, n30_adj_4826, n29_adj_4827, 
        n28_adj_4828, n27_adj_4829, n26_adj_4830, n25_adj_4831, n24_adj_4832, 
        n2425, n16067, n16066, n2824, n16065, n16318, n16064, 
        n16063, n16062, n16241, n16061, n12563, n16060, n16059, 
        n16317, n16058, n16316, n16057, n16718, n16056, n17_adj_4833, 
        n16_adj_4834, n16055, n18_adj_4835, n35_adj_4836, n34_adj_4837, 
        n33_adj_4838, n32_adj_4839, n31_adj_4840, n30_adj_4841, n29_adj_4842, 
        n28_adj_4843, n27_adj_4844, n26_adj_4845, n25_adj_4846, n24_adj_4847, 
        n23_adj_4848, n22_adj_4849, n21_adj_4850, n20_adj_4851, n19_adj_4852, 
        n36_adj_4853, n37_adj_4854, n16054, n16053, n16052, n16051, 
        n32_adj_4855, n16050, n23_adj_4856, n16315, n16471, n16049, 
        n16239, n23_adj_4857, n22_adj_4858, n21_adj_4859, n20_adj_4860, 
        n19_adj_4861, n18_adj_4862, n17_adj_4863, n16_adj_4864, n15_adj_4865, 
        n14_adj_4866, n13_adj_4867, n12_adj_4868, n11_adj_4869, n10_adj_4870, 
        n9_adj_4871, n8_adj_4872, n7_adj_4873, n6_adj_4874, n5_adj_4875, 
        n4_adj_4876, n3_adj_4877, n2_adj_4878, n22_adj_4879, n16470, 
        n78_adj_4880, n81_adj_4881, n84_adj_4882, n87_adj_4883, n90_adj_4884, 
        n93_adj_4885, n96_adj_4886, n99_adj_4887, n102_adj_4888, n105_adj_4889, 
        n108_adj_4890, n111_adj_4891, n114_adj_4892, n117_adj_4893, 
        n120_adj_4894, n123_adj_4895, n126_adj_4896, n129_adj_4897, 
        n132_adj_4898, n135_adj_4899, n138_adj_4900, n141_adj_4901, 
        n144_adj_4902, n147_adj_4903, n150_adj_4904, n153_adj_4905, 
        n156_adj_4906, n159_adj_4907, n162_adj_4908, n165_adj_4909, 
        n168_adj_4910, n171_adj_4911, n174_adj_4912, n177_adj_4913, 
        n180_adj_4914, n183_adj_4915, n78_adj_4916, n81_adj_4917, n84_adj_4918, 
        n87_adj_4919, n90_adj_4920, n93_adj_4921, n96_adj_4922, n99_adj_4923, 
        n102_adj_4924, n105_adj_4925, n108_adj_4926, n111_adj_4927, 
        n114_adj_4928, n117_adj_4929, n120_adj_4930, n123_adj_4931, 
        n126_adj_4932, n129_adj_4933, n132_adj_4934, n135_adj_4935, 
        n138_adj_4936, n141_adj_4937, n144_adj_4938, n147_adj_4939, 
        n150_adj_4940, n153_adj_4941, n156_adj_4942, n159_adj_4943, 
        n162_adj_4944, n165_adj_4945, n168_adj_4946, n171_adj_4947, 
        n174_adj_4948, n177_adj_4949, n180_adj_4950, n183_adj_4951, 
        n78_adj_4952, n81_adj_4953, n84_adj_4954, n87_adj_4955, n90_adj_4956, 
        n93_adj_4957, n96_adj_4958, n99_adj_4959, n102_adj_4960, n105_adj_4961, 
        n108_adj_4962, n111_adj_4963, n114_adj_4964, n117_adj_4965, 
        n120_adj_4966, n123_adj_4967, n126_adj_4968, n129_adj_4969, 
        n132_adj_4970, n135_adj_4971, n138_adj_4972, n141_adj_4973, 
        n144_adj_4974, n147_adj_4975, n150_adj_4976, n153_adj_4977, 
        n156_adj_4978, n159_adj_4979, n162_adj_4980, n165_adj_4981, 
        n168_adj_4982, n171_adj_4983, n174_adj_4984, n177_adj_4985, 
        n180_adj_4986, n183_adj_4987, n78_adj_4988, n81_adj_4989, n84_adj_4990, 
        n87_adj_4991, n90_adj_4992, n93_adj_4993, n96_adj_4994, n99_adj_4995, 
        n102_adj_4996, n105_adj_4997, n108_adj_4998, n111_adj_4999, 
        n114_adj_5000, n117_adj_5001, n120_adj_5002, n123_adj_5003, 
        n126_adj_5004, n129_adj_5005, n132_adj_5006, n135_adj_5007, 
        n138_adj_5008, n141_adj_5009, n144_adj_5010, n147_adj_5011, 
        n150_adj_5012, n153_adj_5013, n156_adj_5014, n159_adj_5015, 
        n162_adj_5016, n165_adj_5017, n168_adj_5018, n171_adj_5019, 
        n174_adj_5020, n177_adj_5021, n180_adj_5022, n183_adj_5023, 
        n78_adj_5024, n81_adj_5025, n84_adj_5026, n87_adj_5027, n90_adj_5028, 
        n93_adj_5029, n96_adj_5030, n99_adj_5031, n102_adj_5032, n105_adj_5033, 
        n108_adj_5034, n111_adj_5035, n114_adj_5036, n117_adj_5037, 
        n120_adj_5038, n78_adj_5039, n81_adj_5040, n84_adj_5041, n87_adj_5042, 
        n90_adj_5043, n93_adj_5044, n96_adj_5045, n99_adj_5046, n102_adj_5047, 
        n105_adj_5048, n108_adj_5049, n111_adj_5050, n114_adj_5051, 
        n117_adj_5052, n120_adj_5053, n123_adj_5054, n126_adj_5055, 
        n129_adj_5056, n132_adj_5057, n135_adj_5058, n138_adj_5059, 
        n141_adj_5060, n144_adj_5061, n147_adj_5062, n150_adj_5063, 
        n153_adj_5064, n156_adj_5065, n159_adj_5066, n162_adj_5067, 
        n165_adj_5068, n168_adj_5069, n171_adj_5070, n174_adj_5071, 
        n177_adj_5072, n180_adj_5073, n183_adj_5074, n78_adj_5075, n81_adj_5076, 
        n84_adj_5077, n87_adj_5078, n90_adj_5079, n93_adj_5080, n96_adj_5081, 
        n99_adj_5082, n102_adj_5083, n105_adj_5084, n108_adj_5085, n111_adj_5086, 
        n114_adj_5087, n117_adj_5088, n120_adj_5089, n123_adj_5090, 
        n126_adj_5091, n129_adj_5092, n132_adj_5093, n135_adj_5094, 
        n138_adj_5095, n141_adj_5096, n144_adj_5097, n147_adj_5098, 
        n150_adj_5099, n153_adj_5100, n156_adj_5101, n159_adj_5102, 
        n162_adj_5103, n165_adj_5104, n168_adj_5105, n171_adj_5106, 
        n174_adj_5107, n177_adj_5108, n180_adj_5109, n183_adj_5110, 
        n134_adj_5111, n137, n140, n143, n146, n149, n152, n155, 
        n158, n161, n164, n167, n170, n173, n176, n179, n182, 
        n185, n188, n191, n194, n197, n200, n203, n206, n209, 
        n212, n215, n218, n221, n224, n227, n230, n233, n236, 
        n239, n242, n245, n248, n251, n254, n257, n260, n263, 
        n266, n269, n272, n275, n278, n281, n284, n287, n290, 
        n293, n296, n299, n302, n305, n308, n311, n314, n317, 
        n320, n323, n16048, n16047, n16046, n16045, n16044, n16043, 
        n16042, n16041, n16040, n16039, cout_adj_5112, cout_adj_5113, 
        n78_adj_5114, n81_adj_5115, n84_adj_5116, n87_adj_5117, n90_adj_5118, 
        n93_adj_5119, n96_adj_5120, n99_adj_5121, n102_adj_5122, n105_adj_5123, 
        n108_adj_5124, n111_adj_5125, n114_adj_5126, n117_adj_5127, 
        n120_adj_5128, n123_adj_5129, n126_adj_5130, n129_adj_5131, 
        n132_adj_5132, n135_adj_5133, n138_adj_5134, n141_adj_5135, 
        n144_adj_5136, n147_adj_5137, n150_adj_5138, n153_adj_5139, 
        n156_adj_5140, n159_adj_5141, n162_adj_5142, n165_adj_5143, 
        n168_adj_5144, n171_adj_5145, n174_adj_5146, n177_adj_5147, 
        n180_adj_5148, n183_adj_5149, n78_adj_5150, n81_adj_5151, n84_adj_5152, 
        n87_adj_5153, n90_adj_5154, n93_adj_5155, n96_adj_5156, n99_adj_5157, 
        n102_adj_5158, n105_adj_5159, n108_adj_5160, n111_adj_5161, 
        n114_adj_5162, n117_adj_5163, n120_adj_5164, n123_adj_5165, 
        n126_adj_5166, n129_adj_5167, n132_adj_5168, n135_adj_5169, 
        n138_adj_5170, n141_adj_5171, n144_adj_5172, n147_adj_5173, 
        n150_adj_5174, n153_adj_5175, n156_adj_5176, n159_adj_5177, 
        n162_adj_5178, n165_adj_5179, n168_adj_5180, n171_adj_5181, 
        n174_adj_5182, n177_adj_5183, n180_adj_5184, n183_adj_5185, 
        n33_adj_5186, n36_adj_5187, n39, n42, n45, n48, n51, n54, 
        n57, n60, n78_adj_5188, n81_adj_5189, n84_adj_5190, n87_adj_5191, 
        n90_adj_5192, n93_adj_5193, n96_adj_5194, n99_adj_5195, n102_adj_5196, 
        n105_adj_5197, n108_adj_5198, n111_adj_5199, n114_adj_5200, 
        n117_adj_5201, n120_adj_5202, n123_adj_5203, n126_adj_5204, 
        n129_adj_5205, n132_adj_5206, n135_adj_5207, n138_adj_5208, 
        n141_adj_5209, n144_adj_5210, n147_adj_5211, n150_adj_5212, 
        n153_adj_5213, n156_adj_5214, n159_adj_5215, n162_adj_5216, 
        n165_adj_5217, n168_adj_5218, n171_adj_5219, n174_adj_5220, 
        n177_adj_5221, n180_adj_5222, n183_adj_5223, n78_adj_5224, n81_adj_5225, 
        n84_adj_5226, n87_adj_5227, n90_adj_5228, n93_adj_5229, n96_adj_5230, 
        n99_adj_5231, n102_adj_5232, n105_adj_5233, n108_adj_5234, n111_adj_5235, 
        n114_adj_5236, n117_adj_5237, n120_adj_5238, n123_adj_5239, 
        n126_adj_5240, n129_adj_5241, n132_adj_5242, n135_adj_5243, 
        n138_adj_5244, n141_adj_5245, n144_adj_5246, n147_adj_5247, 
        n150_adj_5248, n153_adj_5249, n156_adj_5250, n159_adj_5251, 
        n162_adj_5252, n165_adj_5253, n168_adj_5254, n171_adj_5255, 
        n174_adj_5256, n177_adj_5257, n180_adj_5258, n183_adj_5259, 
        n78_adj_5260, n81_adj_5261, n84_adj_5262, n87_adj_5263, n90_adj_5264, 
        n93_adj_5265, n96_adj_5266, n99_adj_5267, n102_adj_5268, n105_adj_5269, 
        n108_adj_5270, n111_adj_5271, n114_adj_5272, n117_adj_5273, 
        n120_adj_5274, n45_adj_5275, n48_adj_5276, n51_adj_5277, n54_adj_5278, 
        n57_adj_5279, n60_adj_5280, n63_adj_5281, n66_adj_5282, n69, 
        n72, n75, n78_adj_5283, n81_adj_5284, n84_adj_5285, n87_adj_5286, 
        n90_adj_5287, cout_adj_5288, n78_adj_5289, n81_adj_5290, n84_adj_5291, 
        n87_adj_5292, n90_adj_5293, n93_adj_5294, n96_adj_5295, n99_adj_5296, 
        n102_adj_5297, n105_adj_5298, n108_adj_5299, n111_adj_5300, 
        n114_adj_5301, n117_adj_5302, n120_adj_5303, n123_adj_5304, 
        n126_adj_5305, n129_adj_5306, n132_adj_5307, n135_adj_5308, 
        n138_adj_5309, n141_adj_5310, n144_adj_5311, n147_adj_5312, 
        n150_adj_5313, n153_adj_5314, n156_adj_5315, n159_adj_5316, 
        n162_adj_5317, n165_adj_5318, n168_adj_5319, n171_adj_5320, 
        n174_adj_5321, n177_adj_5322, n180_adj_5323, n183_adj_5324, 
        cout_adj_5325, cout_adj_5326, cout_adj_5327, n36_adj_5328, n39_adj_5329, 
        n42_adj_5330, n45_adj_5331, n48_adj_5332, n51_adj_5333, n54_adj_5334, 
        n57_adj_5335, n60_adj_5336, n63_adj_5337, n66_adj_5338, n69_adj_5339, 
        n72_adj_5340, n75_adj_5341, n78_adj_5342, n81_adj_5343, cout_adj_5344, 
        cout_adj_5345, n45_adj_5346, n48_adj_5347, n51_adj_5348, n54_adj_5349, 
        n57_adj_5350, n60_adj_5351, n63_adj_5352, n66_adj_5353, n69_adj_5354, 
        n72_adj_5355, n75_adj_5356, n78_adj_5357, n81_adj_5358, n84_adj_5359, 
        n87_adj_5360, n90_adj_5361, cout_adj_5362, cout_adj_5363, n78_adj_5364, 
        n81_adj_5365, n84_adj_5366, n87_adj_5367, n90_adj_5368, n93_adj_5369, 
        n96_adj_5370, n99_adj_5371, n102_adj_5372, n105_adj_5373, n108_adj_5374, 
        n111_adj_5375, n114_adj_5376, n117_adj_5377, n120_adj_5378, 
        n123_adj_5379, n126_adj_5380, n129_adj_5381, n132_adj_5382, 
        n135_adj_5383, n138_adj_5384, n141_adj_5385, n144_adj_5386, 
        n147_adj_5387, n150_adj_5388, n153_adj_5389, n156_adj_5390, 
        n159_adj_5391, n162_adj_5392, n165_adj_5393, n168_adj_5394, 
        n171_adj_5395, n174_adj_5396, n177_adj_5397, n180_adj_5398, 
        n183_adj_5399, n36_adj_5400, n39_adj_5401, n42_adj_5402, n45_adj_5403, 
        n48_adj_5404, n51_adj_5405, n54_adj_5406, n57_adj_5407, n60_adj_5408, 
        n63_adj_5409, n66_adj_5410, n69_adj_5411, n72_adj_5412, n75_adj_5413, 
        n78_adj_5414, n81_adj_5415, n130, n133_adj_5416, n136_adj_5417, 
        n139, n142, n145, n148, n151, n154, n157, n160, n163, 
        n166, n169, n172, n175, n178, n181, n184, n187, n190, 
        n193, n196, n199, n202, n205, n208, n211, n214, n217, 
        n220, n223, n226, n229, n232, n235, n238, n241, n244, 
        n247, n250, n253, n256, n259, n262, n265, n268, n271, 
        n274, n277, n280, n283, n286, n289, n292, n295, n298, 
        n301, n304, n307, n310, n313, n316, n76, n79, n82, 
        n85, n88, n91, n94, n97, n100, n103, n106, n109, n112, 
        n115, n118, n54_adj_5418, n57_adj_5419, n60_adj_5420, n63_adj_5421, 
        n66_adj_5422, n69_adj_5423, n72_adj_5424, n75_adj_5425, n78_adj_5426, 
        n81_adj_5427, n84_adj_5428, n87_adj_5429, n90_adj_5430, n93_adj_5431, 
        n96_adj_5432, n99_adj_5433, n102_adj_5434, n105_adj_5435, n108_adj_5436, 
        n111_adj_5437, n114_adj_5438, n117_adj_5439, n120_adj_5440, 
        n123_adj_5441, n126_adj_5442, cout_adj_5443, n78_adj_5444, n81_adj_5445, 
        n84_adj_5446, n87_adj_5447, n90_adj_5448, n93_adj_5449, n96_adj_5450, 
        n99_adj_5451, n102_adj_5452, n105_adj_5453, n108_adj_5454, n111_adj_5455, 
        n114_adj_5456, n117_adj_5457, n120_adj_5458, n123_adj_5459, 
        n126_adj_5460, n129_adj_5461, n132_adj_5462, n135_adj_5463, 
        n138_adj_5464, n141_adj_5465, n144_adj_5466, n147_adj_5467, 
        n150_adj_5468, n153_adj_5469, n156_adj_5470, n159_adj_5471, 
        n162_adj_5472, n165_adj_5473, n168_adj_5474, n171_adj_5475, 
        n174_adj_5476, n177_adj_5477, n180_adj_5478, n183_adj_5479, 
        n78_adj_5480, n81_adj_5481, n84_adj_5482, n87_adj_5483, n90_adj_5484, 
        n93_adj_5485, n96_adj_5486, n99_adj_5487, n102_adj_5488, n105_adj_5489, 
        n108_adj_5490, n111_adj_5491, n114_adj_5492, n117_adj_5493, 
        n120_adj_5494, n123_adj_5495, n126_adj_5496, n129_adj_5497, 
        n132_adj_5498, n135_adj_5499, n138_adj_5500, n141_adj_5501, 
        n144_adj_5502, n147_adj_5503, n150_adj_5504, n153_adj_5505, 
        n156_adj_5506, n159_adj_5507, n162_adj_5508, n165_adj_5509, 
        n168_adj_5510, n171_adj_5511, n174_adj_5512, n177_adj_5513, 
        n180_adj_5514, n183_adj_5515, n16038, n16037, n16036, n16035, 
        n16034, n16033, n16032, n16031, n16030, n16029, n16028, 
        n16027, n16026, n16025, n16024, n16023, n16022, n16021, 
        n16020, n16019, n16018, n16017, n16016, n16015, n16014, 
        n16013, n16012, n16011, n16010, n16009, n16008, n16007, 
        n16006, n16005, n16004, n16003, cout_adj_5516, n16428, n16469, 
        n16427, n16468, n16426, n16314, n16467, n16425, n16466, 
        n17940, n16465, n16238, n16389, n16461, n16460, clk_80mhz_enable_1407, 
        cout_adj_5517, n16420, n16419, n16418, n16417, n16416, n16415, 
        n16414, n16313, n16312, n16311, n16310, n16309, n16308, 
        n16307, n12290, n12172, n12170, n12168, n12294, n12162, 
        n12160, n16172, n12156, n12152, n12150, n12148, n12146, 
        n12144, n12142, n12138, n12136, n12134, n12132, n12130, 
        n12128, n12126, n12124, n12122, n12120, n16171, n12116, 
        n12114, n12112, n12110, n12108, n12106, n12102, n12098, 
        n12094, n12092, n12086, n12084, n12082, n12078, n12076, 
        n16413, n17939, n17955, n15224, n16237, n16459, n16458, 
        n16404, n17094, n16457, n16456, n16306, n16305, n16455, 
        n16454, n16304, n45_adj_5518, n48_adj_5519, n51_adj_5520, 
        n54_adj_5521, n16412, n57_adj_5522, n60_adj_5523, n16453, 
        n63_adj_5524, n16394, n66_adj_5525, n16452, n69_adj_5526, 
        n72_adj_5527, n75_adj_5528, n16302, n78_adj_5529, n16393, 
        n81_adj_5530, n16451, n84_adj_5531, n87_adj_5532, n16450, 
        n90_adj_5533, n16301, n11804, n16449, n16448, n16236, n16300, 
        n16191, n16447, n16446, n16299, n16403, n16445, n16444, 
        n16218, n16442, n16298, n16441, n16392, n16440, n16297, 
        n16235, n16002, n16001, n16000, n15999, n15998, n15997, 
        n15996, n15995, n15994, n15993, n15992, n15991, n15990, 
        n15989, n15988, n15987, n15223, n15222, n16439, n16438, 
        n16437, n16436, n16391, n16234, n16435, n16434, n16296, 
        n16433, n16390, n16295, n17663, n15221, n16233, n16432, 
        n16431, n16294, n16293, n16292, n16291, n16290, n16289, 
        n16288, n16287, n16286, n16285, n16284, n16283, n16282, 
        n16281, n16280, n16279, n16222, n16278, n16277, n16276, 
        n16275, n16274, n16273, n16272, n16271, n16270, n16269, 
        n16268, n16267, n16266, n16265, n16411, n16264, n16173, 
        n16219, n16263, n16262, n16261, n16260, n16259, n16258, 
        n16257, n16256, n16255, n16254, n16253, n16252, n16251, 
        n16249, n16698, n15220, n16697, n16696, n16695, n16694, 
        n16693, n16692, n16691, n16690, cout_adj_5534, clk_80mhz_enable_1469, 
        n16684, clk_80mhz_enable_1471, n16683, n16682, n16681, n16680, 
        n15986, n16679, n16678, n16677, n16676, n15985, n16670, 
        n15984, n16669, n16668, n16667, n16666, n16665, n16664, 
        n16663, n45_adj_5535, n16410, n48_adj_5536, n17097, n51_adj_5537, 
        n54_adj_5538, n16409, n57_adj_5539, n60_adj_5540, n16408, 
        n63_adj_5541, n16657, n66_adj_5542, n69_adj_5543, n16656, 
        n72_adj_5544, n16407, n75_adj_5545, n16655, n78_adj_5546, 
        n81_adj_5547, n16232, n84_adj_5548, n16654, n87_adj_5549, 
        n16398, n90_adj_5550, n16653, n16231, n16652, n16651, n16650, 
        n16649, n16230, n16229, n16643, n16406, n16397, n16642, 
        n16641, n16640, n16639, n16228, n16638, n16637, n16396, 
        n16636, n16635, n16634, n16227, n16633, n16632, n16631, 
        n16395, n16630, n15219, n16629, n16430, n16429, n16628, 
        n16627, n15983, n15982, n15981, n15980, n15979, n15978, 
        n15977, n15976, n15975, n15974, n15973, n15972, n15971, 
        n15970, n15969, n15968, n15967, n15966, n15965, n15964, 
        n15963, n15962, n15961, n15960, n15959, n15958, n15957, 
        n15956, n15955, n15953, n15952, n15951, n15950, n15949, 
        n15948, n15947, n15946, n15945, n15944, n15943, n15942, 
        cout_adj_5551, n15941, n15940, n15939, n15938, n15937, n15936, 
        n15935, n15934, n15933, n15932, n15931, n15930, n15929, 
        n15928, n15927, n15926, n15925, n15924, n15923, n15921, 
        n15920, n15919, n15918, n15917, n15916, n15915, n15914, 
        n15913, n15912, n15911, n15910, n15909, n15908, n15907, 
        n15906, n15905, n15904, n15903, n15902, n15901, n15900, 
        n15899, n15898, n15897, n15896, n15895, n15894, n15893, 
        n15892, n15891, n15890, n15889, n15888, n15887, n15886, 
        n15885, n15884, n15883, n15882, n15881, n15880, n15879, 
        n15878, n15876, n15875, n15874, n15873, n15872, n15871, 
        n15870, n15869, n15868, n15867, n78_adj_5552, n15866, n81_adj_5553, 
        n15865, n84_adj_5554, n15864, n87_adj_5555, n15863, n90_adj_5556, 
        n15862, n93_adj_5557, n15861, n96_adj_5558, n15860, n99_adj_5559, 
        n15859, n102_adj_5560, n105_adj_5561, n108_adj_5562, n15855, 
        n111_adj_5563, n15854, n114_adj_5564, n15853, n117_adj_5565, 
        n15852, n120_adj_5566, n15851, n123_adj_5567, n15850, n126_adj_5568, 
        n15849, n129_adj_5569, n15848, n132_adj_5570, n15847, n135_adj_5571, 
        n15846, n138_adj_5572, n15845, n141_adj_5573, n15844, n144_adj_5574, 
        n15843, n147_adj_5575, n15842, n150_adj_5576, n15841, n153_adj_5577, 
        n15840, n156_adj_5578, n15839, n159_adj_5579, n15838, n162_adj_5580, 
        n165_adj_5581, n15836, n168_adj_5582, n15835, n171_adj_5583, 
        n15834, n174_adj_5584, n15833, n177_adj_5585, n15832, n180_adj_5586, 
        n15831, n183_adj_5587, n15830, n15829, n15828, n15827, n15826, 
        n15825, n15824, n15823, n15822, n15821, n15820, n15819, 
        n15815, n15814, n15813, n15812, n15811, n15810, n15809, 
        n15808, n15807, n15806, n15805, n15804, n15803, n15802, 
        n15801, n15800, n15799, n15798, n15797, n15796, n15795, 
        n15794, n15793, n15792, n15791, n15790, n15789, n15788, 
        n15787, n15786, n15785, n15784, n15783, n15782, n15781, 
        n15780, n15778, n15777, n15776, n15775, n15774, n15773, 
        n15772, n15771, n15770, n15769, n15768, n15767, n15766, 
        n15765, n15764, n15763, n15762, n15761, n15757, n15756, 
        n15755, n15754, n15753, n15752, n15751, n15750, n15749, 
        n15748, n15747, n15746, n15745, n15744, n15743, n15742, 
        n15741, n15740, n15738, n15737, n15736, n15735, n15734, 
        n15733, n15732, n15731, n15730, n15729, n15728, n15727, 
        n15726, n15725, n15724, n15723, n15722, n15721, n15720, 
        n15719, n15718, n15717, n15716, n15715, n15714, n15713, 
        n15712, n15711, n15710, n15709, n15708, n15706, n15705, 
        n15704, n15703, n15702, n15701, n15700, n15699, n15698, 
        n15697, n15696, n15695, n15694, n15693, n15692, n15691, 
        n15690, n15689, n15685, n15684, n15683, n15682, n15681, 
        n15680, n15679, n15678, n15677, n15676, n15675, n15674, 
        n15673, n15672, n15671, n15670, n15669, n15668, n15666, 
        n15665, n45_adj_5588, n15664, n48_adj_5589, n15663, n51_adj_5590, 
        n15662, n54_adj_5591, n15661, n57_adj_5592, n15660, n60_adj_5593, 
        n15659, n63_adj_5594, n15658, n66_adj_5595, n15657, n69_adj_5596, 
        n15656, n72_adj_5597, n15655, n75_adj_5598, n15654, n78_adj_5599, 
        n15653, n81_adj_5600, n15652, n84_adj_5601, n15651, n87_adj_5602, 
        n15650, n90_adj_5603, n15649, n15645, n15644, n15643, n15642, 
        n15641, n15640, n15639, n15638, n15637, n15636, n15635, 
        n15634, n15633, n15632, n15631, n15630, n15629, n15628, 
        n15627, n15626, n15625, n15624, n15623, n15622, n15621, 
        n15620, n15619, n15618, n15617, n15616, n15613, n41, n44, 
        n15612, n47, n15611, n50, n15610, n53, n15609, n56, 
        n15608, n59, n15607, n62, n15606, n65_adj_5604, n15605, 
        n68, n15604, n71, n15603, n74, n15602, n77, n15601, 
        n80, n15600, n15599, n15598, n15597, n15596, n15592, n15591, 
        n15590, n15589, n15588, n15587, n15586, n15585, n15584, 
        n15583, n15582, n15581, n15580, n15579, n15578, n15577, 
        n15576, n15575, n15573, n15572, n15571, n15570, n15569, 
        n15568, n15567, n15566, n15565, n15564, n15563, n15562, 
        n15561, n15560, n15559, n15558, n15557, n15556, n15552, 
        n15551, n15550, n15549, n15548, n15547, n15546, n15545, 
        n15544, n15543, n15542, n15541, n15540, n15539, n15538, 
        n15537, n15536, n15535, n15534, n15533, n15532, n15531, 
        n15530, n15529, n15527, n15526, n15525, n15524, n15523, 
        n15522, n15521, n15520, n15519, n15518, n15517, n15516, 
        n15515, n15514, n15513, n15512, n15511, n15510, n15505, 
        n15504, n15503, n15502, n15501, n15500, cout_adj_5605, n15499, 
        n15498, n15497, n15492, n15491, n15490, n15489, n15488, 
        n15487, n15486, n15485, n15484, n15483, n15482, n15481, 
        n15480, n15479, n15478, n15477, n15476, n15475, n15474, 
        n15473, n15472, n15471, n15470, n15469, n15468, n15467, 
        n15466, n15465, n15464, n15463, n15462, n15461, n15460, 
        n15459, n15458, n15457, n15456, n15455, n15454, n15453, 
        n15452, n15451, n15450, n15449, n15448, n15447, n15446, 
        n15445, n15444, n15443, n15442, n15441, n15440, n15439, 
        n15438, n15437, n15436, n15435, n15434, n15433, n15432, 
        n15431, n15430, n15429, n15428, n15427, n15426, n15425, 
        n15424, n15423, n15422, n15421, n15420, n15419, n15418, 
        n15417, n15416, n15415, n15414, n15413, n15412, n15411, 
        n15410, n15409, n15408, n15407, n15406, n15405, n15404, 
        n15403, n15402, n15401, n15400, n15399, n15398, n15397, 
        n15396, n15395, n15394, n15392, n15391, n15390, n15389, 
        n15388, n15387, n15386, n15385, n15384, n15383, n15382, 
        n15381, n15380, n15379, n15378, n15377, n15376, n15375, 
        n15374, n15373, n15372, n15371, n15370, n15369, n15368, 
        n15367, n15366, n15365, n15364, n15363, n15362, n15361, 
        n15360, n15359, n15358, n15357, n15354, n15353, n15352, 
        n15351, n15350, n15349, n15348, n15347, n15346, n15345, 
        n29_adj_5606, n32_adj_5607, n15344, n35_adj_5608, n15343, 
        n38, n15342, n41_adj_5609, n15341, n44_adj_5610, n15340, 
        n47_adj_5611, n15339, n50_adj_5612, n15338, n15337, n15332, 
        n15331, n15330, n15329, n15328, n15327, n15326, n15325, 
        n15324, n15323, n15322, n15321, n15320, n15319, n15318, 
        n15317, n15316, n15315, n15311, n15310, n15309, n15308, 
        n15307, n15306, n15305, n15304, n15303, n15302, n15301, 
        n15300, n15299, n15298, n15297, n15296, n15295, n15294, 
        n15292, n15291, n15290, n15289, n15288, n15287, n15286, 
        n15285, n15284, n15283, n15282, n15281, n15280, n16405, 
        n15279, n15278, n15277, n15276, n15275, n15274, n15273, 
        n15272, n15271, n15270, n15269, n15268, n15267, n15266, 
        n15265, n15264, n15263, n15262, n15261, n15260, n15259, 
        n15258, n15257, n15256, n15255, n15254, n15253, n15252, 
        n15251, n15250, n15249, n15248, n15247, n15246, n15245, 
        cout_adj_5613, n15244, n15243, n15242, n15241, n15240, n15239, 
        n15238, n15237, n15236, n15235, n15234, n15233, n15232, 
        n15231, n15230, n15229, n15228, n17205, n17925, clk_80mhz_enable_1459, 
        n37_adj_5614, n40, n18121, n43, n46, n49, n52, n55, 
        n58, n61, n64_adj_5615, n67, n70, n76_adj_5616, n79_adj_5617, 
        n82_adj_5618, n85_adj_5619, n88_adj_5620, n91_adj_5621, n94_adj_5622, 
        n97_adj_5623, n100_adj_5624, n103_adj_5625, n106_adj_5626, n109_adj_5627, 
        n112_adj_5628, n115_adj_5629, n118_adj_5630, n124, n127, n130_adj_5631, 
        n133_adj_5632, n136_adj_5633, n139_adj_5634, n142_adj_5635, 
        n145_adj_5636, n148_adj_5637, n151_adj_5638, n154_adj_5639, 
        n157_adj_5640, n160_adj_5641, n163_adj_5642, n166_adj_5643, 
        n169_adj_5644, n172_adj_5645, n175_adj_5646, n178_adj_5647, 
        n181_adj_5648, n184_adj_5649, n187_adj_5650, n190_adj_5651, 
        n193_adj_5652, n196_adj_5653, n199_adj_5654, n202_adj_5655, 
        n205_adj_5656, n208_adj_5657, n211_adj_5658, n214_adj_5659, 
        n217_adj_5660, n220_adj_5661, n223_adj_5662, n226_adj_5663, 
        n229_adj_5664, n232_adj_5665, n235_adj_5666, n238_adj_5667, 
        n241_adj_5668, n244_adj_5669, n247_adj_5670, n250_adj_5671, 
        n253_adj_5672, n256_adj_5673, n259_adj_5674, n262_adj_5675, 
        n265_adj_5676, n268_adj_5677, n271_adj_5678, n274_adj_5679, 
        n17777, n277_adj_5680, n280_adj_5681, n283_adj_5682, n286_adj_5683, 
        n289_adj_5684, n292_adj_5685, n295_adj_5686, n298_adj_5687, 
        n301_adj_5688, n17401, n15218, n15217, n15216, n15215, n17397, 
        n17610, n78_adj_5689, n81_adj_5690, n84_adj_5691, n87_adj_5692, 
        n90_adj_5693, n93_adj_5694, n96_adj_5695, n99_adj_5696, n102_adj_5697, 
        n105_adj_5698, n108_adj_5699, n111_adj_5700, n114_adj_5701, 
        n117_adj_5702, n120_adj_5703, n123_adj_5704, n126_adj_5705, 
        n129_adj_5706, n17938, n132_adj_5707, n135_adj_5708, n138_adj_5709, 
        n141_adj_5710, n144_adj_5711, n147_adj_5712, n150_adj_5713, 
        n153_adj_5714, n156_adj_5715, n159_adj_5716, n162_adj_5717, 
        n165_adj_5718, n168_adj_5719, n171_adj_5720, n174_adj_5721, 
        n177_adj_5722, n180_adj_5723, n183_adj_5724, n11_adj_5725, n13_adj_5726, 
        n17937, n17069, n15214, n15213, n15212, n27_adj_5727, n40_adj_5728, 
        n21_adj_5729, n15211, n15210, n15208, n15203, n15202, n17961, 
        n17960, n17317, n18075, clk_80mhz_enable_1470, n12983, n15173, 
        n15205, n15206, n29_adj_5730, n17959, n15198, n15201, n15200, 
        n15199, n15209, n17953, n17952, n15207, n15204, n17090, 
        n17934, n17933, n17954, n17932, n17906, n17905, n17951, 
        n17664, n18076;
    
    VHI i2 (.Z(VCC_net));
    \uart_rx(CLKS_PER_BIT=87)  uart_rx_inst (.clk_80mhz(clk_80mhz), .i_Rx_Serial_c(i_Rx_Serial_c), 
            .r_Rx_Data(r_Rx_Data), .o_Rx_Byte1({o_Rx_Byte1}), .\r_Rx_Byte[4] (r_Rx_Byte[4]), 
            .n17663(n17663), .GND_net(GND_net), .VCC_net(VCC_net), .o_Rx_DV1(o_Rx_DV1), 
            .n17943(n17943), .\r_Rx_Byte[6] (r_Rx_Byte[6]), .n17945(n17945), 
            .n17397(n17397), .n17946(n17946), .n17664(n17664)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(179[33] 184[5])
    CCU2C _add_1_1424_add_4_12 (.A0(d1_adj_5740[10]), .B0(MixerOutCos[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[11]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16308), .COUT(n16309), .S0(d1_71__N_418_adj_5756[10]), 
          .S1(d1_71__N_418_adj_5756[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_10 (.A0(d1_adj_5740[8]), .B0(MixerOutCos[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[9]), .B1(MixerOutCos[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16307), .COUT(n16308), .S0(d1_71__N_418_adj_5756[8]), 
          .S1(d1_71__N_418_adj_5756[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_10.INJECT1_1 = "NO";
    LUT4 i2354_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(n18076), .D(n169_adj_5644), 
         .Z(n12152)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2354_3_lut_4_lut.init = 16'hf808;
    CCU2C _add_1_1436_add_4_28 (.A0(d4_adj_5743[26]), .B0(d3_adj_5742[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[27]), .B1(d3_adj_5742[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16171), .COUT(n16172), .S0(d4_71__N_634_adj_5759[26]), 
          .S1(d4_71__N_634_adj_5759[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_28.INJECT1_1 = "NO";
    Mixer Mixer_inst (.MixerOutCos({MixerOutCos}), .clk_80mhz(clk_80mhz), 
          .MixerOutSin({MixerOutSin}), .DiffOut_c(DiffOut_c), .RFIn_c(RFIn_c), 
          .\LOCosine[10] (LOCosine[10]), .MixerOutCos_11__N_250({MixerOutCos_11__N_250}), 
          .\LOCosine[7] (LOCosine[7]), .\LOCosine[6] (LOCosine[6]), .\LOCosine[11] (LOCosine[11]), 
          .\LOCosine[5] (LOCosine[5]), .\LOCosine[4] (LOCosine[4]), .\LOCosine[3] (LOCosine[3]), 
          .\LOSine[1] (LOSine[1]), .MixerOutSin_11__N_236({MixerOutSin_11__N_236}), 
          .\LOCosine[2] (LOCosine[2]), .\LOCosine[12] (LOCosine[12]), .\LOCosine[1] (LOCosine[1]), 
          .\LOSine[12] (LOSine[12]), .\LOCosine[9] (LOCosine[9]), .\LOCosine[8] (LOCosine[8]), 
          .\LOSine[11] (LOSine[11]), .\LOSine[10] (LOSine[10]), .\LOSine[9] (LOSine[9]), 
          .\LOSine[8] (LOSine[8]), .\LOSine[7] (LOSine[7]), .\LOSine[6] (LOSine[6]), 
          .\LOSine[5] (LOSine[5]), .\LOSine[4] (LOSine[4]), .\LOSine[3] (LOSine[3]), 
          .\LOSine[2] (LOSine[2])) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(122[10] 130[5])
    CCU2C _add_1_1436_add_4_26 (.A0(d4_adj_5743[24]), .B0(d3_adj_5742[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[25]), .B1(d3_adj_5742[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16170), .COUT(n16171), .S0(d4_71__N_634_adj_5759[24]), 
          .S1(d4_71__N_634_adj_5759[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_26.INJECT1_1 = "NO";
    CCU2C add_3836_19 (.A0(d_out_d_11__N_1884[17]), .B0(n48_adj_5519), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n45_adj_5518), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16551), .S0(n45_adj_5535), 
          .S1(d_out_d_11__N_1886[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3836_19.INIT0 = 16'h9995;
    defparam add_3836_19.INIT1 = 16'h9995;
    defparam add_3836_19.INJECT1_0 = "NO";
    defparam add_3836_19.INJECT1_1 = "NO";
    FD1S3AX o_Rx_Byte_i1 (.D(o_Rx_Byte1[0]), .CK(clk_80mhz), .Q(led_c_0));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    CCU2C _add_1_1406_add_4_6 (.A0(d1[4]), .B0(MixerOutSin[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[5]), .B1(MixerOutSin[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16324), .COUT(n16325), .S0(d1_71__N_418[4]), 
          .S1(d1_71__N_418[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_4 (.A0(d1[2]), .B0(MixerOutSin[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[3]), .B1(MixerOutSin[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16323), .COUT(n16324), .S0(d1_71__N_418[2]), 
          .S1(d1_71__N_418[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_31 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n99_adj_5296), .D0(d1[64]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n96_adj_5295), .D1(d1[65]), .CIN(n16194), .COUT(n16195), 
          .S0(d1_71__N_418[64]), .S1(d1_71__N_418[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_31.INJECT1_1 = "NO";
    CCU2C add_3836_17 (.A0(d_out_d_11__N_1884[17]), .B0(n54_adj_5521), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n51_adj_5520), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16550), .COUT(n16551), .S0(n51_adj_5537), 
          .S1(n48_adj_5536));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3836_17.INIT0 = 16'h9995;
    defparam add_3836_17.INIT1 = 16'h9995;
    defparam add_3836_17.INJECT1_0 = "NO";
    defparam add_3836_17.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_25 (.A0(d7_adj_5747[58]), .B0(cout_adj_5613), 
          .C0(n117_adj_4965), .D0(n15_adj_4700), .A1(d7_adj_5747[59]), 
          .B1(cout_adj_5613), .C1(n114_adj_4964), .D1(n14_adj_4701), .CIN(n16213), 
          .COUT(n16214), .S0(d8_71__N_1603_adj_5774[58]), .S1(d8_71__N_1603_adj_5774[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_25.INJECT1_1 = "NO";
    FD1S3AX o_Rx_DV_40 (.D(o_Rx_DV1), .CK(clk_80mhz), .Q(o_Rx_DV));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam o_Rx_DV_40.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i0 (.D(phase_inc_carrGen[0]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i0.GSR = "ENABLED";
    CCU2C _add_1_1439_add_4_24 (.A0(d5_adj_5744[22]), .B0(d4_adj_5743[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[23]), .B1(d4_adj_5743[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16110), .COUT(n16111), .S0(d5_71__N_706_adj_5760[22]), 
          .S1(d5_71__N_706_adj_5760[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_24 (.A0(d4_adj_5743[22]), .B0(d3_adj_5742[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[23]), .B1(d3_adj_5742[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16169), .COUT(n16170), .S0(d4_71__N_634_adj_5759[22]), 
          .S1(d4_71__N_634_adj_5759[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_28 (.A0(d1_adj_5740[26]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[27]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16316), .COUT(n16317), .S0(d1_71__N_418_adj_5756[26]), 
          .S1(d1_71__N_418_adj_5756[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_22 (.A0(d4_adj_5743[20]), .B0(d3_adj_5742[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[21]), .B1(d3_adj_5742[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16168), .COUT(n16169), .S0(d4_71__N_634_adj_5759[20]), 
          .S1(d4_71__N_634_adj_5759[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_22.INJECT1_1 = "NO";
    PWM PWM_inst (.\DataInReg[0] (DataInReg[0]), .clk_80mhz(clk_80mhz), 
        .\DataInReg_11__N_1856[0] (DataInReg_11__N_1856[0]), .counter({counter}), 
        .GND_net(GND_net), .VCC_net(VCC_net), .\DataInReg[1] (DataInReg[1]), 
        .\DataInReg_11__N_1856[1] (DataInReg_11__N_1856[1]), .\DataInReg[2] (DataInReg[2]), 
        .\DataInReg_11__N_1856[2] (DataInReg_11__N_1856[2]), .\DataInReg[3] (DataInReg[3]), 
        .\DataInReg_11__N_1856[3] (DataInReg_11__N_1856[3]), .\DataInReg[4] (DataInReg[4]), 
        .\DataInReg_11__N_1856[4] (DataInReg_11__N_1856[4]), .\DataInReg[5] (DataInReg[5]), 
        .\DataInReg_11__N_1856[5] (DataInReg_11__N_1856[5]), .\DataInReg[6] (DataInReg[6]), 
        .\DataInReg_11__N_1856[6] (DataInReg_11__N_1856[6]), .\DataInReg[7] (DataInReg[7]), 
        .\DataInReg_11__N_1856[7] (DataInReg_11__N_1856[7]), .\DataInReg[8] (DataInReg[8]), 
        .\DataInReg_11__N_1856[8] (DataInReg_11__N_1856[8]), .\DataInReg[9] (DataInReg[9]), 
        .\DemodOut[9] (DemodOut[9])) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(156[8] 160[5])
    CCU2C _add_1_1436_add_4_20 (.A0(d4_adj_5743[18]), .B0(d3_adj_5742[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[19]), .B1(d3_adj_5742[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16167), .COUT(n16168), .S0(d4_71__N_634_adj_5759[18]), 
          .S1(d4_71__N_634_adj_5759[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_32 (.A0(d_d9[29]), .B0(d9[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[30]), .B1(d9[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16291), .COUT(n16292));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_22 (.A0(d5_adj_5744[20]), .B0(d4_adj_5743[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[21]), .B1(d4_adj_5743[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16109), .COUT(n16110), .S0(d5_71__N_706_adj_5760[20]), 
          .S1(d5_71__N_706_adj_5760[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_18 (.A0(d4_adj_5743[16]), .B0(d3_adj_5742[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[17]), .B1(d3_adj_5742[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16166), .COUT(n16167), .S0(d4_71__N_634_adj_5759[16]), 
          .S1(d4_71__N_634_adj_5759[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_4 (.A0(d_d7_adj_5748[37]), .B0(d7_adj_5747[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[38]), .B1(d7_adj_5747[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16118), .COUT(n16119), .S0(n180_adj_4986), 
          .S1(n177_adj_4985));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_28 (.A0(d_d9[25]), .B0(d9[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[26]), .B1(d9[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16289), .COUT(n16290));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_20 (.A0(d5_adj_5744[18]), .B0(d4_adj_5743[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[19]), .B1(d4_adj_5743[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16108), .COUT(n16109), .S0(d5_71__N_706_adj_5760[18]), 
          .S1(d5_71__N_706_adj_5760[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_23 (.A0(d7_adj_5747[56]), .B0(cout_adj_5613), 
          .C0(n123_adj_4967), .D0(n17_adj_4698), .A1(d7_adj_5747[57]), 
          .B1(cout_adj_5613), .C1(n120_adj_4966), .D1(n16_adj_4699), .CIN(n16212), 
          .COUT(n16213), .S0(d8_71__N_1603_adj_5774[56]), .S1(d8_71__N_1603_adj_5774[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_16 (.A0(d4_adj_5743[14]), .B0(d3_adj_5742[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[15]), .B1(d3_adj_5742[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16165), .COUT(n16166), .S0(d4_71__N_634_adj_5759[14]), 
          .S1(d4_71__N_634_adj_5759[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_34 (.A0(d3[67]), .B0(d2[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[68]), .B1(d2[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15893), .COUT(n15894), .S0(n90_adj_5556), .S1(n87_adj_5555));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_34.INJECT1_1 = "NO";
    FD1P3AX CICGain__i1 (.D(led_c_0), .SP(clk_80mhz_enable_1407), .CK(clk_80mhz), 
            .Q(CICGain[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam CICGain__i1.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i1 (.D(n126_adj_5442), .CK(CIC1_out_clkSin), .Q(ISquare[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i1.GSR = "ENABLED";
    CCU2C _add_1_1424_add_4_8 (.A0(d1_adj_5740[6]), .B0(MixerOutCos[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[7]), .B1(MixerOutCos[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16306), .COUT(n16307), .S0(d1_71__N_418_adj_5756[6]), 
          .S1(d1_71__N_418_adj_5756[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_2 (.A0(d1[0]), .B0(MixerOutSin[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[1]), .B1(MixerOutSin[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16323), .S1(d1_71__N_418[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1406_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_3 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n183_adj_5324), .D0(d1[36]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n180_adj_5323), .D1(d1[37]), .CIN(n16180), .COUT(n16181), 
          .S0(d1_71__N_418[36]), .S1(d1_71__N_418[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_32 (.A0(d3[65]), .B0(d2[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[66]), .B1(d2[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15892), .COUT(n15893), .S0(n96_adj_5558), .S1(n93_adj_5557));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_26 (.A0(d1_adj_5740[24]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[25]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16315), .COUT(n16316), .S0(d1_71__N_418_adj_5756[24]), 
          .S1(d1_71__N_418_adj_5756[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_30 (.A0(d3[63]), .B0(d2[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[64]), .B1(d2[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15891), .COUT(n15892), .S0(n102_adj_5560), .S1(n99_adj_5559));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_24 (.A0(d1_adj_5740[22]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[23]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16314), .COUT(n16315), .S0(d1_71__N_418_adj_5756[22]), 
          .S1(d1_71__N_418_adj_5756[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_22 (.A0(d1_adj_5740[20]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[21]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16313), .COUT(n16314), .S0(d1_71__N_418_adj_5756[20]), 
          .S1(d1_71__N_418_adj_5756[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_20 (.A0(d1_adj_5740[18]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[19]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16312), .COUT(n16313), .S0(d1_71__N_418_adj_5756[18]), 
          .S1(d1_71__N_418_adj_5756[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_18 (.A0(d1_adj_5740[16]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[17]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16311), .COUT(n16312), .S0(d1_71__N_418_adj_5756[16]), 
          .S1(d1_71__N_418_adj_5756[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_21 (.A0(d7_adj_5747[54]), .B0(cout_adj_5613), 
          .C0(n129_adj_4969), .D0(n19_adj_4696), .A1(d7_adj_5747[55]), 
          .B1(cout_adj_5613), .C1(n126_adj_4968), .D1(n18_adj_4697), .CIN(n16211), 
          .COUT(n16212), .S0(d8_71__N_1603_adj_5774[54]), .S1(d8_71__N_1603_adj_5774[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_14 (.A0(d4_adj_5743[12]), .B0(d3_adj_5742[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[13]), .B1(d3_adj_5742[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16164), .COUT(n16165), .S0(d4_71__N_634_adj_5759[12]), 
          .S1(d4_71__N_634_adj_5759[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_12 (.A0(d4_adj_5743[10]), .B0(d3_adj_5742[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[11]), .B1(d3_adj_5742[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16163), .COUT(n16164), .S0(d4_71__N_634_adj_5759[10]), 
          .S1(d4_71__N_634_adj_5759[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_10 (.A0(d4_adj_5743[8]), .B0(d3_adj_5742[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[9]), .B1(d3_adj_5742[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16162), .COUT(n16163), .S0(d4_71__N_634_adj_5759[8]), 
          .S1(d4_71__N_634_adj_5759[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_19 (.A0(d7_adj_5747[52]), .B0(cout_adj_5613), 
          .C0(n135_adj_4971), .D0(n21_adj_4694), .A1(d7_adj_5747[53]), 
          .B1(cout_adj_5613), .C1(n132_adj_4970), .D1(n20_adj_4695), .CIN(n16210), 
          .COUT(n16211), .S0(d8_71__N_1603_adj_5774[52]), .S1(d8_71__N_1603_adj_5774[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_19.INJECT1_1 = "NO";
    LUT4 mux_325_i33_4_lut (.A(n12124), .B(n223), .C(n17925), .D(n2572), 
         .Z(n2339)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i33_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1424_add_4_16 (.A0(d1_adj_5740[14]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[15]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16310), .COUT(n16311), .S0(d1_71__N_418_adj_5756[14]), 
          .S1(d1_71__N_418_adj_5756[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_14 (.A0(d1_adj_5740[12]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[13]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16309), .COUT(n16310), .S0(d1_71__N_418_adj_5756[12]), 
          .S1(d1_71__N_418_adj_5756[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_14.INJECT1_1 = "NO";
    CCU2C add_3836_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1884[17]), .C0(n60_adj_5523), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n57_adj_5522), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16549), .COUT(n16550), .S0(n57_adj_5539), 
          .S1(n54_adj_5538));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3836_15.INIT0 = 16'h6969;
    defparam add_3836_15.INIT1 = 16'h9995;
    defparam add_3836_15.INJECT1_0 = "NO";
    defparam add_3836_15.INJECT1_1 = "NO";
    CCU2C add_3836_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1884[17]), .C0(n66_adj_5525), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1884[17]), 
          .C1(n63_adj_5524), .D1(VCC_net), .CIN(n16548), .COUT(n16549), 
          .S0(n63_adj_5541), .S1(n60_adj_5540));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3836_13.INIT0 = 16'h6969;
    defparam add_3836_13.INIT1 = 16'h6969;
    defparam add_3836_13.INJECT1_0 = "NO";
    defparam add_3836_13.INJECT1_1 = "NO";
    CCU2C add_3836_11 (.A0(d_out_d_11__N_1884[17]), .B0(n17938), .C0(n72_adj_5527), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n69_adj_5526), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16547), .COUT(n16548), .S0(n69_adj_5543), 
          .S1(n66_adj_5542));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3836_11.INIT0 = 16'h6969;
    defparam add_3836_11.INIT1 = 16'h9995;
    defparam add_3836_11.INJECT1_0 = "NO";
    defparam add_3836_11.INJECT1_1 = "NO";
    CCU2C add_3836_9 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(n78_adj_5529), .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), 
          .B1(d_out_d_11__N_1884[17]), .C1(n75_adj_5528), .D1(VCC_net), 
          .CIN(n16546), .COUT(n16547), .S0(n75_adj_5545), .S1(n72_adj_5544));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3836_9.INIT0 = 16'h9696;
    defparam add_3836_9.INIT1 = 16'h9696;
    defparam add_3836_9.INJECT1_0 = "NO";
    defparam add_3836_9.INJECT1_1 = "NO";
    CCU2C add_3836_7 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1884[17]), 
          .C0(n84_adj_5531), .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(d_out_d_11__N_1884[17]), .C1(n81_adj_5530), .D1(VCC_net), 
          .CIN(n16545), .COUT(n16546), .S0(n81_adj_5547), .S1(n78_adj_5546));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3836_7.INIT0 = 16'h9696;
    defparam add_3836_7.INIT1 = 16'h9696;
    defparam add_3836_7.INJECT1_0 = "NO";
    defparam add_3836_7.INJECT1_1 = "NO";
    CCU2C add_3836_5 (.A0(n90_adj_5533), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1882[17]), .B1(d_out_d_11__N_1884[17]), .C1(n87_adj_5532), 
          .D1(VCC_net), .CIN(n16544), .COUT(n16545), .S0(n87_adj_5549), 
          .S1(n84_adj_5548));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3836_5.INIT0 = 16'haaa0;
    defparam add_3836_5.INIT1 = 16'h9696;
    defparam add_3836_5.INJECT1_0 = "NO";
    defparam add_3836_5.INJECT1_1 = "NO";
    CCU2C add_3836_3 (.A0(d_out_d_11__N_1884[17]), .B0(ISquare[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16543), .COUT(n16544), .S1(n90_adj_5550));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3836_3.INIT0 = 16'h666a;
    defparam add_3836_3.INIT1 = 16'h555f;
    defparam add_3836_3.INJECT1_0 = "NO";
    defparam add_3836_3.INJECT1_1 = "NO";
    CCU2C add_3836_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1884[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16543));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3836_1.INIT0 = 16'h0000;
    defparam add_3836_1.INIT1 = 16'haaaf;
    defparam add_3836_1.INJECT1_0 = "NO";
    defparam add_3836_1.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_17 (.A0(d7_adj_5747[50]), .B0(cout_adj_5613), 
          .C0(n141_adj_4973), .D0(n23_adj_4692), .A1(d7_adj_5747[51]), 
          .B1(cout_adj_5613), .C1(n138_adj_4972), .D1(n22_adj_4693), .CIN(n16209), 
          .COUT(n16210), .S0(d8_71__N_1603_adj_5774[50]), .S1(d8_71__N_1603_adj_5774[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_2 (.A0(d1_adj_5740[0]), .B0(MixerOutCos[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[1]), .B1(MixerOutCos[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16304), .S1(d1_71__N_418_adj_5756[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1424_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_34 (.A0(d1[32]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[33]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16338), .COUT(n16339), .S0(d1_71__N_418[32]), 
          .S1(d1_71__N_418[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_8 (.A0(d4_adj_5743[6]), .B0(d3_adj_5742[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[7]), .B1(d3_adj_5742[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16161), .COUT(n16162), .S0(d4_71__N_634_adj_5759[6]), 
          .S1(d4_71__N_634_adj_5759[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_18 (.A0(d5_adj_5744[16]), .B0(d4_adj_5743[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[17]), .B1(d4_adj_5743[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16107), .COUT(n16108), .S0(d5_71__N_706_adj_5760[16]), 
          .S1(d5_71__N_706_adj_5760[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_29 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n105_adj_5298), .D0(d1[62]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n102_adj_5297), .D1(d1[63]), .CIN(n16193), .COUT(n16194), 
          .S0(d1_71__N_418[62]), .S1(d1_71__N_418[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_15 (.A0(d7_adj_5747[48]), .B0(cout_adj_5613), 
          .C0(n147_adj_4975), .D0(n25_adj_4690), .A1(d7_adj_5747[49]), 
          .B1(cout_adj_5613), .C1(n144_adj_4974), .D1(n24_adj_4691), .CIN(n16208), 
          .COUT(n16209), .S0(d8_71__N_1603_adj_5774[48]), .S1(d8_71__N_1603_adj_5774[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_27 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n111_adj_5300), .D0(d1[60]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n108_adj_5299), .D1(d1[61]), .CIN(n16192), .COUT(n16193), 
          .S0(d1_71__N_418[60]), .S1(d1_71__N_418[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_22 (.A0(d_d9[19]), .B0(d9[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[20]), .B1(d9[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16286), .COUT(n16287));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_6 (.A0(d4_adj_5743[4]), .B0(d3_adj_5742[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[5]), .B1(d3_adj_5742[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16160), .COUT(n16161), .S0(d4_71__N_634_adj_5759[4]), 
          .S1(d4_71__N_634_adj_5759[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_20 (.A0(d_d9[17]), .B0(d9[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[18]), .B1(d9[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16285), .COUT(n16286));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_14 (.A0(d_d9[11]), .B0(d9[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[12]), .B1(d9[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16282), .COUT(n16283));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_8 (.A0(d_d9[5]), .B0(d9[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[6]), .B1(d9[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16279), .COUT(n16280));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_13 (.A0(d7_adj_5747[46]), .B0(cout_adj_5613), 
          .C0(n153_adj_4977), .D0(n27_adj_4688), .A1(d7_adj_5747[47]), 
          .B1(cout_adj_5613), .C1(n150_adj_4976), .D1(n26_adj_4689), .CIN(n16207), 
          .COUT(n16208), .S0(d8_71__N_1603_adj_5774[46]), .S1(d8_71__N_1603_adj_5774[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_12 (.A0(d_d9[9]), .B0(d9[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[10]), .B1(d9[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16281), .COUT(n16282));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_18 (.A0(d_d9[15]), .B0(d9[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[16]), .B1(d9[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16284), .COUT(n16285));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_10 (.A0(d_d9[7]), .B0(d9[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[8]), .B1(d9[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16280), .COUT(n16281));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_6 (.A0(d_d9[3]), .B0(d9[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[4]), .B1(d9[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16278), .COUT(n16279));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_16 (.A0(d_d9[13]), .B0(d9[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[14]), .B1(d9[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16283), .COUT(n16284));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_28 (.A0(d3[61]), .B0(d2[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[62]), .B1(d2[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15890), .COUT(n15891), .S0(n108_adj_5562), .S1(n105_adj_5561));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_26 (.A0(d3[59]), .B0(d2[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[60]), .B1(d2[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15889), .COUT(n15890), .S0(n114_adj_5564), .S1(n111_adj_5563));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_24 (.A0(d3[57]), .B0(d2[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[58]), .B1(d2[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15888), .COUT(n15889), .S0(n120_adj_5566), .S1(n117_adj_5565));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_22 (.A0(d3[55]), .B0(d2[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[56]), .B1(d2[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15887), .COUT(n15888), .S0(n126_adj_5568), .S1(n123_adj_5567));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_20 (.A0(d3[53]), .B0(d2[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[54]), .B1(d2[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15886), .COUT(n15887), .S0(n132_adj_5570), .S1(n129_adj_5569));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_18 (.A0(d3[51]), .B0(d2[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[52]), .B1(d2[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15885), .COUT(n15886), .S0(n138_adj_5572), .S1(n135_adj_5571));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_11 (.A0(d7_adj_5747[44]), .B0(cout_adj_5613), 
          .C0(n159_adj_4979), .D0(n29_adj_4686), .A1(d7_adj_5747[45]), 
          .B1(cout_adj_5613), .C1(n156_adj_4978), .D1(n28_adj_4687), .CIN(n16206), 
          .COUT(n16207), .S0(d8_71__N_1603_adj_5774[44]), .S1(d8_71__N_1603_adj_5774[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_16 (.A0(d3[49]), .B0(d2[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[50]), .B1(d2[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15884), .COUT(n15885), .S0(n144_adj_5574), .S1(n141_adj_5573));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_14 (.A0(d3[47]), .B0(d2[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[48]), .B1(d2[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15883), .COUT(n15884), .S0(n150_adj_5576), .S1(n147_adj_5575));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_22 (.A0(d_d_tmp[19]), .B0(d_tmp[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[20]), .B1(d_tmp[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16268), .COUT(n16269), .S0(d6_71__N_1459[19]), 
          .S1(d6_71__N_1459[20]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_16 (.A0(d5_adj_5744[14]), .B0(d4_adj_5743[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[15]), .B1(d4_adj_5743[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16106), .COUT(n16107), .S0(d5_71__N_706_adj_5760[14]), 
          .S1(d5_71__N_706_adj_5760[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_24 (.A0(d_d9[21]), .B0(d9[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[22]), .B1(d9[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16287), .COUT(n16288));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_25 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n117_adj_5302), .D0(d1[58]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n114_adj_5301), .D1(d1[59]), .CIN(n16191), .COUT(n16192), 
          .S0(d1_71__N_418[58]), .S1(d1_71__N_418[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_4 (.A0(d_d9[1]), .B0(d9[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[2]), .B1(d9[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16277), .COUT(n16278));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[0]), .B1(d9[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16277));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1627_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_38 (.A0(d_d_tmp[35]), .B0(d_tmp[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16276), .S0(d6_71__N_1459[35]), .S1(cout_adj_5551));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1531_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_23 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n123_adj_5304), .D0(d1[56]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n120_adj_5303), .D1(d1[57]), .CIN(n16190), .COUT(n16191), 
          .S0(d1_71__N_418[56]), .S1(d1_71__N_418[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_36 (.A0(d_d_tmp[33]), .B0(d_tmp[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[34]), .B1(d_tmp[34]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16275), .COUT(n16276), .S0(d6_71__N_1459[33]), 
          .S1(d6_71__N_1459[34]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_32 (.A0(d_d_tmp[29]), .B0(d_tmp[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[30]), .B1(d_tmp[30]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16273), .COUT(n16274), .S0(d6_71__N_1459[29]), 
          .S1(d6_71__N_1459[30]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_32.INJECT1_1 = "NO";
    LUT4 mux_325_i34_4_lut (.A(n12126), .B(n220), .C(n17925), .D(n2572), 
         .Z(n2338)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i34_4_lut.init = 16'hcfca;
    CCU2C _add_1_1531_add_4_34 (.A0(d_d_tmp[31]), .B0(d_tmp[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[32]), .B1(d_tmp[32]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16274), .COUT(n16275), .S0(d6_71__N_1459[31]), 
          .S1(d6_71__N_1459[32]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_9 (.A0(d7_adj_5747[42]), .B0(cout_adj_5613), 
          .C0(n165_adj_4981), .D0(n31_adj_4683), .A1(d7_adj_5747[43]), 
          .B1(cout_adj_5613), .C1(n162_adj_4980), .D1(n30_adj_4685), .CIN(n16205), 
          .COUT(n16206), .S0(d8_71__N_1603_adj_5774[42]), .S1(d8_71__N_1603_adj_5774[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_9.INJECT1_1 = "NO";
    LUT4 i2372_3_lut_4_lut (.A(n18075), .B(n17937), .C(n18076), .D(n136_adj_5633), 
         .Z(n12170)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2372_3_lut_4_lut.init = 16'hfb0b;
    CCU2C _add_1_1436_add_4_4 (.A0(d4_adj_5743[2]), .B0(d3_adj_5742[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[3]), .B1(d3_adj_5742[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16159), .COUT(n16160), .S0(d4_71__N_634_adj_5759[2]), 
          .S1(d4_71__N_634_adj_5759[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_12 (.A0(d3[45]), .B0(d2[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[46]), .B1(d2[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15882), .COUT(n15883), .S0(n156_adj_5578), .S1(n153_adj_5577));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_10 (.A0(d3[43]), .B0(d2[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[44]), .B1(d2[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15881), .COUT(n15882), .S0(n162_adj_5580), .S1(n159_adj_5579));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_36 (.A0(d_d9[33]), .B0(d9[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[34]), .B1(d9[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16293), .COUT(n16294));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_13 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n153_adj_5314), .D0(d1[46]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n150_adj_5313), .D1(d1[47]), .CIN(n16185), .COUT(n16186), 
          .S0(d1_71__N_418[46]), .S1(d1_71__N_418[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_2 (.A0(d4_adj_5743[0]), .B0(d3_adj_5742[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[1]), .B1(d3_adj_5742[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16159), .S1(d4_71__N_634_adj_5759[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1436_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_6 (.A0(d1_adj_5740[4]), .B0(MixerOutCos[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[5]), .B1(MixerOutCos[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16305), .COUT(n16306), .S0(d1_71__N_418_adj_5756[4]), 
          .S1(d1_71__N_418_adj_5756[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_6.INJECT1_1 = "NO";
    FD1S3AX phase_accum_e3_i0_i0 (.D(n321), .CK(clk_80mhz), .Q(phase_accum_adj_5732[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i0.GSR = "ENABLED";
    CCU2C _add_1_1531_add_4_30 (.A0(d_d_tmp[27]), .B0(d_tmp[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[28]), .B1(d_tmp[28]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16272), .COUT(n16273), .S0(d6_71__N_1459[27]), 
          .S1(d6_71__N_1459[28]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_8 (.A0(d3[41]), .B0(d2[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[42]), .B1(d2[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15880), .COUT(n15881), .S0(n168_adj_5582), .S1(n165_adj_5581));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_37 (.A0(d6_adj_5745[70]), .B0(cout_adj_4625), 
          .C0(n81_adj_4917), .D0(n3), .A1(d6_adj_5745[71]), .B1(cout_adj_4625), 
          .C1(n78_adj_4916), .D1(n2), .CIN(n16156), .S0(d7_71__N_1531_adj_5773[70]), 
          .S1(d7_71__N_1531_adj_5773[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_35 (.A0(d6_adj_5745[68]), .B0(cout_adj_4625), 
          .C0(n87_adj_4919), .D0(n5), .A1(d6_adj_5745[69]), .B1(cout_adj_4625), 
          .C1(n84_adj_4918), .D1(n4), .CIN(n16155), .COUT(n16156), .S0(d7_71__N_1531_adj_5773[68]), 
          .S1(d7_71__N_1531_adj_5773[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_4 (.A0(d1_adj_5740[2]), .B0(MixerOutCos[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[3]), .B1(MixerOutCos[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16304), .COUT(n16305), .S0(d1_71__N_418_adj_5756[2]), 
          .S1(d1_71__N_418_adj_5756[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_33 (.A0(d6_adj_5745[66]), .B0(cout_adj_4625), 
          .C0(n93_adj_4921), .D0(n7), .A1(d6_adj_5745[67]), .B1(cout_adj_4625), 
          .C1(n90_adj_4920), .D1(n6), .CIN(n16154), .COUT(n16155), .S0(d7_71__N_1531_adj_5773[66]), 
          .S1(d7_71__N_1531_adj_5773[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_31 (.A0(d6_adj_5745[64]), .B0(cout_adj_4625), 
          .C0(n99_adj_4923), .D0(n9_adj_4741), .A1(d6_adj_5745[65]), .B1(cout_adj_4625), 
          .C1(n96_adj_4922), .D1(n8_adj_4745), .CIN(n16153), .COUT(n16154), 
          .S0(d7_71__N_1531_adj_5773[64]), .S1(d7_71__N_1531_adj_5773[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_8 (.A0(d_d_tmp[5]), .B0(d_tmp[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[6]), .B1(d_tmp[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16261), .COUT(n16262), .S0(d6_71__N_1459[5]), 
          .S1(d6_71__N_1459[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_20 (.A0(d_d_tmp[17]), .B0(d_tmp[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[18]), .B1(d_tmp[18]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16267), .COUT(n16268), .S0(d6_71__N_1459[17]), 
          .S1(d6_71__N_1459[18]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_4 (.A0(d_d_tmp[1]), .B0(d_tmp[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[2]), .B1(d_tmp[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16259), .COUT(n16260), .S0(d6_71__N_1459[1]), 
          .S1(d6_71__N_1459[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_6 (.A0(d3[39]), .B0(d2[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[40]), .B1(d2[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15879), .COUT(n15880), .S0(n174_adj_5584), .S1(n171_adj_5583));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_29 (.A0(d6_adj_5745[62]), .B0(cout_adj_4625), 
          .C0(n105_adj_4925), .D0(n11_adj_4743), .A1(d6_adj_5745[63]), 
          .B1(cout_adj_4625), .C1(n102_adj_4924), .D1(n10_adj_4742), .CIN(n16152), 
          .COUT(n16153), .S0(d7_71__N_1531_adj_5773[62]), .S1(d7_71__N_1531_adj_5773[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_27 (.A0(d6_adj_5745[60]), .B0(cout_adj_4625), 
          .C0(n111_adj_4927), .D0(n13_adj_4740), .A1(d6_adj_5745[61]), 
          .B1(cout_adj_4625), .C1(n108_adj_4926), .D1(n12_adj_4744), .CIN(n16151), 
          .COUT(n16152), .S0(d7_71__N_1531_adj_5773[60]), .S1(d7_71__N_1531_adj_5773[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_25 (.A0(d6_adj_5745[58]), .B0(cout_adj_4625), 
          .C0(n117_adj_4929), .D0(n15_adj_4738), .A1(d6_adj_5745[59]), 
          .B1(cout_adj_4625), .C1(n114_adj_4928), .D1(n14_adj_4739), .CIN(n16150), 
          .COUT(n16151), .S0(d7_71__N_1531_adj_5773[58]), .S1(d7_71__N_1531_adj_5773[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_23 (.A0(d6_adj_5745[56]), .B0(cout_adj_4625), 
          .C0(n123_adj_4931), .D0(n17_adj_4736), .A1(d6_adj_5745[57]), 
          .B1(cout_adj_4625), .C1(n120_adj_4930), .D1(n16_adj_4737), .CIN(n16149), 
          .COUT(n16150), .S0(d7_71__N_1531_adj_5773[56]), .S1(d7_71__N_1531_adj_5773[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_21 (.A0(d6_adj_5745[54]), .B0(cout_adj_4625), 
          .C0(n129_adj_4933), .D0(n19_adj_4734), .A1(d6_adj_5745[55]), 
          .B1(cout_adj_4625), .C1(n126_adj_4932), .D1(n18_adj_4735), .CIN(n16148), 
          .COUT(n16149), .S0(d7_71__N_1531_adj_5773[54]), .S1(d7_71__N_1531_adj_5773[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_19 (.A0(d6_adj_5745[52]), .B0(cout_adj_4625), 
          .C0(n135_adj_4935), .D0(n21_adj_4732), .A1(d6_adj_5745[53]), 
          .B1(cout_adj_4625), .C1(n132_adj_4934), .D1(n20_adj_4733), .CIN(n16147), 
          .COUT(n16148), .S0(d7_71__N_1531_adj_5773[52]), .S1(d7_71__N_1531_adj_5773[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_17 (.A0(d6_adj_5745[50]), .B0(cout_adj_4625), 
          .C0(n141_adj_4937), .D0(n23_adj_4730), .A1(d6_adj_5745[51]), 
          .B1(cout_adj_4625), .C1(n138_adj_4936), .D1(n22_adj_4731), .CIN(n16146), 
          .COUT(n16147), .S0(d7_71__N_1531_adj_5773[50]), .S1(d7_71__N_1531_adj_5773[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_15 (.A0(d6_adj_5745[48]), .B0(cout_adj_4625), 
          .C0(n147_adj_4939), .D0(n25_adj_4728), .A1(d6_adj_5745[49]), 
          .B1(cout_adj_4625), .C1(n144_adj_4938), .D1(n24_adj_4729), .CIN(n16145), 
          .COUT(n16146), .S0(d7_71__N_1531_adj_5773[48]), .S1(d7_71__N_1531_adj_5773[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_13 (.A0(d6_adj_5745[46]), .B0(cout_adj_4625), 
          .C0(n153_adj_4941), .D0(n27_adj_4726), .A1(d6_adj_5745[47]), 
          .B1(cout_adj_4625), .C1(n150_adj_4940), .D1(n26_adj_4727), .CIN(n16144), 
          .COUT(n16145), .S0(d7_71__N_1531_adj_5773[46]), .S1(d7_71__N_1531_adj_5773[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_11 (.A0(d6_adj_5745[44]), .B0(cout_adj_4625), 
          .C0(n159_adj_4943), .D0(n29_adj_4724), .A1(d6_adj_5745[45]), 
          .B1(cout_adj_4625), .C1(n156_adj_4942), .D1(n28_adj_4725), .CIN(n16143), 
          .COUT(n16144), .S0(d7_71__N_1531_adj_5773[44]), .S1(d7_71__N_1531_adj_5773[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[0]), .B1(d_tmp[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16259), .S1(d6_71__N_1459[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1531_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_9 (.A0(d6_adj_5745[42]), .B0(cout_adj_4625), 
          .C0(n165_adj_4945), .D0(n31_adj_4722), .A1(d6_adj_5745[43]), 
          .B1(cout_adj_4625), .C1(n162_adj_4944), .D1(n30_adj_4723), .CIN(n16142), 
          .COUT(n16143), .S0(d7_71__N_1531_adj_5773[42]), .S1(d7_71__N_1531_adj_5773[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_32 (.A0(d2_adj_5741[30]), .B0(d1_adj_5740[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[31]), .B1(d1_adj_5740[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16255), .COUT(n16256), .S0(d2_71__N_490_adj_5757[30]), 
          .S1(d2_71__N_490_adj_5757[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_8 (.A0(d2_adj_5741[6]), .B0(d1_adj_5740[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[7]), .B1(d1_adj_5740[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16243), .COUT(n16244), .S0(d2_71__N_490_adj_5757[6]), 
          .S1(d2_71__N_490_adj_5757[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_20 (.A0(d2_adj_5741[18]), .B0(d1_adj_5740[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[19]), .B1(d1_adj_5740[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16249), .COUT(n16250), .S0(d2_71__N_490_adj_5757[18]), 
          .S1(d2_71__N_490_adj_5757[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_2 (.A0(d2_adj_5741[0]), .B0(d1_adj_5740[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[1]), .B1(d1_adj_5740[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16241), .S1(d2_71__N_490_adj_5757[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1430_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_18 (.A0(d2_adj_5741[16]), .B0(d1_adj_5740[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[17]), .B1(d1_adj_5740[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16248), .COUT(n16249), .S0(d2_71__N_490_adj_5757[16]), 
          .S1(d2_71__N_490_adj_5757[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_30 (.A0(d2_adj_5741[28]), .B0(d1_adj_5740[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[29]), .B1(d1_adj_5740[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16254), .COUT(n16255), .S0(d2_71__N_490_adj_5757[28]), 
          .S1(d2_71__N_490_adj_5757[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_4 (.A0(d3[37]), .B0(d2[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[38]), .B1(d2[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15878), .COUT(n15879), .S0(n180_adj_5586), .S1(n177_adj_5585));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_4 (.A0(d2_adj_5741[2]), .B0(d1_adj_5740[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[3]), .B1(d1_adj_5740[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16241), .COUT(n16242), .S0(d2_71__N_490_adj_5757[2]), 
          .S1(d2_71__N_490_adj_5757[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_16 (.A0(d2_adj_5741[14]), .B0(d1_adj_5740[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[15]), .B1(d1_adj_5740[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16247), .COUT(n16248), .S0(d2_71__N_490_adj_5757[14]), 
          .S1(d2_71__N_490_adj_5757[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_28 (.A0(d2_adj_5741[26]), .B0(d1_adj_5740[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[27]), .B1(d1_adj_5740[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16253), .COUT(n16254), .S0(d2_71__N_490_adj_5757[26]), 
          .S1(d2_71__N_490_adj_5757[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_28.INJECT1_1 = "NO";
    LUT4 mux_325_i31_4_lut (.A(n12120), .B(n229), .C(n17925), .D(n2572), 
         .Z(n2341)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i31_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1430_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16258), .S0(cout_adj_5344));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1430_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1430_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_12 (.A0(d2_adj_5741[10]), .B0(d1_adj_5740[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[11]), .B1(d1_adj_5740[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16245), .COUT(n16246), .S0(d2_71__N_490_adj_5757[10]), 
          .S1(d2_71__N_490_adj_5757[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_26 (.A0(d2_adj_5741[24]), .B0(d1_adj_5740[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[25]), .B1(d1_adj_5740[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16252), .COUT(n16253), .S0(d2_71__N_490_adj_5757[24]), 
          .S1(d2_71__N_490_adj_5757[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_14 (.A0(d2_adj_5741[12]), .B0(d1_adj_5740[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[13]), .B1(d1_adj_5740[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16246), .COUT(n16247), .S0(d2_71__N_490_adj_5757[12]), 
          .S1(d2_71__N_490_adj_5757[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_24 (.A0(d2_adj_5741[22]), .B0(d1_adj_5740[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[23]), .B1(d1_adj_5740[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16251), .COUT(n16252), .S0(d2_71__N_490_adj_5757[22]), 
          .S1(d2_71__N_490_adj_5757[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_36 (.A0(d2_adj_5741[34]), .B0(d1_adj_5740[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[35]), .B1(d1_adj_5740[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16257), .COUT(n16258), .S0(d2_71__N_490_adj_5757[34]), 
          .S1(d2_71__N_490_adj_5757[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_22 (.A0(d2_adj_5741[20]), .B0(d1_adj_5740[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[21]), .B1(d1_adj_5740[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16250), .COUT(n16251), .S0(d2_71__N_490_adj_5757[20]), 
          .S1(d2_71__N_490_adj_5757[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_34 (.A0(d2_adj_5741[32]), .B0(d1_adj_5740[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[33]), .B1(d1_adj_5740[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16256), .COUT(n16257), .S0(d2_71__N_490_adj_5757[32]), 
          .S1(d2_71__N_490_adj_5757[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_15 (.A0(count[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16301), .COUT(n16302), .S0(n42_adj_5330), 
          .S1(n39_adj_5329));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1427_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1427_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1427_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16300), .COUT(n16301), .S0(n48_adj_5332), 
          .S1(n45_adj_5331));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1427_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1427_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1427_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_13.INJECT1_1 = "NO";
    LUT4 i2364_3_lut_4_lut (.A(n18075), .B(n17937), .C(n18076), .D(n151_adj_5638), 
         .Z(n12162)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2364_3_lut_4_lut.init = 16'hfb0b;
    CCU2C _add_1_1427_add_4_17 (.A0(count[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16302), .S0(n36_adj_5328));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1427_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1427_add_4_17.INIT1 = 16'h0000;
    defparam _add_1_1427_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16299), .COUT(n16300), .S0(n54_adj_5334), 
          .S1(n51_adj_5333));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1427_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1427_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1427_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16298), .COUT(n16299), .S0(n60_adj_5336), .S1(n57_adj_5335));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1427_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1427_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1427_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16297), .COUT(n16298), .S0(n66_adj_5338), .S1(n63_adj_5337));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1427_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1427_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1427_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16296), .COUT(n16297), .S0(n72_adj_5340), .S1(n69_adj_5339));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1427_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1427_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1427_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5534), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16180));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1519_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1519_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_21 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n129_adj_5306), .D0(d1[54]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n126_adj_5305), .D1(d1[55]), .CIN(n16189), .COUT(n16190), 
          .S0(d1_71__N_418[54]), .S1(d1_71__N_418[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_16 (.A0(d_d_tmp[13]), .B0(d_tmp[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[14]), .B1(d_tmp[14]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16265), .COUT(n16266), .S0(d6_71__N_1459[13]), 
          .S1(d6_71__N_1459[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_6 (.A0(d_d_tmp[3]), .B0(d_tmp[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[4]), .B1(d_tmp[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16260), .COUT(n16261), .S0(d6_71__N_1459[3]), 
          .S1(d6_71__N_1459[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_6.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i63 (.D(phase_inc_carrGen[63]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i63.GSR = "ENABLED";
    CCU2C _add_1_1477_add_4_7 (.A0(d6_adj_5745[40]), .B0(cout_adj_4625), 
          .C0(n171_adj_4947), .D0(n33_adj_4720), .A1(d6_adj_5745[41]), 
          .B1(cout_adj_4625), .C1(n168_adj_4946), .D1(n32_adj_4721), .CIN(n16141), 
          .COUT(n16142), .S0(d7_71__N_1531_adj_5773[40]), .S1(d7_71__N_1531_adj_5773[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_5 (.A0(d6_adj_5745[38]), .B0(cout_adj_4625), 
          .C0(n177_adj_4949), .D0(n35_adj_4718), .A1(d6_adj_5745[39]), 
          .B1(cout_adj_4625), .C1(n174_adj_4948), .D1(n34_adj_4719), .CIN(n16140), 
          .COUT(n16141), .S0(d7_71__N_1531_adj_5773[38]), .S1(d7_71__N_1531_adj_5773[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_5.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i62 (.D(phase_inc_carrGen[62]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[62]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i62.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i61 (.D(phase_inc_carrGen[61]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i61.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i60 (.D(phase_inc_carrGen[60]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[60]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i60.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i59 (.D(phase_inc_carrGen[59]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i59.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i58 (.D(phase_inc_carrGen[58]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[58]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i58.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i57 (.D(phase_inc_carrGen[57]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i57.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i56 (.D(phase_inc_carrGen[56]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[56]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i56.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i55 (.D(phase_inc_carrGen[55]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i55.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i54 (.D(phase_inc_carrGen[54]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[54]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i54.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i53 (.D(phase_inc_carrGen[53]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i53.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i52 (.D(phase_inc_carrGen[52]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[52]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i52.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i51 (.D(phase_inc_carrGen[51]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i51.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i50 (.D(phase_inc_carrGen[50]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[50]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i50.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i49 (.D(phase_inc_carrGen[49]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i49.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i48 (.D(phase_inc_carrGen[48]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[48]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i48.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i47 (.D(phase_inc_carrGen[47]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i47.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i46 (.D(phase_inc_carrGen[46]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[46]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i46.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i45 (.D(phase_inc_carrGen[45]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i45.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i44 (.D(phase_inc_carrGen[44]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[44]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i44.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i43 (.D(phase_inc_carrGen[43]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i43.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i42 (.D(phase_inc_carrGen[42]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[42]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i42.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i41 (.D(phase_inc_carrGen[41]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i41.GSR = "ENABLED";
    CCU2C _add_1_1474_add_4_7 (.A0(d7_adj_5747[40]), .B0(cout_adj_5613), 
          .C0(n171_adj_4983), .D0(n33_adj_4681), .A1(d7_adj_5747[41]), 
          .B1(cout_adj_5613), .C1(n168_adj_4982), .D1(n32_adj_4682), .CIN(n16204), 
          .COUT(n16205), .S0(d8_71__N_1603_adj_5774[40]), .S1(d8_71__N_1603_adj_5774[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[36]), .B1(d2[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15878), .S1(n183_adj_5587));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1561_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_2.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i40 (.D(phase_inc_carrGen[40]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[40]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i40.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i39 (.D(phase_inc_carrGen[39]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i39.GSR = "ENABLED";
    CCU2C _add_1_1480_add_4_37 (.A0(d_tmp_adj_5738[70]), .B0(cout_adj_5605), 
          .C0(n81_adj_4881), .D0(n3_adj_2820), .A1(d_tmp_adj_5738[71]), 
          .B1(cout_adj_5605), .C1(n78_adj_4880), .D1(n2_adj_2821), .CIN(n15876), 
          .S0(d6_71__N_1459_adj_5772[70]), .S1(d6_71__N_1459_adj_5772[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_37.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i38 (.D(phase_inc_carrGen[38]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[38]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i38.GSR = "ENABLED";
    LUT4 mux_325_i32_4_lut (.A(n12122), .B(n226), .C(n17925), .D(n2572), 
         .Z(n2340)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i32_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1480_add_4_35 (.A0(d_tmp_adj_5738[68]), .B0(cout_adj_5605), 
          .C0(n87_adj_4883), .D0(n5_adj_2818), .A1(d_tmp_adj_5738[69]), 
          .B1(cout_adj_5605), .C1(n84_adj_4882), .D1(n4_adj_2819), .CIN(n15875), 
          .COUT(n15876), .S0(d6_71__N_1459_adj_5772[68]), .S1(d6_71__N_1459_adj_5772[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_35.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i37 (.D(phase_inc_carrGen[37]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i37.GSR = "ENABLED";
    CCU2C _add_1_1430_add_4_6 (.A0(d2_adj_5741[4]), .B0(d1_adj_5740[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[5]), .B1(d1_adj_5740[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16242), .COUT(n16243), .S0(d2_71__N_490_adj_5757[4]), 
          .S1(d2_71__N_490_adj_5757[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1480_add_4_33 (.A0(d_tmp_adj_5738[66]), .B0(cout_adj_5605), 
          .C0(n93_adj_4885), .D0(n7_adj_2816), .A1(d_tmp_adj_5738[67]), 
          .B1(cout_adj_5605), .C1(n90_adj_4884), .D1(n6_adj_2817), .CIN(n15874), 
          .COUT(n15875), .S0(d6_71__N_1459_adj_5772[66]), .S1(d6_71__N_1459_adj_5772[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_33.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i36 (.D(phase_inc_carrGen[36]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[36]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i36.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i35 (.D(phase_inc_carrGen[35]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i35.GSR = "ENABLED";
    CCU2C _add_1_1480_add_4_31 (.A0(d_tmp_adj_5738[64]), .B0(cout_adj_5605), 
          .C0(n99_adj_4887), .D0(n9), .A1(d_tmp_adj_5738[65]), .B1(cout_adj_5605), 
          .C1(n96_adj_4886), .D1(n8), .CIN(n15873), .COUT(n15874), .S0(d6_71__N_1459_adj_5772[64]), 
          .S1(d6_71__N_1459_adj_5772[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_31.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i34 (.D(phase_inc_carrGen[34]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[34]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i34.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i33 (.D(phase_inc_carrGen[33]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i33.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i32 (.D(phase_inc_carrGen[32]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[32]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i32.GSR = "ENABLED";
    CCU2C _add_1_1480_add_4_29 (.A0(d_tmp_adj_5738[62]), .B0(cout_adj_5605), 
          .C0(n105_adj_4889), .D0(n11), .A1(d_tmp_adj_5738[63]), .B1(cout_adj_5605), 
          .C1(n102_adj_4888), .D1(n10), .CIN(n15872), .COUT(n15873), 
          .S0(d6_71__N_1459_adj_5772[62]), .S1(d6_71__N_1459_adj_5772[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_29.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i31 (.D(phase_inc_carrGen[31]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i31.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i30 (.D(phase_inc_carrGen[30]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[30]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i30.GSR = "ENABLED";
    CCU2C _add_1_1519_add_4_19 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n135_adj_5308), .D0(d1[52]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n132_adj_5307), .D1(d1[53]), .CIN(n16188), .COUT(n16189), 
          .S0(d1_71__N_418[52]), .S1(d1_71__N_418[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1480_add_4_27 (.A0(d_tmp_adj_5738[60]), .B0(cout_adj_5605), 
          .C0(n111_adj_4891), .D0(n13), .A1(d_tmp_adj_5738[61]), .B1(cout_adj_5605), 
          .C1(n108_adj_4890), .D1(n12), .CIN(n15871), .COUT(n15872), 
          .S0(d6_71__N_1459_adj_5772[60]), .S1(d6_71__N_1459_adj_5772[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_27.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i29 (.D(phase_inc_carrGen[29]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i29.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i28 (.D(phase_inc_carrGen[28]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[28]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i28.GSR = "ENABLED";
    CCU2C _add_1_1480_add_4_25 (.A0(d_tmp_adj_5738[58]), .B0(cout_adj_5605), 
          .C0(n117_adj_4893), .D0(n15), .A1(d_tmp_adj_5738[59]), .B1(cout_adj_5605), 
          .C1(n114_adj_4892), .D1(n14), .CIN(n15870), .COUT(n15871), 
          .S0(d6_71__N_1459_adj_5772[58]), .S1(d6_71__N_1459_adj_5772[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_25.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i27 (.D(phase_inc_carrGen[27]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i27.GSR = "ENABLED";
    CCU2C _add_1_1480_add_4_23 (.A0(d_tmp_adj_5738[56]), .B0(cout_adj_5605), 
          .C0(n123_adj_4895), .D0(n17), .A1(d_tmp_adj_5738[57]), .B1(cout_adj_5605), 
          .C1(n120_adj_4894), .D1(n16), .CIN(n15869), .COUT(n15870), 
          .S0(d6_71__N_1459_adj_5772[56]), .S1(d6_71__N_1459_adj_5772[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1480_add_4_21 (.A0(d_tmp_adj_5738[54]), .B0(cout_adj_5605), 
          .C0(n129_adj_4897), .D0(n19), .A1(d_tmp_adj_5738[55]), .B1(cout_adj_5605), 
          .C1(n126_adj_4896), .D1(n18), .CIN(n15868), .COUT(n15869), 
          .S0(d6_71__N_1459_adj_5772[54]), .S1(d6_71__N_1459_adj_5772[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_21.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i26 (.D(phase_inc_carrGen[26]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[26]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i26.GSR = "ENABLED";
    CCU2C _add_1_1480_add_4_19 (.A0(d_tmp_adj_5738[52]), .B0(cout_adj_5605), 
          .C0(n135_adj_4899), .D0(n21), .A1(d_tmp_adj_5738[53]), .B1(cout_adj_5605), 
          .C1(n132_adj_4898), .D1(n20), .CIN(n15867), .COUT(n15868), 
          .S0(d6_71__N_1459_adj_5772[52]), .S1(d6_71__N_1459_adj_5772[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_14 (.A0(d5_adj_5744[12]), .B0(d4_adj_5743[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[13]), .B1(d4_adj_5743[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16105), .COUT(n16106), .S0(d5_71__N_706_adj_5760[12]), 
          .S1(d5_71__N_706_adj_5760[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_14.INJECT1_1 = "NO";
    LUT4 mux_750_i2_3_lut (.A(led_c_2), .B(led_c_4), .C(n2824), .Z(n3692)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_750_i2_3_lut.init = 16'hc5c5;
    CCU2C _add_1_1439_add_4_12 (.A0(d5_adj_5744[10]), .B0(d4_adj_5743[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[11]), .B1(d4_adj_5743[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16104), .COUT(n16105), .S0(d5_71__N_706_adj_5760[10]), 
          .S1(d5_71__N_706_adj_5760[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_12.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i25 (.D(phase_inc_carrGen[25]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i25.GSR = "ENABLED";
    LUT4 mux_325_i29_4_lut (.A(n12116), .B(n235), .C(n17925), .D(n2572), 
         .Z(n2343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i29_4_lut.init = 16'hcfca;
    LUT4 mux_325_i10_4_lut (.A(n12084), .B(n292), .C(n17925), .D(n2572), 
         .Z(n2362)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i10_4_lut.init = 16'hcfca;
    CCU2C _add_1_1636_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7_adj_5748[36]), .B1(d7_adj_5747[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16118), .S1(n183_adj_4987));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1636_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1430_add_4_10 (.A0(d2_adj_5741[8]), .B0(d1_adj_5740[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[9]), .B1(d1_adj_5740[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16244), .COUT(n16245), .S0(d2_71__N_490_adj_5757[8]), 
          .S1(d2_71__N_490_adj_5757[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1430_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1430_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1430_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1430_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_17 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n141_adj_5310), .D0(d1[50]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n138_adj_5309), .D1(d1[51]), .CIN(n16187), .COUT(n16188), 
          .S0(d1_71__N_418[50]), .S1(d1_71__N_418[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_5 (.A0(d7_adj_5747[38]), .B0(cout_adj_5613), 
          .C0(n177_adj_4985), .D0(n35_adj_4679), .A1(d7_adj_5747[39]), 
          .B1(cout_adj_5613), .C1(n174_adj_4984), .D1(n34_adj_4680), .CIN(n16203), 
          .COUT(n16204), .S0(d8_71__N_1603_adj_5774[38]), .S1(d8_71__N_1603_adj_5774[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_5.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i24 (.D(phase_inc_carrGen[24]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[24]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i24.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i23 (.D(phase_inc_carrGen[23]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i23.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i22 (.D(phase_inc_carrGen[22]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[22]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i22.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i21 (.D(phase_inc_carrGen[21]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i21.GSR = "ENABLED";
    LUT4 i45_4_lut_4_lut_4_lut (.A(led_c_3), .B(led_c_0), .C(led_c_1), 
         .D(led_c_2), .Z(n29_adj_5730)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i45_4_lut_4_lut_4_lut.init = 16'h6014;
    LUT4 led_c_3_bdd_4_lut_6449 (.A(led_c_3), .B(n313), .C(n17069), .D(led_c_4), 
         .Z(n17955)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !(C)))) */ ;
    defparam led_c_3_bdd_4_lut_6449.init = 16'h4505;
    LUT4 PWMOut_I_0_1_lut (.A(PWMOutP4_c), .Z(PWMOutN4_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(92[22:29])
    defparam PWMOut_I_0_1_lut.init = 16'h5555;
    CCU2C _add_1_1480_add_4_17 (.A0(d_tmp_adj_5738[50]), .B0(cout_adj_5605), 
          .C0(n141_adj_4901), .D0(n23), .A1(d_tmp_adj_5738[51]), .B1(cout_adj_5605), 
          .C1(n138_adj_4900), .D1(n22), .CIN(n15866), .COUT(n15867), 
          .S0(d6_71__N_1459_adj_5772[50]), .S1(d6_71__N_1459_adj_5772[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_17.INJECT1_1 = "NO";
    LUT4 CIC_out_clkSin_c_bdd_2_lut_6409_rep_154_3_lut_4_lut (.A(led_c_4), 
         .B(n17940), .C(n12563), .D(n17900), .Z(n17926)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;
    defparam CIC_out_clkSin_c_bdd_2_lut_6409_rep_154_3_lut_4_lut.init = 16'hf0b0;
    SinCos SinCos_inst (.clk_80mhz(clk_80mhz), .VCC_net(VCC_net), .GND_net(GND_net), 
           .\phase_accum[57] (phase_accum[57]), .\phase_accum[58] (phase_accum[58]), 
           .\phase_accum[59] (phase_accum[59]), .\phase_accum[60] (phase_accum[60]), 
           .\phase_accum[61] (phase_accum[61]), .\phase_accum[62] (phase_accum[62]), 
           .\phase_accum[63] (phase_accum[63]), .\LOSine[1] (LOSine[1]), 
           .\LOSine[2] (LOSine[2]), .\LOSine[3] (LOSine[3]), .\LOSine[4] (LOSine[4]), 
           .\LOSine[5] (LOSine[5]), .\LOSine[6] (LOSine[6]), .\LOSine[7] (LOSine[7]), 
           .\LOSine[8] (LOSine[8]), .\LOSine[9] (LOSine[9]), .\LOSine[10] (LOSine[10]), 
           .\LOSine[11] (LOSine[11]), .\LOSine[12] (LOSine[12]), .\LOCosine[1] (LOCosine[1]), 
           .\LOCosine[2] (LOCosine[2]), .\LOCosine[3] (LOCosine[3]), .\LOCosine[4] (LOCosine[4]), 
           .\LOCosine[5] (LOCosine[5]), .\LOCosine[6] (LOCosine[6]), .\LOCosine[7] (LOCosine[7]), 
           .\LOCosine[8] (LOCosine[8]), .\LOCosine[9] (LOCosine[9]), .\LOCosine[10] (LOCosine[10]), 
           .\LOCosine[11] (LOCosine[11]), .\LOCosine[12] (LOCosine[12]), 
           .\phase_accum[56] (phase_accum[56])) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    LUT4 mux_325_i4_4_lut_4_lut_4_lut_then_3_lut (.A(led_c_3), .B(n310), 
         .C(led_c_4), .Z(n17960)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam mux_325_i4_4_lut_4_lut_4_lut_then_3_lut.init = 16'h4545;
    LUT4 mux_325_i4_4_lut_4_lut_4_lut_else_3_lut (.A(led_c_3), .B(n17937), 
         .C(led_c_2), .Z(n17959)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam mux_325_i4_4_lut_4_lut_4_lut_else_3_lut.init = 16'h4040;
    FD1S3AX phase_inc_carrGen1_i20 (.D(phase_inc_carrGen[20]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[20]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i20.GSR = "ENABLED";
    CCU2C _add_1_1477_add_4_3 (.A0(d6_adj_5745[36]), .B0(cout_adj_4625), 
          .C0(n183_adj_4951), .D0(n37_adj_4715), .A1(d6_adj_5745[37]), 
          .B1(cout_adj_4625), .C1(n180_adj_4950), .D1(n36_adj_4716), .CIN(n16139), 
          .COUT(n16140), .S0(d7_71__N_1531_adj_5773[36]), .S1(d7_71__N_1531_adj_5773[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1477_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1477_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_3.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i19 (.D(phase_inc_carrGen[19]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i19.GSR = "ENABLED";
    CCU2C _add_1_1531_add_4_10 (.A0(d_d_tmp[7]), .B0(d_tmp[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[8]), .B1(d_tmp[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16262), .COUT(n16263), .S0(d6_71__N_1459[7]), 
          .S1(d6_71__N_1459[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_10.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i18 (.D(phase_inc_carrGen[18]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[18]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i18.GSR = "ENABLED";
    CCU2C _add_1_1531_add_4_24 (.A0(d_d_tmp[21]), .B0(d_tmp[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[22]), .B1(d_tmp[22]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16269), .COUT(n16270), .S0(d6_71__N_1459[21]), 
          .S1(d6_71__N_1459[22]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_24.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut (.A(led_c_4), .B(n17948), .C(led_c_6), .D(n17097), 
         .Z(n12563)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff7f;
    CCU2C _add_1_1531_add_4_18 (.A0(d_d_tmp[15]), .B0(d_tmp[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[16]), .B1(d_tmp[16]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16266), .COUT(n16267), .S0(d6_71__N_1459[15]), 
          .S1(d6_71__N_1459[16]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_28 (.A0(d_d_tmp[25]), .B0(d_tmp[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[26]), .B1(d_tmp[26]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16271), .COUT(n16272), .S0(d6_71__N_1459[25]), 
          .S1(d6_71__N_1459[26]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_12 (.A0(d_d_tmp[9]), .B0(d_tmp[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[10]), .B1(d_tmp[10]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16263), .COUT(n16264), .S0(d6_71__N_1459[9]), 
          .S1(d6_71__N_1459[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1531_add_4_26 (.A0(d_d_tmp[23]), .B0(d_tmp[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[24]), .B1(d_tmp[24]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16270), .COUT(n16271), .S0(d6_71__N_1459[23]), 
          .S1(d6_71__N_1459[24]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_26.INJECT1_1 = "NO";
    LUT4 i6357_3_lut_4_lut (.A(led_c_6), .B(n17948), .C(led_c_4), .D(n29_adj_5730), 
         .Z(n17205)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i6357_3_lut_4_lut.init = 16'hf7ff;
    CCU2C _add_1_1531_add_4_14 (.A0(d_d_tmp[11]), .B0(d_tmp[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[12]), .B1(d_tmp[12]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16264), .COUT(n16265), .S0(d6_71__N_1459[11]), 
          .S1(d6_71__N_1459[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1531_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1531_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1531_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1531_add_4_14.INJECT1_1 = "NO";
    LUT4 n17900_bdd_2_lut_rep_162_3_lut_4_lut (.A(led_c_6), .B(n17948), 
         .C(n17900), .D(led_c_4), .Z(n17934)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam n17900_bdd_2_lut_rep_162_3_lut_4_lut.init = 16'hfff7;
    FD1S3AX phase_inc_carrGen1_i17 (.D(phase_inc_carrGen[17]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i17.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i16 (.D(phase_inc_carrGen[16]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[16]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i16.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i15 (.D(phase_inc_carrGen[15]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i15.GSR = "ENABLED";
    CCU2C _add_1_1424_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16321), .S0(cout_adj_5327));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1424_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1424_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_36 (.A0(d1_adj_5740[34]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[35]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16320), .COUT(n16321), .S0(d1_71__N_418_adj_5756[34]), 
          .S1(d1_71__N_418_adj_5756[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1480_add_4_15 (.A0(d_tmp_adj_5738[48]), .B0(cout_adj_5605), 
          .C0(n147_adj_4903), .D0(n25_adj_2814), .A1(d_tmp_adj_5738[49]), 
          .B1(cout_adj_5605), .C1(n144_adj_4902), .D1(n24_adj_2815), .CIN(n15865), 
          .COUT(n15866), .S0(d6_71__N_1459_adj_5772[48]), .S1(d6_71__N_1459_adj_5772[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_34 (.A0(d1_adj_5740[32]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[33]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16319), .COUT(n16320), .S0(d1_71__N_418_adj_5756[32]), 
          .S1(d1_71__N_418_adj_5756[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_10 (.A0(d5_adj_5744[8]), .B0(d4_adj_5743[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[9]), .B1(d4_adj_5743[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16103), .COUT(n16104), .S0(d5_71__N_706_adj_5760[8]), 
          .S1(d5_71__N_706_adj_5760[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16295), .COUT(n16296), .S0(n78_adj_5342), .S1(n75_adj_5341));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1427_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1427_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1427_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1477_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_4625), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16139));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1477_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1477_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1477_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1477_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_38 (.A0(d_d7_adj_5748[71]), .B0(d7_adj_5747[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16135), .S0(n78_adj_4952));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1636_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_38.INJECT1_1 = "NO";
    LUT4 i3143_2_lut_rep_157 (.A(led_c_4), .B(n2824), .Z(n17929)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i3143_2_lut_rep_157.init = 16'h8888;
    CCU2C _add_1_1439_add_4_8 (.A0(d5_adj_5744[6]), .B0(d4_adj_5743[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[7]), .B1(d4_adj_5743[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16102), .COUT(n16103), .S0(d5_71__N_706_adj_5760[6]), 
          .S1(d5_71__N_706_adj_5760[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_36 (.A0(d_d7_adj_5748[69]), .B0(d7_adj_5747[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[70]), .B1(d7_adj_5747[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16134), .COUT(n16135), .S0(n84_adj_4954), 
          .S1(n81_adj_4953));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_34 (.A0(d_d7_adj_5748[67]), .B0(d7_adj_5747[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[68]), .B1(d7_adj_5747[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16133), .COUT(n16134), .S0(n90_adj_4956), 
          .S1(n87_adj_4955));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_32 (.A0(d_d7_adj_5748[65]), .B0(d7_adj_5747[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[66]), .B1(d7_adj_5747[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16132), .COUT(n16133), .S0(n96_adj_4958), 
          .S1(n93_adj_4957));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_30 (.A0(d_d7_adj_5748[63]), .B0(d7_adj_5747[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[64]), .B1(d7_adj_5747[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16131), .COUT(n16132), .S0(n102_adj_4960), 
          .S1(n99_adj_4959));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_38 (.A0(d_d9[35]), .B0(d9[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16294), .S1(cout_adj_4756));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1627_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1480_add_4_13 (.A0(d_tmp_adj_5738[46]), .B0(cout_adj_5605), 
          .C0(n153_adj_4905), .D0(n27_adj_2812), .A1(d_tmp_adj_5738[47]), 
          .B1(cout_adj_5605), .C1(n150_adj_4904), .D1(n26_adj_2813), .CIN(n15864), 
          .COUT(n15865), .S0(d6_71__N_1459_adj_5772[46]), .S1(d6_71__N_1459_adj_5772[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_13.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i14 (.D(phase_inc_carrGen[14]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i14.GSR = "ENABLED";
    CCU2C _add_1_1636_add_4_28 (.A0(d_d7_adj_5748[61]), .B0(d7_adj_5747[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[62]), .B1(d7_adj_5747[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16130), .COUT(n16131), .S0(n108_adj_4962), 
          .S1(n105_adj_4961));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_26 (.A0(d_d7_adj_5748[59]), .B0(d7_adj_5747[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[60]), .B1(d7_adj_5747[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16129), .COUT(n16130), .S0(n114_adj_4964), 
          .S1(n111_adj_4963));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_24 (.A0(d_d7_adj_5748[57]), .B0(d7_adj_5747[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[58]), .B1(d7_adj_5747[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16128), .COUT(n16129), .S0(n120_adj_4966), 
          .S1(n117_adj_4965));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_22 (.A0(d_d7_adj_5748[55]), .B0(d7_adj_5747[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[56]), .B1(d7_adj_5747[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16127), .COUT(n16128), .S0(n126_adj_4968), 
          .S1(n123_adj_4967));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_20 (.A0(d_d7_adj_5748[53]), .B0(d7_adj_5747[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[54]), .B1(d7_adj_5747[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16126), .COUT(n16127), .S0(n132_adj_4970), 
          .S1(n129_adj_4969));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_18 (.A0(d_d7_adj_5748[51]), .B0(d7_adj_5747[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[52]), .B1(d7_adj_5747[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16125), .COUT(n16126), .S0(n138_adj_4972), 
          .S1(n135_adj_4971));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_16 (.A0(d_d7_adj_5748[49]), .B0(d7_adj_5747[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[50]), .B1(d7_adj_5747[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16124), .COUT(n16125), .S0(n144_adj_4974), 
          .S1(n141_adj_4973));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_16.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i13 (.D(phase_inc_carrGen[13]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i13.GSR = "ENABLED";
    CCU2C _add_1_1636_add_4_14 (.A0(d_d7_adj_5748[47]), .B0(d7_adj_5747[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[48]), .B1(d7_adj_5747[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16123), .COUT(n16124), .S0(n150_adj_4976), 
          .S1(n147_adj_4975));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_14.INJECT1_1 = "NO";
    FD1S3AX _add_1_1654_i7 (.D(cout_adj_5112), .CK(clk_80mhz), .Q(PWMOutP4_c));
    defparam _add_1_1654_i7.GSR = "ENABLED";
    OB led_pad_6 (.I(led_c_6), .O(led[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    CCU2C _add_1_1439_add_4_6 (.A0(d5_adj_5744[4]), .B0(d4_adj_5743[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[5]), .B1(d4_adj_5743[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16101), .COUT(n16102), .S0(d5_71__N_706_adj_5760[4]), 
          .S1(d5_71__N_706_adj_5760[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_4 (.A0(d5_adj_5744[2]), .B0(d4_adj_5743[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[3]), .B1(d4_adj_5743[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16100), .COUT(n16101), .S0(d5_71__N_706_adj_5760[2]), 
          .S1(d5_71__N_706_adj_5760[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_2 (.A0(d5_adj_5744[0]), .B0(d4_adj_5743[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[1]), .B1(d4_adj_5743[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16100), .S1(d5_71__N_706_adj_5760[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1439_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_38 (.A0(d5[71]), .B0(d4[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16098), .S0(n78_adj_5364));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1567_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_36 (.A0(d5[69]), .B0(d4[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[70]), .B1(d4[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16097), .COUT(n16098), .S0(n84_adj_5366), .S1(n81_adj_5365));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_34 (.A0(d5[67]), .B0(d4[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[68]), .B1(d4[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16096), .COUT(n16097), .S0(n90_adj_5368), .S1(n87_adj_5367));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_32 (.A0(d5[65]), .B0(d4[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[66]), .B1(d4[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16095), .COUT(n16096), .S0(n96_adj_5370), .S1(n93_adj_5369));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_30 (.A0(d5[63]), .B0(d4[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[64]), .B1(d4[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16094), .COUT(n16095), .S0(n102_adj_5372), .S1(n99_adj_5371));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_28 (.A0(d5[61]), .B0(d4[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[62]), .B1(d4[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16093), .COUT(n16094), .S0(n108_adj_5374), .S1(n105_adj_5373));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_26 (.A0(d5[59]), .B0(d4[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[60]), .B1(d4[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16092), .COUT(n16093), .S0(n114_adj_5376), .S1(n111_adj_5375));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1480_add_4_11 (.A0(d_tmp_adj_5738[44]), .B0(cout_adj_5605), 
          .C0(n159_adj_4907), .D0(n29_adj_2810), .A1(d_tmp_adj_5738[45]), 
          .B1(cout_adj_5605), .C1(n156_adj_4906), .D1(n28_adj_2811), .CIN(n15863), 
          .COUT(n15864), .S0(d6_71__N_1459_adj_5772[44]), .S1(d6_71__N_1459_adj_5772[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_24 (.A0(d5[57]), .B0(d4[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[58]), .B1(d4[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16091), .COUT(n16092), .S0(n120_adj_5378), .S1(n117_adj_5377));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_24.INJECT1_1 = "NO";
    LUT4 i3242_1_lut_2_lut (.A(led_c_4), .B(n2824), .Z(n3677)) /* synthesis lut_function=(!(A (B))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i3242_1_lut_2_lut.init = 16'h7777;
    LUT4 i2352_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(led_c_3), .D(n172_adj_5645), 
         .Z(n12150)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2352_3_lut_4_lut.init = 16'hfb0b;
    CCU2C _add_1_1627_add_4_30 (.A0(d_d9[27]), .B0(d9[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[28]), .B1(d9[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16290), .COUT(n16291));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_22 (.A0(d5[55]), .B0(d4[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[56]), .B1(d4[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16090), .COUT(n16091), .S0(n126_adj_5380), .S1(n123_adj_5379));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_20 (.A0(d5[53]), .B0(d4[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[54]), .B1(d4[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16089), .COUT(n16090), .S0(n132_adj_5382), .S1(n129_adj_5381));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_20.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i12 (.D(phase_inc_carrGen[12]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i12.GSR = "ENABLED";
    CCU2C _add_1_1567_add_4_18 (.A0(d5[51]), .B0(d4[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[52]), .B1(d4[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16088), .COUT(n16089), .S0(n138_adj_5384), .S1(n135_adj_5383));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1427_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16295), .S1(n81_adj_5343));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1427_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1427_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1427_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1427_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_32 (.A0(d1_adj_5740[30]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[31]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16318), .COUT(n16319), .S0(d1_71__N_418_adj_5756[30]), 
          .S1(d1_71__N_418_adj_5756[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_16 (.A0(d5[49]), .B0(d4[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[50]), .B1(d4[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16087), .COUT(n16088), .S0(n144_adj_5386), .S1(n141_adj_5385));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_14 (.A0(d5[47]), .B0(d4[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[48]), .B1(d4[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16086), .COUT(n16087), .S0(n150_adj_5388), .S1(n147_adj_5387));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_12 (.A0(d_d7_adj_5748[45]), .B0(d7_adj_5747[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[46]), .B1(d7_adj_5747[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16122), .COUT(n16123), .S0(n156_adj_4978), 
          .S1(n153_adj_4977));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_12 (.A0(d5[45]), .B0(d4[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[46]), .B1(d4[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16085), .COUT(n16086), .S0(n156_adj_5390), .S1(n153_adj_5389));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1424_add_4_30 (.A0(d1_adj_5740[28]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[29]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16317), .COUT(n16318), .S0(d1_71__N_418_adj_5756[28]), 
          .S1(d1_71__N_418_adj_5756[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1424_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1424_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1424_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1424_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_3 (.A0(d7_adj_5747[36]), .B0(cout_adj_5613), 
          .C0(n183_adj_4987), .D0(n37_adj_4677), .A1(d7_adj_5747[37]), 
          .B1(cout_adj_5613), .C1(n180_adj_4986), .D1(n36_adj_4678), .CIN(n16202), 
          .COUT(n16203), .S0(d8_71__N_1603_adj_5774[36]), .S1(d8_71__N_1603_adj_5774[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_10 (.A0(d5[43]), .B0(d4[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[44]), .B1(d4[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16084), .COUT(n16085), .S0(n162_adj_5392), .S1(n159_adj_5391));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_8 (.A0(d5[41]), .B0(d4[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[42]), .B1(d4[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16083), .COUT(n16084), .S0(n168_adj_5394), .S1(n165_adj_5393));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_8.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i11 (.D(phase_inc_carrGen[11]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i11.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i10 (.D(phase_inc_carrGen[10]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i10.GSR = "ENABLED";
    CCU2C _add_1_1567_add_4_6 (.A0(d5[39]), .B0(d4[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[40]), .B1(d4[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16082), .COUT(n16083), .S0(n174_adj_5396), .S1(n171_adj_5395));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_6.INJECT1_1 = "NO";
    LUT4 i5289_2_lut_rep_170 (.A(ISquare[23]), .B(ISquare[22]), .Z(n17942)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam i5289_2_lut_rep_170.init = 16'heeee;
    LUT4 led_c_4_bdd_4_lut (.A(n18075), .B(led_c_0), .C(n18076), .D(led_c_1), 
         .Z(n17905)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !(B+(C (D)+!C !(D)))) */ ;
    defparam led_c_4_bdd_4_lut.init = 16'hab90;
    LUT4 i5418_4_lut (.A(n17401), .B(n17940), .C(n17906), .D(n17777), 
         .Z(clk_80mhz_enable_1469)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C))) */ ;
    defparam i5418_4_lut.init = 16'hc0c8;
    LUT4 mux_750_i3_3_lut_rep_158 (.A(led_c_2), .B(led_c_4), .C(n2824), 
         .Z(n17930)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_750_i3_3_lut_rep_158.init = 16'hcaca;
    LUT4 i2011_1_lut_3_lut (.A(led_c_2), .B(led_c_4), .C(n2824), .Z(n11804)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2011_1_lut_3_lut.init = 16'h3535;
    LUT4 n17905_bdd_2_lut (.A(n17905), .B(led_c_4), .Z(n17906)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n17905_bdd_2_lut.init = 16'h2222;
    FD1S3AX phase_inc_carrGen1_i9 (.D(phase_inc_carrGen[9]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i9.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i8 (.D(phase_inc_carrGen[8]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i8.GSR = "ENABLED";
    LUT4 i3146_rep_114_2_lut (.A(led_c_2), .B(led_c_1), .Z(n17777)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3146_rep_114_2_lut.init = 16'heeee;
    CCU2C _add_1_1567_add_4_4 (.A0(d5[37]), .B0(d4[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[38]), .B1(d4[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16081), .COUT(n16082), .S0(n180_adj_5398), .S1(n177_adj_5397));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1567_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1567_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[36]), .B1(d4[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16081), .S1(n183_adj_5399));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1567_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1567_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1567_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1567_add_4_2.INJECT1_1 = "NO";
    FD1S3AX phase_inc_carrGen1_i7 (.D(phase_inc_carrGen[7]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i7.GSR = "ENABLED";
    LUT4 i5333_1_lut_2_lut_3_lut (.A(ISquare[23]), .B(ISquare[22]), .C(ISquare[31]), 
         .Z(n23_adj_2823)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam i5333_1_lut_2_lut_3_lut.init = 16'h0101;
    OB led_pad_7 (.I(led_c_7), .O(led[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    OB o_Tx_Serial_pad (.I(GND_net), .O(o_Tx_Serial));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(43[22:33])
    FD1S3AX phase_inc_carrGen1_i6 (.D(phase_inc_carrGen[6]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i6.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i5 (.D(phase_inc_carrGen[5]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i5.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i4 (.D(phase_inc_carrGen[4]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i4.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i3 (.D(phase_inc_carrGen[3]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i3.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i2 (.D(phase_inc_carrGen[2]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i2.GSR = "ENABLED";
    FD1S3AX phase_inc_carrGen1_i1 (.D(phase_inc_carrGen[1]), .CK(clk_80mhz), 
            .Q(phase_inc_carrGen1[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen1_i1.GSR = "ENABLED";
    CCU2C _add_1_1615_add_4_38 (.A0(d_d6_adj_5746[35]), .B0(d6_adj_5745[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16080), .S0(d7_71__N_1531_adj_5773[35]), 
          .S1(cout_adj_4625));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1615_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_38.INJECT1_1 = "NO";
    OB led_pad_5 (.I(led_c_5), .O(led[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    FD1S3AX o_Rx_Byte_i8 (.D(o_Rx_Byte1[7]), .CK(clk_80mhz), .Q(led_c_7));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam o_Rx_Byte_i8.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i7 (.D(o_Rx_Byte1[6]), .CK(clk_80mhz), .Q(led_c_6));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i6 (.D(o_Rx_Byte1[5]), .CK(clk_80mhz), .Q(led_c_5));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i5 (.D(o_Rx_Byte1[4]), .CK(clk_80mhz), .Q(led_c_4));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i4 (.D(o_Rx_Byte1[3]), .CK(clk_80mhz), .Q(led_c_3));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i3 (.D(o_Rx_Byte1[2]), .CK(clk_80mhz), .Q(led_c_2));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1S3AX o_Rx_Byte_i2 (.D(o_Rx_Byte1[1]), .CK(clk_80mhz), .Q(led_c_1));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    CCU2C _add_1_1406_add_4_32 (.A0(d1[30]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[31]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16337), .COUT(n16338), .S0(d1_71__N_418[30]), 
          .S1(d1_71__N_418[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5613), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16202));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1474_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1474_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1627_add_4_26 (.A0(d_d9[23]), .B0(d9[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[24]), .B1(d9[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16288), .COUT(n16289));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_36 (.A0(d_d6_adj_5746[33]), .B0(d6_adj_5745[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[34]), .B1(d6_adj_5745[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16079), .COUT(n16080), .S0(d7_71__N_1531_adj_5773[33]), 
          .S1(d7_71__N_1531_adj_5773[34]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_36.INJECT1_1 = "NO";
    LUT4 mux_325_i30_4_lut (.A(n2542), .B(n232), .C(n17925), .D(n2572), 
         .Z(n2342)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i30_4_lut.init = 16'hc0ca;
    LUT4 i1_2_lut_rep_166_3_lut (.A(ISquare[23]), .B(ISquare[22]), .C(ISquare[31]), 
         .Z(n17938)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam i1_2_lut_rep_166_3_lut.init = 16'hfefe;
    OB led_pad_4 (.I(led_c_4), .O(led[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    OB led_pad_3 (.I(led_c_3), .O(led[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    OB led_pad_2 (.I(led_c_2), .O(led[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    OB led_pad_1 (.I(led_c_1), .O(led[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    OB led_pad_0 (.I(led_c_0), .O(led[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    OB XOut_pad (.I(GND_net), .O(XOut));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(45[22:26])
    OB DiffOut_pad (.I(DiffOut_c), .O(DiffOut));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(46[22:29])
    OB PWMOut_pad (.I(PWMOutP4_c), .O(PWMOut));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(47[22:28])
    OB PWMOutP1_pad (.I(PWMOutP4_c), .O(PWMOutP1));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(48[22:30])
    OB PWMOutP2_pad (.I(PWMOutP4_c), .O(PWMOutP2));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(49[22:30])
    OB PWMOutP3_pad (.I(PWMOutP4_c), .O(PWMOutP3));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(50[22:30])
    OB PWMOutP4_pad (.I(PWMOutP4_c), .O(PWMOutP4));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(51[22:30])
    OB PWMOutN1_pad (.I(PWMOutN4_c), .O(PWMOutN1));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(52[22:30])
    OB PWMOutN2_pad (.I(PWMOutN4_c), .O(PWMOutN2));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(53[22:30])
    OB PWMOutN3_pad (.I(PWMOutN4_c), .O(PWMOutN3));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(54[22:30])
    OB PWMOutN4_pad (.I(PWMOutN4_c), .O(PWMOutN4));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(55[22:30])
    OB sinGen_pad (.I(sinGen_c), .O(sinGen));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(56[22:28])
    OB sin_out_pad (.I(GND_net), .O(sin_out));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(57[22:29])
    OB CIC_out_clkSin_pad (.I(GND_net), .O(CIC_out_clkSin));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(58[22:36])
    IB clk_25mhz_pad (.I(clk_25mhz), .O(clk_25mhz_c));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(40[22:31])
    IB i_Rx_Serial_pad (.I(i_Rx_Serial), .O(i_Rx_Serial_c));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(41[22:33])
    IB RFIn_pad (.I(RFIn), .O(RFIn_c));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(42[22:26])
    CCU2C _add_1_1433_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16239), .S0(cout_adj_5345));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1433_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1433_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_36 (.A0(d3_adj_5742[34]), .B0(d2_adj_5741[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[35]), .B1(d2_adj_5741[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16238), .COUT(n16239), .S0(d3_71__N_562_adj_5758[34]), 
          .S1(d3_71__N_562_adj_5758[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_34 (.A0(d3_adj_5742[32]), .B0(d2_adj_5741[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[33]), .B1(d2_adj_5741[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16237), .COUT(n16238), .S0(d3_71__N_562_adj_5758[32]), 
          .S1(d3_71__N_562_adj_5758[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_34.INJECT1_1 = "NO";
    LUT4 i5317_2_lut_3_lut (.A(ISquare[23]), .B(ISquare[22]), .C(ISquare[31]), 
         .Z(n15173)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam i5317_2_lut_3_lut.init = 16'h0e0e;
    CCU2C _add_1_1433_add_4_32 (.A0(d3_adj_5742[30]), .B0(d2_adj_5741[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[31]), .B1(d2_adj_5741[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16236), .COUT(n16237), .S0(d3_71__N_562_adj_5758[30]), 
          .S1(d3_71__N_562_adj_5758[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_30 (.A0(d3_adj_5742[28]), .B0(d2_adj_5741[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[29]), .B1(d2_adj_5741[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16235), .COUT(n16236), .S0(d3_71__N_562_adj_5758[28]), 
          .S1(d3_71__N_562_adj_5758[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_30.INJECT1_1 = "NO";
    LUT4 n17317_bdd_4_lut (.A(n17317), .B(n17090), .C(n18075), .D(n17940), 
         .Z(n2824)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n17317_bdd_4_lut.init = 16'hca00;
    CCU2C _add_1_1433_add_4_28 (.A0(d3_adj_5742[26]), .B0(d2_adj_5741[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[27]), .B1(d2_adj_5741[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16234), .COUT(n16235), .S0(d3_71__N_562_adj_5758[26]), 
          .S1(d3_71__N_562_adj_5758[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_26 (.A0(d3_adj_5742[24]), .B0(d2_adj_5741[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[25]), .B1(d2_adj_5741[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16233), .COUT(n16234), .S0(d3_71__N_562_adj_5758[24]), 
          .S1(d3_71__N_562_adj_5758[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_26.INJECT1_1 = "NO";
    LUT4 i2322_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(led_c_3), .D(n223_adj_5662), 
         .Z(n12120)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2322_3_lut_4_lut.init = 16'hf808;
    CCU2C _add_1_1433_add_4_24 (.A0(d3_adj_5742[22]), .B0(d2_adj_5741[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[23]), .B1(d2_adj_5741[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16232), .COUT(n16233), .S0(d3_71__N_562_adj_5758[22]), 
          .S1(d3_71__N_562_adj_5758[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_24.INJECT1_1 = "NO";
    LUT4 i5307_1_lut_2_lut (.A(ISquare[23]), .B(ISquare[22]), .Z(n32_adj_2822)) /* synthesis lut_function=(!(A+(B))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam i5307_1_lut_2_lut.init = 16'h1111;
    CCU2C _add_1_1433_add_4_22 (.A0(d3_adj_5742[20]), .B0(d2_adj_5741[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[21]), .B1(d2_adj_5741[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16231), .COUT(n16232), .S0(d3_71__N_562_adj_5758[20]), 
          .S1(d3_71__N_562_adj_5758[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_20 (.A0(d3_adj_5742[18]), .B0(d2_adj_5741[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[19]), .B1(d2_adj_5741[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16230), .COUT(n16231), .S0(d3_71__N_562_adj_5758[18]), 
          .S1(d3_71__N_562_adj_5758[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_18 (.A0(d3_adj_5742[16]), .B0(d2_adj_5741[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[17]), .B1(d2_adj_5741[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16229), .COUT(n16230), .S0(d3_71__N_562_adj_5758[16]), 
          .S1(d3_71__N_562_adj_5758[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_16 (.A0(d3_adj_5742[14]), .B0(d2_adj_5741[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[15]), .B1(d2_adj_5741[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16228), .COUT(n16229), .S0(d3_71__N_562_adj_5758[14]), 
          .S1(d3_71__N_562_adj_5758[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_14 (.A0(d3_adj_5742[12]), .B0(d2_adj_5741[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[13]), .B1(d2_adj_5741[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16227), .COUT(n16228), .S0(d3_71__N_562_adj_5758[12]), 
          .S1(d3_71__N_562_adj_5758[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_12 (.A0(d3_adj_5742[10]), .B0(d2_adj_5741[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[11]), .B1(d2_adj_5741[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16226), .COUT(n16227), .S0(d3_71__N_562_adj_5758[10]), 
          .S1(d3_71__N_562_adj_5758[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_10 (.A0(d3_adj_5742[8]), .B0(d2_adj_5741[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[9]), .B1(d2_adj_5741[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16225), .COUT(n16226), .S0(d3_71__N_562_adj_5758[8]), 
          .S1(d3_71__N_562_adj_5758[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_8 (.A0(d3_adj_5742[6]), .B0(d2_adj_5741[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[7]), .B1(d2_adj_5741[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16224), .COUT(n16225), .S0(d3_71__N_562_adj_5758[6]), 
          .S1(d3_71__N_562_adj_5758[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_6 (.A0(d3_adj_5742[4]), .B0(d2_adj_5741[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[5]), .B1(d2_adj_5741[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16223), .COUT(n16224), .S0(d3_71__N_562_adj_5758[4]), 
          .S1(d3_71__N_562_adj_5758[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_6.INJECT1_1 = "NO";
    LUT4 i2346_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(n18076), .D(n184_adj_5649), 
         .Z(n12144)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2346_3_lut_4_lut.init = 16'hfb0b;
    CCU2C _add_1_1433_add_4_4 (.A0(d3_adj_5742[2]), .B0(d2_adj_5741[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[3]), .B1(d2_adj_5741[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16222), .COUT(n16223), .S0(d3_71__N_562_adj_5758[2]), 
          .S1(d3_71__N_562_adj_5758[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1433_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1433_add_4_2 (.A0(d3_adj_5742[0]), .B0(d2_adj_5741[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[1]), .B1(d2_adj_5741[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16222), .S1(d3_71__N_562_adj_5758[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1433_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1433_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1433_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1433_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_37 (.A0(d7_adj_5747[70]), .B0(cout_adj_5613), 
          .C0(n81_adj_4953), .D0(n3_adj_4712), .A1(d7_adj_5747[71]), .B1(cout_adj_5613), 
          .C1(n78_adj_4952), .D1(n2_adj_4713), .CIN(n16219), .S0(d8_71__N_1603_adj_5774[70]), 
          .S1(d8_71__N_1603_adj_5774[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_35 (.A0(d7_adj_5747[68]), .B0(cout_adj_5613), 
          .C0(n87_adj_4955), .D0(n5_adj_4710), .A1(d7_adj_5747[69]), .B1(cout_adj_5613), 
          .C1(n84_adj_4954), .D1(n4_adj_4711), .CIN(n16218), .COUT(n16219), 
          .S0(d8_71__N_1603_adj_5774[68]), .S1(d8_71__N_1603_adj_5774[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_33 (.A0(d7_adj_5747[66]), .B0(cout_adj_5613), 
          .C0(n93_adj_4957), .D0(n7_adj_4708), .A1(d7_adj_5747[67]), .B1(cout_adj_5613), 
          .C1(n90_adj_4956), .D1(n6_adj_4709), .CIN(n16217), .COUT(n16218), 
          .S0(d8_71__N_1603_adj_5774[66]), .S1(d8_71__N_1603_adj_5774[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_31 (.A0(d7_adj_5747[64]), .B0(cout_adj_5613), 
          .C0(n99_adj_4959), .D0(n9_adj_4706), .A1(d7_adj_5747[65]), .B1(cout_adj_5613), 
          .C1(n96_adj_4958), .D1(n8_adj_4707), .CIN(n16216), .COUT(n16217), 
          .S0(d8_71__N_1603_adj_5774[64]), .S1(d8_71__N_1603_adj_5774[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_29 (.A0(d7_adj_5747[62]), .B0(cout_adj_5613), 
          .C0(n105_adj_4961), .D0(n11_adj_4704), .A1(d7_adj_5747[63]), 
          .B1(cout_adj_5613), .C1(n102_adj_4960), .D1(n10_adj_4705), .CIN(n16215), 
          .COUT(n16216), .S0(d8_71__N_1603_adj_5774[62]), .S1(d8_71__N_1603_adj_5774[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1474_add_4_27 (.A0(d7_adj_5747[60]), .B0(cout_adj_5613), 
          .C0(n111_adj_4963), .D0(n13_adj_4702), .A1(d7_adj_5747[61]), 
          .B1(cout_adj_5613), .C1(n108_adj_4962), .D1(n12_adj_4703), .CIN(n16214), 
          .COUT(n16215), .S0(d8_71__N_1603_adj_5774[60]), .S1(d8_71__N_1603_adj_5774[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1474_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1474_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1474_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1474_add_4_27.INJECT1_1 = "NO";
    LUT4 i3164_3_lut_4_lut (.A(led_c_0), .B(n17933), .C(n17094), .D(n12563), 
         .Z(n12983)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i3164_3_lut_4_lut.init = 16'hfe00;
    CCU2C _add_1_1519_add_4_15 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n147_adj_5312), .D0(d1[48]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n144_adj_5311), .D1(d1[49]), .CIN(n16186), .COUT(n16187), 
          .S0(d1_71__N_418[48]), .S1(d1_71__N_418[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_7 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n171_adj_5320), .D0(d1[40]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n168_adj_5319), .D1(d1[41]), .CIN(n16182), .COUT(n16183), 
          .S0(d1_71__N_418[40]), .S1(d1_71__N_418[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_7.INJECT1_1 = "NO";
    LUT4 mux_325_i27_4_lut (.A(n12112), .B(n241), .C(n17925), .D(n2572), 
         .Z(n2345)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i27_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1519_add_4_11 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n159_adj_5316), .D0(d1[44]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n156_adj_5315), .D1(d1[45]), .CIN(n16184), .COUT(n16185), 
          .S0(d1_71__N_418[44]), .S1(d1_71__N_418[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_11.INJECT1_1 = "NO";
    LUT4 i2358_3_lut_4_lut (.A(n18075), .B(n17937), .C(led_c_3), .D(n160_adj_5641), 
         .Z(n12156)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2358_3_lut_4_lut.init = 16'hf404;
    CCU2C _add_1_1436_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16176), .S0(cout_adj_5362));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1436_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1436_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_5 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n177_adj_5322), .D0(d1[38]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n174_adj_5321), .D1(d1[39]), .CIN(n16181), .COUT(n16182), 
          .S0(d1_71__N_418[38]), .S1(d1_71__N_418[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_5.INJECT1_1 = "NO";
    LUT4 i2348_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(n18076), .D(n178_adj_5647), 
         .Z(n12146)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2348_3_lut_4_lut.init = 16'hf404;
    CCU2C _add_1_1406_add_4_16 (.A0(d1[14]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[15]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16329), .COUT(n16330), .S0(d1_71__N_418[14]), 
          .S1(d1_71__N_418[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_36 (.A0(d4_adj_5743[34]), .B0(d3_adj_5742[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[35]), .B1(d3_adj_5742[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16175), .COUT(n16176), .S0(d4_71__N_634_adj_5759[34]), 
          .S1(d4_71__N_634_adj_5759[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_38 (.A0(d_d7[35]), .B0(d7[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16523), .S0(d8_71__N_1603[35]), .S1(cout_adj_5325));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1594_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_36 (.A0(d_d7[33]), .B0(d7[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[34]), .B1(d7[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16522), .COUT(n16523), .S0(d8_71__N_1603[33]), .S1(d8_71__N_1603[34]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_34 (.A0(d_d7[31]), .B0(d7[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[32]), .B1(d7[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16521), .COUT(n16522), .S0(d8_71__N_1603[31]), .S1(d8_71__N_1603[32]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_32 (.A0(d_d7[29]), .B0(d7[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[30]), .B1(d7[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16520), .COUT(n16521), .S0(d8_71__N_1603[29]), .S1(d8_71__N_1603[30]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_30 (.A0(d_d7[27]), .B0(d7[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[28]), .B1(d7[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16519), .COUT(n16520), .S0(d8_71__N_1603[27]), .S1(d8_71__N_1603[28]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_28 (.A0(d_d7[25]), .B0(d7[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[26]), .B1(d7[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16518), .COUT(n16519), .S0(d8_71__N_1603[25]), .S1(d8_71__N_1603[26]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_14 (.A0(d1[12]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[13]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16328), .COUT(n16329), .S0(d1_71__N_418[12]), 
          .S1(d1_71__N_418[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_34 (.A0(d4_adj_5743[32]), .B0(d3_adj_5742[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[33]), .B1(d3_adj_5742[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16174), .COUT(n16175), .S0(d4_71__N_634_adj_5759[32]), 
          .S1(d4_71__N_634_adj_5759[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_12 (.A0(d1[10]), .B0(MixerOutSin[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[11]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16327), .COUT(n16328), .S0(d1_71__N_418[10]), 
          .S1(d1_71__N_418[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_26 (.A0(d_d7[23]), .B0(d7[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[24]), .B1(d7[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16517), .COUT(n16518), .S0(d8_71__N_1603[23]), .S1(d8_71__N_1603[24]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_24 (.A0(d_d7[21]), .B0(d7[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[22]), .B1(d7[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16516), .COUT(n16517), .S0(d8_71__N_1603[21]), .S1(d8_71__N_1603[22]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_22 (.A0(d_d7[19]), .B0(d7[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[20]), .B1(d7[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16515), .COUT(n16516), .S0(d8_71__N_1603[19]), .S1(d8_71__N_1603[20]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_20 (.A0(d_d7[17]), .B0(d7[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[18]), .B1(d7[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16514), .COUT(n16515), .S0(d8_71__N_1603[17]), .S1(d8_71__N_1603[18]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_18 (.A0(d_d7[15]), .B0(d7[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[16]), .B1(d7[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16513), .COUT(n16514), .S0(d8_71__N_1603[15]), .S1(d8_71__N_1603[16]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_16 (.A0(d_d7[13]), .B0(d7[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[14]), .B1(d7[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16512), .COUT(n16513), .S0(d8_71__N_1603[13]), .S1(d8_71__N_1603[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_14 (.A0(d_d7[11]), .B0(d7[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[12]), .B1(d7[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16511), .COUT(n16512), .S0(d8_71__N_1603[11]), .S1(d8_71__N_1603[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_12 (.A0(d_d7[9]), .B0(d7[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[10]), .B1(d7[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16510), .COUT(n16511), .S0(d8_71__N_1603[9]), .S1(d8_71__N_1603[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_10 (.A0(d_d7[7]), .B0(d7[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[8]), .B1(d7[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16509), .COUT(n16510), .S0(d8_71__N_1603[7]), .S1(d8_71__N_1603[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_8 (.A0(d_d7[5]), .B0(d7[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[6]), .B1(d7[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16508), .COUT(n16509), .S0(d8_71__N_1603[5]), .S1(d8_71__N_1603[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_6 (.A0(d_d7[3]), .B0(d7[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[4]), .B1(d7[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16507), .COUT(n16508), .S0(d8_71__N_1603[3]), .S1(d8_71__N_1603[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_4 (.A0(d_d7[1]), .B0(d7[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[2]), .B1(d7[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16506), .COUT(n16507), .S0(d8_71__N_1603[1]), .S1(d8_71__N_1603[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1594_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1594_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[0]), .B1(d7[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16506), .S1(d8_71__N_1603[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1594_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1594_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1594_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1594_add_4_2.INJECT1_1 = "NO";
    FD1P3AX CICGain__i2 (.D(led_c_1), .SP(clk_80mhz_enable_1407), .CK(clk_80mhz), 
            .Q(CICGain[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam CICGain__i2.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i2 (.D(n123_adj_5441), .CK(CIC1_out_clkSin), .Q(ISquare[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i2.GSR = "ENABLED";
    CCU2C _add_1_1436_add_4_32 (.A0(d4_adj_5743[30]), .B0(d3_adj_5742[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[31]), .B1(d3_adj_5742[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16173), .COUT(n16174), .S0(d4_71__N_634_adj_5759[30]), 
          .S1(d4_71__N_634_adj_5759[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_37 (.A0(d1_adj_5740[70]), .B0(cout_adj_5344), 
          .C0(n81), .D0(d2_adj_5741[70]), .A1(d1_adj_5740[71]), .B1(cout_adj_5344), 
          .C1(n78), .D1(d2_adj_5741[71]), .CIN(n16504), .S0(d2_71__N_490_adj_5757[70]), 
          .S1(d2_71__N_490_adj_5757[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_37.INJECT1_1 = "NO";
    FD1S3AX ISquare_e3__i3 (.D(n120_adj_5440), .CK(CIC1_out_clkSin), .Q(ISquare[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i3.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i4 (.D(n117_adj_5439), .CK(CIC1_out_clkSin), .Q(ISquare[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i4.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i5 (.D(n114_adj_5438), .CK(CIC1_out_clkSin), .Q(ISquare[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i5.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i6 (.D(n111_adj_5437), .CK(CIC1_out_clkSin), .Q(ISquare[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i6.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i7 (.D(n108_adj_5436), .CK(CIC1_out_clkSin), .Q(ISquare[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i7.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i8 (.D(n105_adj_5435), .CK(CIC1_out_clkSin), .Q(ISquare[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i8.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i9 (.D(n102_adj_5434), .CK(CIC1_out_clkSin), .Q(ISquare[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i9.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i10 (.D(n99_adj_5433), .CK(CIC1_out_clkSin), .Q(ISquare[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i10.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i11 (.D(n96_adj_5432), .CK(CIC1_out_clkSin), .Q(ISquare[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i11.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i12 (.D(n93_adj_5431), .CK(CIC1_out_clkSin), .Q(ISquare[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i12.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i13 (.D(n90_adj_5430), .CK(CIC1_out_clkSin), .Q(ISquare[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i13.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i14 (.D(n87_adj_5429), .CK(CIC1_out_clkSin), .Q(ISquare[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i14.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i15 (.D(n84_adj_5428), .CK(CIC1_out_clkSin), .Q(ISquare[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i15.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i16 (.D(n81_adj_5427), .CK(CIC1_out_clkSin), .Q(ISquare[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i16.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i17 (.D(n78_adj_5426), .CK(CIC1_out_clkSin), .Q(ISquare[16]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i17.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i18 (.D(n75_adj_5425), .CK(CIC1_out_clkSin), .Q(ISquare[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i18.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i19 (.D(n72_adj_5424), .CK(CIC1_out_clkSin), .Q(ISquare[18]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i19.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i20 (.D(n69_adj_5423), .CK(CIC1_out_clkSin), .Q(ISquare[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i20.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i21 (.D(n66_adj_5422), .CK(CIC1_out_clkSin), .Q(ISquare[20]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i21.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i22 (.D(n63_adj_5421), .CK(CIC1_out_clkSin), .Q(ISquare[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i22.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i23 (.D(n60_adj_5420), .CK(CIC1_out_clkSin), .Q(ISquare[22]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i23.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i24 (.D(n57_adj_5419), .CK(CIC1_out_clkSin), .Q(ISquare[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i24.GSR = "ENABLED";
    FD1S3AX ISquare_e3__i25 (.D(n54_adj_5418), .CK(CIC1_out_clkSin), .Q(ISquare[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_e3__i25.GSR = "ENABLED";
    CCU2C _add_1_1406_add_4_10 (.A0(d1[8]), .B0(MixerOutSin[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[9]), .B1(MixerOutSin[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16326), .COUT(n16327), .S0(d1_71__N_418[8]), 
          .S1(d1_71__N_418[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_34 (.A0(d_d6_adj_5746[31]), .B0(d6_adj_5745[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[32]), .B1(d6_adj_5745[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16078), .COUT(n16079), .S0(d7_71__N_1531_adj_5773[31]), 
          .S1(d7_71__N_1531_adj_5773[32]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_35 (.A0(d1_adj_5740[68]), .B0(cout_adj_5344), 
          .C0(n87), .D0(d2_adj_5741[68]), .A1(d1_adj_5740[69]), .B1(cout_adj_5344), 
          .C1(n84), .D1(d2_adj_5741[69]), .CIN(n16503), .COUT(n16504), 
          .S0(d2_71__N_490_adj_5757[68]), .S1(d2_71__N_490_adj_5757[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_33 (.A0(d1_adj_5740[66]), .B0(cout_adj_5344), 
          .C0(n93), .D0(d2_adj_5741[66]), .A1(d1_adj_5740[67]), .B1(cout_adj_5344), 
          .C1(n90), .D1(d2_adj_5741[67]), .CIN(n16502), .COUT(n16503), 
          .S0(d2_71__N_490_adj_5757[66]), .S1(d2_71__N_490_adj_5757[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_31 (.A0(d1_adj_5740[64]), .B0(cout_adj_5344), 
          .C0(n99), .D0(d2_adj_5741[64]), .A1(d1_adj_5740[65]), .B1(cout_adj_5344), 
          .C1(n96), .D1(d2_adj_5741[65]), .CIN(n16501), .COUT(n16502), 
          .S0(d2_71__N_490_adj_5757[64]), .S1(d2_71__N_490_adj_5757[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_29 (.A0(d1_adj_5740[62]), .B0(cout_adj_5344), 
          .C0(n105), .D0(d2_adj_5741[62]), .A1(d1_adj_5740[63]), .B1(cout_adj_5344), 
          .C1(n102), .D1(d2_adj_5741[63]), .CIN(n16500), .COUT(n16501), 
          .S0(d2_71__N_490_adj_5757[62]), .S1(d2_71__N_490_adj_5757[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_27 (.A0(d1_adj_5740[60]), .B0(cout_adj_5344), 
          .C0(n111), .D0(d2_adj_5741[60]), .A1(d1_adj_5740[61]), .B1(cout_adj_5344), 
          .C1(n108), .D1(d2_adj_5741[61]), .CIN(n16499), .COUT(n16500), 
          .S0(d2_71__N_490_adj_5757[60]), .S1(d2_71__N_490_adj_5757[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_25 (.A0(d1_adj_5740[58]), .B0(cout_adj_5344), 
          .C0(n117), .D0(d2_adj_5741[58]), .A1(d1_adj_5740[59]), .B1(cout_adj_5344), 
          .C1(n114), .D1(d2_adj_5741[59]), .CIN(n16498), .COUT(n16499), 
          .S0(d2_71__N_490_adj_5757[58]), .S1(d2_71__N_490_adj_5757[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_23 (.A0(d1_adj_5740[56]), .B0(cout_adj_5344), 
          .C0(n123), .D0(d2_adj_5741[56]), .A1(d1_adj_5740[57]), .B1(cout_adj_5344), 
          .C1(n120), .D1(d2_adj_5741[57]), .CIN(n16497), .COUT(n16498), 
          .S0(d2_71__N_490_adj_5757[56]), .S1(d2_71__N_490_adj_5757[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_21 (.A0(d1_adj_5740[54]), .B0(cout_adj_5344), 
          .C0(n129), .D0(d2_adj_5741[54]), .A1(d1_adj_5740[55]), .B1(cout_adj_5344), 
          .C1(n126), .D1(d2_adj_5741[55]), .CIN(n16496), .COUT(n16497), 
          .S0(d2_71__N_490_adj_5757[54]), .S1(d2_71__N_490_adj_5757[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_19 (.A0(d1_adj_5740[52]), .B0(cout_adj_5344), 
          .C0(n135), .D0(d2_adj_5741[52]), .A1(d1_adj_5740[53]), .B1(cout_adj_5344), 
          .C1(n132), .D1(d2_adj_5741[53]), .CIN(n16495), .COUT(n16496), 
          .S0(d2_71__N_490_adj_5757[52]), .S1(d2_71__N_490_adj_5757[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1436_add_4_30 (.A0(d4_adj_5743[28]), .B0(d3_adj_5742[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[29]), .B1(d3_adj_5742[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16172), .COUT(n16173), .S0(d4_71__N_634_adj_5759[28]), 
          .S1(d4_71__N_634_adj_5759[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1436_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1436_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1436_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1436_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16117), .S0(cout_adj_5363));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1439_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1439_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_17 (.A0(d1_adj_5740[50]), .B0(cout_adj_5344), 
          .C0(n141), .D0(d2_adj_5741[50]), .A1(d1_adj_5740[51]), .B1(cout_adj_5344), 
          .C1(n138), .D1(d2_adj_5741[51]), .CIN(n16494), .COUT(n16495), 
          .S0(d2_71__N_490_adj_5757[50]), .S1(d2_71__N_490_adj_5757[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_36 (.A0(d5_adj_5744[34]), .B0(d4_adj_5743[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[35]), .B1(d4_adj_5743[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16116), .COUT(n16117), .S0(d5_71__N_706_adj_5760[34]), 
          .S1(d5_71__N_706_adj_5760[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_8 (.A0(d1[6]), .B0(MixerOutSin[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[7]), .B1(MixerOutSin[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16325), .COUT(n16326), .S0(d1_71__N_418[6]), 
          .S1(d1_71__N_418[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_34 (.A0(d5_adj_5744[32]), .B0(d4_adj_5743[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[33]), .B1(d4_adj_5743[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16115), .COUT(n16116), .S0(d5_71__N_706_adj_5760[32]), 
          .S1(d5_71__N_706_adj_5760[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_32 (.A0(d5_adj_5744[30]), .B0(d4_adj_5743[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[31]), .B1(d4_adj_5743[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16114), .COUT(n16115), .S0(d5_71__N_706_adj_5760[30]), 
          .S1(d5_71__N_706_adj_5760[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_32 (.A0(d_d6_adj_5746[29]), .B0(d6_adj_5745[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[30]), .B1(d6_adj_5745[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16077), .COUT(n16078), .S0(d7_71__N_1531_adj_5773[29]), 
          .S1(d7_71__N_1531_adj_5773[30]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_30 (.A0(d_d6_adj_5746[27]), .B0(d6_adj_5745[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[28]), .B1(d6_adj_5745[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16076), .COUT(n16077), .S0(d7_71__N_1531_adj_5773[27]), 
          .S1(d7_71__N_1531_adj_5773[28]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_28 (.A0(d_d6_adj_5746[25]), .B0(d6_adj_5745[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[26]), .B1(d6_adj_5745[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16075), .COUT(n16076), .S0(d7_71__N_1531_adj_5773[25]), 
          .S1(d7_71__N_1531_adj_5773[26]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_26 (.A0(d_d6_adj_5746[23]), .B0(d6_adj_5745[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[24]), .B1(d6_adj_5745[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16074), .COUT(n16075), .S0(d7_71__N_1531_adj_5773[23]), 
          .S1(d7_71__N_1531_adj_5773[24]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_24 (.A0(d_d6_adj_5746[21]), .B0(d6_adj_5745[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[22]), .B1(d6_adj_5745[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16073), .COUT(n16074), .S0(d7_71__N_1531_adj_5773[21]), 
          .S1(d7_71__N_1531_adj_5773[22]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_22 (.A0(d_d6_adj_5746[19]), .B0(d6_adj_5745[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[20]), .B1(d6_adj_5745[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16072), .COUT(n16073), .S0(d7_71__N_1531_adj_5773[19]), 
          .S1(d7_71__N_1531_adj_5773[20]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_20 (.A0(d_d6_adj_5746[17]), .B0(d6_adj_5745[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[18]), .B1(d6_adj_5745[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16071), .COUT(n16072), .S0(d7_71__N_1531_adj_5773[17]), 
          .S1(d7_71__N_1531_adj_5773[18]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_18 (.A0(d_d6_adj_5746[15]), .B0(d6_adj_5745[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[16]), .B1(d6_adj_5745[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16070), .COUT(n16071), .S0(d7_71__N_1531_adj_5773[15]), 
          .S1(d7_71__N_1531_adj_5773[16]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_16 (.A0(d_d6_adj_5746[13]), .B0(d6_adj_5745[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[14]), .B1(d6_adj_5745[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16069), .COUT(n16070), .S0(d7_71__N_1531_adj_5773[13]), 
          .S1(d7_71__N_1531_adj_5773[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_14 (.A0(d_d6_adj_5746[11]), .B0(d6_adj_5745[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[12]), .B1(d6_adj_5745[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16068), .COUT(n16069), .S0(d7_71__N_1531_adj_5773[11]), 
          .S1(d7_71__N_1531_adj_5773[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_12 (.A0(d_d6_adj_5746[9]), .B0(d6_adj_5745[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[10]), .B1(d6_adj_5745[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16067), .COUT(n16068), .S0(d7_71__N_1531_adj_5773[9]), 
          .S1(d7_71__N_1531_adj_5773[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_10 (.A0(d_d6_adj_5746[7]), .B0(d6_adj_5745[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[8]), .B1(d6_adj_5745[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16066), .COUT(n16067), .S0(d7_71__N_1531_adj_5773[7]), 
          .S1(d7_71__N_1531_adj_5773[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_8 (.A0(d_d6_adj_5746[5]), .B0(d6_adj_5745[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[6]), .B1(d6_adj_5745[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16065), .COUT(n16066), .S0(d7_71__N_1531_adj_5773[5]), 
          .S1(d7_71__N_1531_adj_5773[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_6 (.A0(d_d6_adj_5746[3]), .B0(d6_adj_5745[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[4]), .B1(d6_adj_5745[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16064), .COUT(n16065), .S0(d7_71__N_1531_adj_5773[3]), 
          .S1(d7_71__N_1531_adj_5773[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_4 (.A0(d_d6_adj_5746[1]), .B0(d6_adj_5745[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[2]), .B1(d6_adj_5745[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16063), .COUT(n16064), .S0(d7_71__N_1531_adj_5773[1]), 
          .S1(d7_71__N_1531_adj_5773[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1615_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1615_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6_adj_5746[0]), .B1(d6_adj_5745[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16063), .S1(d7_71__N_1531_adj_5773[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1615_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1615_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1615_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1615_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_38 (.A0(d3_adj_5742[71]), .B0(d2_adj_5741[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16062), .S0(n78_adj_5114));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1576_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_36 (.A0(d3_adj_5742[69]), .B0(d2_adj_5741[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[70]), .B1(d2_adj_5741[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16061), .COUT(n16062), .S0(n84_adj_5116), 
          .S1(n81_adj_5115));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_34 (.A0(d3_adj_5742[67]), .B0(d2_adj_5741[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[68]), .B1(d2_adj_5741[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16060), .COUT(n16061), .S0(n90_adj_5118), 
          .S1(n87_adj_5117));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_32 (.A0(d3_adj_5742[65]), .B0(d2_adj_5741[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[66]), .B1(d2_adj_5741[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16059), .COUT(n16060), .S0(n96_adj_5120), 
          .S1(n93_adj_5119));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_30 (.A0(d3_adj_5742[63]), .B0(d2_adj_5741[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[64]), .B1(d2_adj_5741[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16058), .COUT(n16059), .S0(n102_adj_5122), 
          .S1(n99_adj_5121));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_28 (.A0(d3_adj_5742[61]), .B0(d2_adj_5741[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[62]), .B1(d2_adj_5741[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16057), .COUT(n16058), .S0(n108_adj_5124), 
          .S1(n105_adj_5123));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_26 (.A0(d3_adj_5742[59]), .B0(d2_adj_5741[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[60]), .B1(d2_adj_5741[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16056), .COUT(n16057), .S0(n114_adj_5126), 
          .S1(n111_adj_5125));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_24 (.A0(d3_adj_5742[57]), .B0(d2_adj_5741[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[58]), .B1(d2_adj_5741[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16055), .COUT(n16056), .S0(n120_adj_5128), 
          .S1(n117_adj_5127));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_22 (.A0(d3_adj_5742[55]), .B0(d2_adj_5741[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[56]), .B1(d2_adj_5741[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16054), .COUT(n16055), .S0(n126_adj_5130), 
          .S1(n123_adj_5129));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_20 (.A0(d3_adj_5742[53]), .B0(d2_adj_5741[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[54]), .B1(d2_adj_5741[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16053), .COUT(n16054), .S0(n132_adj_5132), 
          .S1(n129_adj_5131));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_18 (.A0(d3_adj_5742[51]), .B0(d2_adj_5741[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[52]), .B1(d2_adj_5741[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16052), .COUT(n16053), .S0(n138_adj_5134), 
          .S1(n135_adj_5133));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_16 (.A0(d3_adj_5742[49]), .B0(d2_adj_5741[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[50]), .B1(d2_adj_5741[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16051), .COUT(n16052), .S0(n144_adj_5136), 
          .S1(n141_adj_5135));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_14 (.A0(d3_adj_5742[47]), .B0(d2_adj_5741[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[48]), .B1(d2_adj_5741[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16050), .COUT(n16051), .S0(n150_adj_5138), 
          .S1(n147_adj_5137));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_12 (.A0(d3_adj_5742[45]), .B0(d2_adj_5741[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[46]), .B1(d2_adj_5741[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16049), .COUT(n16050), .S0(n156_adj_5140), 
          .S1(n153_adj_5139));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_10 (.A0(d3_adj_5742[43]), .B0(d2_adj_5741[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[44]), .B1(d2_adj_5741[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16048), .COUT(n16049), .S0(n162_adj_5142), 
          .S1(n159_adj_5141));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_8 (.A0(d3_adj_5742[41]), .B0(d2_adj_5741[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[42]), .B1(d2_adj_5741[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16047), .COUT(n16048), .S0(n168_adj_5144), 
          .S1(n165_adj_5143));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_6 (.A0(d3_adj_5742[39]), .B0(d2_adj_5741[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[40]), .B1(d2_adj_5741[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16046), .COUT(n16047), .S0(n174_adj_5146), 
          .S1(n171_adj_5145));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_4 (.A0(d3_adj_5742[37]), .B0(d2_adj_5741[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d3_adj_5742[38]), .B1(d2_adj_5741[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16045), .COUT(n16046), .S0(n180_adj_5148), 
          .S1(n177_adj_5147));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1576_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1576_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d3_adj_5742[36]), .B1(d2_adj_5741[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16045), .S1(n183_adj_5149));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1576_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1576_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1576_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1576_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_38 (.A0(d4_adj_5743[71]), .B0(d3_adj_5742[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16044), .S0(n78_adj_5150));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1579_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_36 (.A0(d4_adj_5743[69]), .B0(d3_adj_5742[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[70]), .B1(d3_adj_5742[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16043), .COUT(n16044), .S0(n84_adj_5152), 
          .S1(n81_adj_5151));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_34 (.A0(d4_adj_5743[67]), .B0(d3_adj_5742[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[68]), .B1(d3_adj_5742[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16042), .COUT(n16043), .S0(n90_adj_5154), 
          .S1(n87_adj_5153));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_32 (.A0(d4_adj_5743[65]), .B0(d3_adj_5742[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[66]), .B1(d3_adj_5742[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16041), .COUT(n16042), .S0(n96_adj_5156), 
          .S1(n93_adj_5155));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_30 (.A0(d4_adj_5743[63]), .B0(d3_adj_5742[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[64]), .B1(d3_adj_5742[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16040), .COUT(n16041), .S0(n102_adj_5158), 
          .S1(n99_adj_5157));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_28 (.A0(d4_adj_5743[61]), .B0(d3_adj_5742[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[62]), .B1(d3_adj_5742[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16039), .COUT(n16040), .S0(n108_adj_5160), 
          .S1(n105_adj_5159));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_26 (.A0(d4_adj_5743[59]), .B0(d3_adj_5742[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[60]), .B1(d3_adj_5742[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16038), .COUT(n16039), .S0(n114_adj_5162), 
          .S1(n111_adj_5161));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_24 (.A0(d4_adj_5743[57]), .B0(d3_adj_5742[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[58]), .B1(d3_adj_5742[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16037), .COUT(n16038), .S0(n120_adj_5164), 
          .S1(n117_adj_5163));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_22 (.A0(d4_adj_5743[55]), .B0(d3_adj_5742[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[56]), .B1(d3_adj_5742[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16036), .COUT(n16037), .S0(n126_adj_5166), 
          .S1(n123_adj_5165));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_20 (.A0(d4_adj_5743[53]), .B0(d3_adj_5742[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[54]), .B1(d3_adj_5742[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16035), .COUT(n16036), .S0(n132_adj_5168), 
          .S1(n129_adj_5167));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_18 (.A0(d4_adj_5743[51]), .B0(d3_adj_5742[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[52]), .B1(d3_adj_5742[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16034), .COUT(n16035), .S0(n138_adj_5170), 
          .S1(n135_adj_5169));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_16 (.A0(d4_adj_5743[49]), .B0(d3_adj_5742[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[50]), .B1(d3_adj_5742[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16033), .COUT(n16034), .S0(n144_adj_5172), 
          .S1(n141_adj_5171));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_14 (.A0(d4_adj_5743[47]), .B0(d3_adj_5742[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[48]), .B1(d3_adj_5742[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16032), .COUT(n16033), .S0(n150_adj_5174), 
          .S1(n147_adj_5173));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_12 (.A0(d4_adj_5743[45]), .B0(d3_adj_5742[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[46]), .B1(d3_adj_5742[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16031), .COUT(n16032), .S0(n156_adj_5176), 
          .S1(n153_adj_5175));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_10 (.A0(d4_adj_5743[43]), .B0(d3_adj_5742[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[44]), .B1(d3_adj_5742[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16030), .COUT(n16031), .S0(n162_adj_5178), 
          .S1(n159_adj_5177));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_8 (.A0(d4_adj_5743[41]), .B0(d3_adj_5742[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[42]), .B1(d3_adj_5742[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16029), .COUT(n16030), .S0(n168_adj_5180), 
          .S1(n165_adj_5179));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_6 (.A0(d4_adj_5743[39]), .B0(d3_adj_5742[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[40]), .B1(d3_adj_5742[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16028), .COUT(n16029), .S0(n174_adj_5182), 
          .S1(n171_adj_5181));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_4 (.A0(d4_adj_5743[37]), .B0(d3_adj_5742[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d4_adj_5743[38]), .B1(d3_adj_5742[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16027), .COUT(n16028), .S0(n180_adj_5184), 
          .S1(n177_adj_5183));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1579_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1579_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d4_adj_5743[36]), .B1(d3_adj_5742[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16027), .S1(n183_adj_5185));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1579_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1579_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1579_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1579_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_38 (.A0(d5_adj_5744[71]), .B0(d4_adj_5743[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16026), .S0(n78_adj_5188));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1582_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_36 (.A0(d5_adj_5744[69]), .B0(d4_adj_5743[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[70]), .B1(d4_adj_5743[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16025), .COUT(n16026), .S0(n84_adj_5190), 
          .S1(n81_adj_5189));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_34 (.A0(d5_adj_5744[67]), .B0(d4_adj_5743[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[68]), .B1(d4_adj_5743[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16024), .COUT(n16025), .S0(n90_adj_5192), 
          .S1(n87_adj_5191));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_32 (.A0(d5_adj_5744[65]), .B0(d4_adj_5743[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[66]), .B1(d4_adj_5743[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16023), .COUT(n16024), .S0(n96_adj_5194), 
          .S1(n93_adj_5193));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_30 (.A0(d5_adj_5744[63]), .B0(d4_adj_5743[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[64]), .B1(d4_adj_5743[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16022), .COUT(n16023), .S0(n102_adj_5196), 
          .S1(n99_adj_5195));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_28 (.A0(d5_adj_5744[61]), .B0(d4_adj_5743[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[62]), .B1(d4_adj_5743[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16021), .COUT(n16022), .S0(n108_adj_5198), 
          .S1(n105_adj_5197));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_26 (.A0(d5_adj_5744[59]), .B0(d4_adj_5743[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[60]), .B1(d4_adj_5743[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16020), .COUT(n16021), .S0(n114_adj_5200), 
          .S1(n111_adj_5199));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_24 (.A0(d5_adj_5744[57]), .B0(d4_adj_5743[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[58]), .B1(d4_adj_5743[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16019), .COUT(n16020), .S0(n120_adj_5202), 
          .S1(n117_adj_5201));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_22 (.A0(d5_adj_5744[55]), .B0(d4_adj_5743[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[56]), .B1(d4_adj_5743[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16018), .COUT(n16019), .S0(n126_adj_5204), 
          .S1(n123_adj_5203));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_20 (.A0(d5_adj_5744[53]), .B0(d4_adj_5743[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[54]), .B1(d4_adj_5743[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16017), .COUT(n16018), .S0(n132_adj_5206), 
          .S1(n129_adj_5205));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_18 (.A0(d5_adj_5744[51]), .B0(d4_adj_5743[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[52]), .B1(d4_adj_5743[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16016), .COUT(n16017), .S0(n138_adj_5208), 
          .S1(n135_adj_5207));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_16 (.A0(d5_adj_5744[49]), .B0(d4_adj_5743[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[50]), .B1(d4_adj_5743[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16015), .COUT(n16016), .S0(n144_adj_5210), 
          .S1(n141_adj_5209));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_14 (.A0(d5_adj_5744[47]), .B0(d4_adj_5743[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[48]), .B1(d4_adj_5743[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16014), .COUT(n16015), .S0(n150_adj_5212), 
          .S1(n147_adj_5211));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_12 (.A0(d5_adj_5744[45]), .B0(d4_adj_5743[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[46]), .B1(d4_adj_5743[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16013), .COUT(n16014), .S0(n156_adj_5214), 
          .S1(n153_adj_5213));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_10 (.A0(d5_adj_5744[43]), .B0(d4_adj_5743[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[44]), .B1(d4_adj_5743[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16012), .COUT(n16013), .S0(n162_adj_5216), 
          .S1(n159_adj_5215));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_8 (.A0(d5_adj_5744[41]), .B0(d4_adj_5743[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[42]), .B1(d4_adj_5743[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16011), .COUT(n16012), .S0(n168_adj_5218), 
          .S1(n165_adj_5217));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_6 (.A0(d5_adj_5744[39]), .B0(d4_adj_5743[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[40]), .B1(d4_adj_5743[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16010), .COUT(n16011), .S0(n174_adj_5220), 
          .S1(n171_adj_5219));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_4 (.A0(d5_adj_5744[37]), .B0(d4_adj_5743[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[38]), .B1(d4_adj_5743[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16009), .COUT(n16010), .S0(n180_adj_5222), 
          .S1(n177_adj_5221));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1582_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1582_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d5_adj_5744[36]), .B1(d4_adj_5743[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16009), .S1(n183_adj_5223));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1582_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1582_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1582_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1582_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_38 (.A0(d_d8_adj_5750[71]), .B0(d8_adj_5749[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16008), .S0(n78_adj_4988));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1639_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1480_add_4_9 (.A0(d_tmp_adj_5738[42]), .B0(cout_adj_5605), 
          .C0(n165_adj_4909), .D0(n31_adj_2808), .A1(d_tmp_adj_5738[43]), 
          .B1(cout_adj_5605), .C1(n162_adj_4908), .D1(n30_adj_2809), .CIN(n15862), 
          .COUT(n15863), .S0(d6_71__N_1459_adj_5772[42]), .S1(d6_71__N_1459_adj_5772[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1480_add_4_7 (.A0(d_tmp_adj_5738[40]), .B0(cout_adj_5605), 
          .C0(n171_adj_4911), .D0(n33), .A1(d_tmp_adj_5738[41]), .B1(cout_adj_5605), 
          .C1(n168_adj_4910), .D1(n32), .CIN(n15861), .COUT(n15862), 
          .S0(d6_71__N_1459_adj_5772[40]), .S1(d6_71__N_1459_adj_5772[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1480_add_4_5 (.A0(d_tmp_adj_5738[38]), .B0(cout_adj_5605), 
          .C0(n177_adj_4913), .D0(n35), .A1(d_tmp_adj_5738[39]), .B1(cout_adj_5605), 
          .C1(n174_adj_4912), .D1(n34), .CIN(n15860), .COUT(n15861), 
          .S0(d6_71__N_1459_adj_5772[38]), .S1(d6_71__N_1459_adj_5772[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1480_add_4_3 (.A0(d_tmp_adj_5738[36]), .B0(cout_adj_5605), 
          .C0(n183_adj_4915), .D0(n37), .A1(d_tmp_adj_5738[37]), .B1(cout_adj_5605), 
          .C1(n180_adj_4914), .D1(n36), .CIN(n15859), .COUT(n15860), 
          .S0(d6_71__N_1459_adj_5772[36]), .S1(d6_71__N_1459_adj_5772[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1480_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1480_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1480_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5605), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15859));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1480_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1480_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1480_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1480_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_38 (.A0(d4[71]), .B0(d3[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15855), .S0(n78_adj_5689));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1564_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_36 (.A0(d4[69]), .B0(d3[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[70]), .B1(d3[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15854), .COUT(n15855), .S0(n84_adj_5691), .S1(n81_adj_5690));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_34 (.A0(d4[67]), .B0(d3[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[68]), .B1(d3[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15853), .COUT(n15854), .S0(n90_adj_5693), .S1(n87_adj_5692));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_32 (.A0(d4[65]), .B0(d3[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[66]), .B1(d3[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15852), .COUT(n15853), .S0(n96_adj_5695), .S1(n93_adj_5694));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_30 (.A0(d4[63]), .B0(d3[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[64]), .B1(d3[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15851), .COUT(n15852), .S0(n102_adj_5697), .S1(n99_adj_5696));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_28 (.A0(d4[61]), .B0(d3[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[62]), .B1(d3[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15850), .COUT(n15851), .S0(n108_adj_5699), .S1(n105_adj_5698));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_26 (.A0(d4[59]), .B0(d3[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[60]), .B1(d3[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15849), .COUT(n15850), .S0(n114_adj_5701), .S1(n111_adj_5700));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_24 (.A0(d4[57]), .B0(d3[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[58]), .B1(d3[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15848), .COUT(n15849), .S0(n120_adj_5703), .S1(n117_adj_5702));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_22 (.A0(d4[55]), .B0(d3[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[56]), .B1(d3[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15847), .COUT(n15848), .S0(n126_adj_5705), .S1(n123_adj_5704));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_20 (.A0(d4[53]), .B0(d3[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[54]), .B1(d3[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15846), .COUT(n15847), .S0(n132_adj_5707), .S1(n129_adj_5706));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_18 (.A0(d4[51]), .B0(d3[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[52]), .B1(d3[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15845), .COUT(n15846), .S0(n138_adj_5709), .S1(n135_adj_5708));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_16 (.A0(d4[49]), .B0(d3[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[50]), .B1(d3[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15844), .COUT(n15845), .S0(n144_adj_5711), .S1(n141_adj_5710));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_14 (.A0(d4[47]), .B0(d3[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[48]), .B1(d3[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15843), .COUT(n15844), .S0(n150_adj_5713), .S1(n147_adj_5712));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_12 (.A0(d4[45]), .B0(d3[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[46]), .B1(d3[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15842), .COUT(n15843), .S0(n156_adj_5715), .S1(n153_adj_5714));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_10 (.A0(d4[43]), .B0(d3[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[44]), .B1(d3[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15841), .COUT(n15842), .S0(n162_adj_5717), .S1(n159_adj_5716));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_8 (.A0(d4[41]), .B0(d3[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[42]), .B1(d3[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15840), .COUT(n15841), .S0(n168_adj_5719), .S1(n165_adj_5718));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_6 (.A0(d4[39]), .B0(d3[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[40]), .B1(d3[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15839), .COUT(n15840), .S0(n174_adj_5721), .S1(n171_adj_5720));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_4 (.A0(d4[37]), .B0(d3[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[38]), .B1(d3[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15838), .COUT(n15839), .S0(n180_adj_5723), .S1(n177_adj_5722));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1564_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1564_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[36]), .B1(d3[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15838), .S1(n183_adj_5724));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1564_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1564_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1564_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1564_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_37 (.A0(d6[70]), .B0(cout_adj_5443), .C0(n81_adj_5076), 
          .D0(n3_adj_4626), .A1(d6[71]), .B1(cout_adj_5443), .C1(n78_adj_5075), 
          .D1(n2_adj_4627), .CIN(n15836), .S0(d7_71__N_1531[70]), .S1(d7_71__N_1531[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_35 (.A0(d6[68]), .B0(cout_adj_5443), .C0(n87_adj_5078), 
          .D0(n5_adj_4789), .A1(d6[69]), .B1(cout_adj_5443), .C1(n84_adj_5077), 
          .D1(n4_adj_4790), .CIN(n15835), .COUT(n15836), .S0(d7_71__N_1531[68]), 
          .S1(d7_71__N_1531[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_33 (.A0(d6[66]), .B0(cout_adj_5443), .C0(n93_adj_5080), 
          .D0(n7_adj_4787), .A1(d6[67]), .B1(cout_adj_5443), .C1(n90_adj_5079), 
          .D1(n6_adj_4788), .CIN(n15834), .COUT(n15835), .S0(d7_71__N_1531[66]), 
          .S1(d7_71__N_1531[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_31 (.A0(d6[64]), .B0(cout_adj_5443), .C0(n99_adj_5082), 
          .D0(n9_adj_4785), .A1(d6[65]), .B1(cout_adj_5443), .C1(n96_adj_5081), 
          .D1(n8_adj_4786), .CIN(n15833), .COUT(n15834), .S0(d7_71__N_1531[64]), 
          .S1(d7_71__N_1531[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_29 (.A0(d6[62]), .B0(cout_adj_5443), .C0(n105_adj_5084), 
          .D0(n11_adj_4783), .A1(d6[63]), .B1(cout_adj_5443), .C1(n102_adj_5083), 
          .D1(n10_adj_4784), .CIN(n15832), .COUT(n15833), .S0(d7_71__N_1531[62]), 
          .S1(d7_71__N_1531[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_27 (.A0(d6[60]), .B0(cout_adj_5443), .C0(n111_adj_5086), 
          .D0(n13_adj_4781), .A1(d6[61]), .B1(cout_adj_5443), .C1(n108_adj_5085), 
          .D1(n12_adj_4782), .CIN(n15831), .COUT(n15832), .S0(d7_71__N_1531[60]), 
          .S1(d7_71__N_1531[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_25 (.A0(d6[58]), .B0(cout_adj_5443), .C0(n117_adj_5088), 
          .D0(n15_adj_4779), .A1(d6[59]), .B1(cout_adj_5443), .C1(n114_adj_5087), 
          .D1(n14_adj_4780), .CIN(n15830), .COUT(n15831), .S0(d7_71__N_1531[58]), 
          .S1(d7_71__N_1531[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_23 (.A0(d6[56]), .B0(cout_adj_5443), .C0(n123_adj_5090), 
          .D0(n17_adj_4777), .A1(d6[57]), .B1(cout_adj_5443), .C1(n120_adj_5089), 
          .D1(n16_adj_4778), .CIN(n15829), .COUT(n15830), .S0(d7_71__N_1531[56]), 
          .S1(d7_71__N_1531[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_21 (.A0(d6[54]), .B0(cout_adj_5443), .C0(n129_adj_5092), 
          .D0(n19_adj_4775), .A1(d6[55]), .B1(cout_adj_5443), .C1(n126_adj_5091), 
          .D1(n18_adj_4776), .CIN(n15828), .COUT(n15829), .S0(d7_71__N_1531[54]), 
          .S1(d7_71__N_1531[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_19 (.A0(d6[52]), .B0(cout_adj_5443), .C0(n135_adj_5094), 
          .D0(n21_adj_4773), .A1(d6[53]), .B1(cout_adj_5443), .C1(n132_adj_5093), 
          .D1(n20_adj_4774), .CIN(n15827), .COUT(n15828), .S0(d7_71__N_1531[52]), 
          .S1(d7_71__N_1531[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_17 (.A0(d6[50]), .B0(cout_adj_5443), .C0(n141_adj_5096), 
          .D0(n23_adj_4771), .A1(d6[51]), .B1(cout_adj_5443), .C1(n138_adj_5095), 
          .D1(n22_adj_4772), .CIN(n15826), .COUT(n15827), .S0(d7_71__N_1531[50]), 
          .S1(d7_71__N_1531[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_15 (.A0(d6[48]), .B0(cout_adj_5443), .C0(n147_adj_5098), 
          .D0(n25_adj_4769), .A1(d6[49]), .B1(cout_adj_5443), .C1(n144_adj_5097), 
          .D1(n24_adj_4770), .CIN(n15825), .COUT(n15826), .S0(d7_71__N_1531[48]), 
          .S1(d7_71__N_1531[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_13 (.A0(d6[46]), .B0(cout_adj_5443), .C0(n153_adj_5100), 
          .D0(n27_adj_4767), .A1(d6[47]), .B1(cout_adj_5443), .C1(n150_adj_5099), 
          .D1(n26_adj_4768), .CIN(n15824), .COUT(n15825), .S0(d7_71__N_1531[46]), 
          .S1(d7_71__N_1531[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_11 (.A0(d6[44]), .B0(cout_adj_5443), .C0(n159_adj_5102), 
          .D0(n29_adj_4765), .A1(d6[45]), .B1(cout_adj_5443), .C1(n156_adj_5101), 
          .D1(n28_adj_4766), .CIN(n15823), .COUT(n15824), .S0(d7_71__N_1531[44]), 
          .S1(d7_71__N_1531[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_9 (.A0(d6[42]), .B0(cout_adj_5443), .C0(n165_adj_5104), 
          .D0(n31_adj_4763), .A1(d6[43]), .B1(cout_adj_5443), .C1(n162_adj_5103), 
          .D1(n30_adj_4764), .CIN(n15822), .COUT(n15823), .S0(d7_71__N_1531[42]), 
          .S1(d7_71__N_1531[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_7 (.A0(d6[40]), .B0(cout_adj_5443), .C0(n171_adj_5106), 
          .D0(n33_adj_4761), .A1(d6[41]), .B1(cout_adj_5443), .C1(n168_adj_5105), 
          .D1(n32_adj_4762), .CIN(n15821), .COUT(n15822), .S0(d7_71__N_1531[40]), 
          .S1(d7_71__N_1531[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_5 (.A0(d6[38]), .B0(cout_adj_5443), .C0(n177_adj_5108), 
          .D0(n35_adj_4759), .A1(d6[39]), .B1(cout_adj_5443), .C1(n174_adj_5107), 
          .D1(n34_adj_4760), .CIN(n15820), .COUT(n15821), .S0(d7_71__N_1531[38]), 
          .S1(d7_71__N_1531[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_3 (.A0(d6[36]), .B0(cout_adj_5443), .C0(n183_adj_5110), 
          .D0(n37_adj_4757), .A1(d6[37]), .B1(cout_adj_5443), .C1(n180_adj_5109), 
          .D1(n36_adj_4758), .CIN(n15819), .COUT(n15820), .S0(d7_71__N_1531[36]), 
          .S1(d7_71__N_1531[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1462_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1462_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1462_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5443), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15819));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1462_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1462_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1462_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1462_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1459_add_4_13 (.A0(LOCosine[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15815), .S0(MixerOutCos_11__N_250[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1459_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_1459_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_1459_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1459_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1459_add_4_11 (.A0(LOCosine[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15814), .COUT(n15815), .S0(MixerOutCos_11__N_250[9]), 
          .S1(MixerOutCos_11__N_250[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1459_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_1459_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_1459_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1459_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1459_add_4_9 (.A0(LOCosine[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15813), .COUT(n15814), .S0(MixerOutCos_11__N_250[7]), 
          .S1(MixerOutCos_11__N_250[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1459_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_1459_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_1459_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1459_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1459_add_4_7 (.A0(LOCosine[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15812), .COUT(n15813), .S0(MixerOutCos_11__N_250[5]), 
          .S1(MixerOutCos_11__N_250[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1459_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_1459_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_1459_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1459_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1459_add_4_5 (.A0(LOCosine[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15811), .COUT(n15812), .S0(MixerOutCos_11__N_250[3]), 
          .S1(MixerOutCos_11__N_250[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1459_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_1459_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_1459_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1459_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1459_add_4_3 (.A0(LOCosine[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15810), .COUT(n15811), .S0(MixerOutCos_11__N_250[1]), 
          .S1(MixerOutCos_11__N_250[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1459_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_1459_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_1459_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1459_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1459_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOCosine[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15810), .S1(MixerOutCos_11__N_250[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(49[22:29])
    defparam _add_1_1459_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1459_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_1459_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1459_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_61 (.A0(phase_inc_carrGen[63]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15809), .S0(n124));
    defparam _add_1_1456_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_61.INIT1 = 16'h0000;
    defparam _add_1_1456_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_61.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_59 (.A0(phase_inc_carrGen[61]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[62]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15808), .COUT(n15809), .S0(n130_adj_5631), 
          .S1(n127));
    defparam _add_1_1456_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_57 (.A0(phase_inc_carrGen[59]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[60]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15807), .COUT(n15808), .S0(n136_adj_5633), 
          .S1(n133_adj_5632));
    defparam _add_1_1456_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_55 (.A0(phase_inc_carrGen[57]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[58]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15806), .COUT(n15807), .S0(n142_adj_5635), 
          .S1(n139_adj_5634));
    defparam _add_1_1456_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_53 (.A0(phase_inc_carrGen[55]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[56]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15805), .COUT(n15806), .S0(n148_adj_5637), 
          .S1(n145_adj_5636));
    defparam _add_1_1456_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_51 (.A0(phase_inc_carrGen[53]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[54]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15804), .COUT(n15805), .S0(n154_adj_5639), 
          .S1(n151_adj_5638));
    defparam _add_1_1456_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_49 (.A0(phase_inc_carrGen[51]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[52]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15803), .COUT(n15804), .S0(n160_adj_5641), 
          .S1(n157_adj_5640));
    defparam _add_1_1456_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_47 (.A0(phase_inc_carrGen[49]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[50]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15802), .COUT(n15803), .S0(n166_adj_5643), 
          .S1(n163_adj_5642));
    defparam _add_1_1456_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_1456_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_45 (.A0(phase_inc_carrGen[47]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[48]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15801), .COUT(n15802), .S0(n172_adj_5645), 
          .S1(n169_adj_5644));
    defparam _add_1_1456_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_45.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_43 (.A0(phase_inc_carrGen[45]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[46]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15800), .COUT(n15801), .S0(n178_adj_5647), 
          .S1(n175_adj_5646));
    defparam _add_1_1456_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_43.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_41 (.A0(phase_inc_carrGen[43]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[44]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15799), .COUT(n15800), .S0(n184_adj_5649), 
          .S1(n181_adj_5648));
    defparam _add_1_1456_add_4_41.INIT0 = 16'haaa0;
    defparam _add_1_1456_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_39 (.A0(phase_inc_carrGen[41]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[42]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15798), .COUT(n15799), .S0(n190_adj_5651), 
          .S1(n187_adj_5650));
    defparam _add_1_1456_add_4_39.INIT0 = 16'haaa0;
    defparam _add_1_1456_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_37 (.A0(phase_inc_carrGen[39]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[40]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15797), .COUT(n15798), .S0(n196_adj_5653), 
          .S1(n193_adj_5652));
    defparam _add_1_1456_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_35 (.A0(phase_inc_carrGen[37]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[38]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15796), .COUT(n15797), .S0(n202_adj_5655), 
          .S1(n199_adj_5654));
    defparam _add_1_1456_add_4_35.INIT0 = 16'haaa0;
    defparam _add_1_1456_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_33 (.A0(phase_inc_carrGen[35]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[36]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15795), .COUT(n15796), .S0(n208_adj_5657), 
          .S1(n205_adj_5656));
    defparam _add_1_1456_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_31 (.A0(phase_inc_carrGen[33]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[34]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15794), .COUT(n15795), .S0(n214_adj_5659), 
          .S1(n211_adj_5658));
    defparam _add_1_1456_add_4_31.INIT0 = 16'haaa0;
    defparam _add_1_1456_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_29 (.A0(phase_inc_carrGen[31]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[32]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15793), .COUT(n15794), .S0(n220_adj_5661), 
          .S1(n217_adj_5660));
    defparam _add_1_1456_add_4_29.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_29.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_29.INJECT1_1 = "NO";
    LUT4 n16_bdd_4_lut_6403 (.A(n18075), .B(led_c_3), .C(led_c_0), .D(led_c_1), 
         .Z(n17900)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n16_bdd_4_lut_6403.init = 16'hd4ef;
    LUT4 i2338_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(led_c_3), .D(n199_adj_5654), 
         .Z(n12136)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2338_3_lut_4_lut.init = 16'hf404;
    LUT4 i2340_3_lut_4_lut (.A(n18075), .B(n17937), .C(n18076), .D(n196_adj_5653), 
         .Z(n12138)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2340_3_lut_4_lut.init = 16'hf404;
    CCU2C _add_1_1456_add_4_27 (.A0(phase_inc_carrGen[29]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[30]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15792), .COUT(n15793), .S0(n226_adj_5663), 
          .S1(n223_adj_5662));
    defparam _add_1_1456_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_25 (.A0(phase_inc_carrGen[27]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[28]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15791), .COUT(n15792), .S0(n232_adj_5665), 
          .S1(n229_adj_5664));
    defparam _add_1_1456_add_4_25.INIT0 = 16'haaa0;
    defparam _add_1_1456_add_4_25.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_23 (.A0(phase_inc_carrGen[25]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[26]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15790), .COUT(n15791), .S0(n238_adj_5667), 
          .S1(n235_adj_5666));
    defparam _add_1_1456_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_21 (.A0(phase_inc_carrGen[23]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[24]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15789), .COUT(n15790), .S0(n244_adj_5669), 
          .S1(n241_adj_5668));
    defparam _add_1_1456_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_19 (.A0(phase_inc_carrGen[21]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[22]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15788), .COUT(n15789), .S0(n250_adj_5671), 
          .S1(n247_adj_5670));
    defparam _add_1_1456_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_1456_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_17 (.A0(phase_inc_carrGen[19]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[20]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15787), .COUT(n15788), .S0(n256_adj_5673), 
          .S1(n253_adj_5672));
    defparam _add_1_1456_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1456_add_4_17.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_15 (.A0(phase_inc_carrGen[17]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[18]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15786), .COUT(n15787), .S0(n262_adj_5675), 
          .S1(n259_adj_5674));
    defparam _add_1_1456_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_15.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_13 (.A0(phase_inc_carrGen[15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[16]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15785), .COUT(n15786), .S0(n268_adj_5677), 
          .S1(n265_adj_5676));
    defparam _add_1_1456_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1456_add_4_13.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_11 (.A0(phase_inc_carrGen[13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15784), .COUT(n15785), .S0(n274_adj_5679), 
          .S1(n271_adj_5678));
    defparam _add_1_1456_add_4_11.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_9 (.A0(phase_inc_carrGen[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15783), .COUT(n15784), .S0(n280_adj_5681), 
          .S1(n277_adj_5680));
    defparam _add_1_1456_add_4_9.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_7 (.A0(phase_inc_carrGen[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15782), .COUT(n15783), .S0(n286_adj_5683), 
          .S1(n283_adj_5682));
    defparam _add_1_1456_add_4_7.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_5 (.A0(phase_inc_carrGen[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15781), .COUT(n15782), .S0(n292_adj_5685), 
          .S1(n289_adj_5684));
    defparam _add_1_1456_add_4_5.INIT0 = 16'h555f;
    defparam _add_1_1456_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_3 (.A0(phase_inc_carrGen[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15780), .COUT(n15781), .S0(n298_adj_5687), 
          .S1(n295_adj_5686));
    defparam _add_1_1456_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1456_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1456_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1456_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15780), .S1(n301_adj_5688));
    defparam _add_1_1456_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1456_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1456_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1456_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_37 (.A0(d_tmp[70]), .B0(cout_adj_5551), .C0(n81_adj_5481), 
          .D0(n3_adj_4817), .A1(d_tmp[71]), .B1(cout_adj_5551), .C1(n78_adj_5480), 
          .D1(n2_adj_4818), .CIN(n15778), .S0(d6_71__N_1459[70]), .S1(d6_71__N_1459[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_35 (.A0(d_tmp[68]), .B0(cout_adj_5551), .C0(n87_adj_5483), 
          .D0(n5_adj_4815), .A1(d_tmp[69]), .B1(cout_adj_5551), .C1(n84_adj_5482), 
          .D1(n4_adj_4816), .CIN(n15777), .COUT(n15778), .S0(d6_71__N_1459[68]), 
          .S1(d6_71__N_1459[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_33 (.A0(d_tmp[66]), .B0(cout_adj_5551), .C0(n93_adj_5485), 
          .D0(n7_adj_4813), .A1(d_tmp[67]), .B1(cout_adj_5551), .C1(n90_adj_5484), 
          .D1(n6_adj_4814), .CIN(n15776), .COUT(n15777), .S0(d6_71__N_1459[66]), 
          .S1(d6_71__N_1459[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_31 (.A0(d_tmp[64]), .B0(cout_adj_5551), .C0(n99_adj_5487), 
          .D0(n9_adj_4811), .A1(d_tmp[65]), .B1(cout_adj_5551), .C1(n96_adj_5486), 
          .D1(n8_adj_4812), .CIN(n15775), .COUT(n15776), .S0(d6_71__N_1459[64]), 
          .S1(d6_71__N_1459[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_29 (.A0(d_tmp[62]), .B0(cout_adj_5551), .C0(n105_adj_5489), 
          .D0(n11_adj_4809), .A1(d_tmp[63]), .B1(cout_adj_5551), .C1(n102_adj_5488), 
          .D1(n10_adj_4810), .CIN(n15774), .COUT(n15775), .S0(d6_71__N_1459[62]), 
          .S1(d6_71__N_1459[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_27 (.A0(d_tmp[60]), .B0(cout_adj_5551), .C0(n111_adj_5491), 
          .D0(n13_adj_4807), .A1(d_tmp[61]), .B1(cout_adj_5551), .C1(n108_adj_5490), 
          .D1(n12_adj_4808), .CIN(n15773), .COUT(n15774), .S0(d6_71__N_1459[60]), 
          .S1(d6_71__N_1459[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_25 (.A0(d_tmp[58]), .B0(cout_adj_5551), .C0(n117_adj_5493), 
          .D0(n15_adj_4805), .A1(d_tmp[59]), .B1(cout_adj_5551), .C1(n114_adj_5492), 
          .D1(n14_adj_4806), .CIN(n15772), .COUT(n15773), .S0(d6_71__N_1459[58]), 
          .S1(d6_71__N_1459[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_23 (.A0(d_tmp[56]), .B0(cout_adj_5551), .C0(n123_adj_5495), 
          .D0(n17_adj_4833), .A1(d_tmp[57]), .B1(cout_adj_5551), .C1(n120_adj_5494), 
          .D1(n16_adj_4834), .CIN(n15771), .COUT(n15772), .S0(d6_71__N_1459[56]), 
          .S1(d6_71__N_1459[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_21 (.A0(d_tmp[54]), .B0(cout_adj_5551), .C0(n129_adj_5497), 
          .D0(n19_adj_4852), .A1(d_tmp[55]), .B1(cout_adj_5551), .C1(n126_adj_5496), 
          .D1(n18_adj_4835), .CIN(n15770), .COUT(n15771), .S0(d6_71__N_1459[54]), 
          .S1(d6_71__N_1459[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_19 (.A0(d_tmp[52]), .B0(cout_adj_5551), .C0(n135_adj_5499), 
          .D0(n21_adj_4850), .A1(d_tmp[53]), .B1(cout_adj_5551), .C1(n132_adj_5498), 
          .D1(n20_adj_4851), .CIN(n15769), .COUT(n15770), .S0(d6_71__N_1459[52]), 
          .S1(d6_71__N_1459[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_17 (.A0(d_tmp[50]), .B0(cout_adj_5551), .C0(n141_adj_5501), 
          .D0(n23_adj_4848), .A1(d_tmp[51]), .B1(cout_adj_5551), .C1(n138_adj_5500), 
          .D1(n22_adj_4849), .CIN(n15768), .COUT(n15769), .S0(d6_71__N_1459[50]), 
          .S1(d6_71__N_1459[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_15 (.A0(d_tmp[48]), .B0(cout_adj_5551), .C0(n147_adj_5503), 
          .D0(n25_adj_4846), .A1(d_tmp[49]), .B1(cout_adj_5551), .C1(n144_adj_5502), 
          .D1(n24_adj_4847), .CIN(n15767), .COUT(n15768), .S0(d6_71__N_1459[48]), 
          .S1(d6_71__N_1459[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_13 (.A0(d_tmp[46]), .B0(cout_adj_5551), .C0(n153_adj_5505), 
          .D0(n27_adj_4844), .A1(d_tmp[47]), .B1(cout_adj_5551), .C1(n150_adj_5504), 
          .D1(n26_adj_4845), .CIN(n15766), .COUT(n15767), .S0(d6_71__N_1459[46]), 
          .S1(d6_71__N_1459[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_11 (.A0(d_tmp[44]), .B0(cout_adj_5551), .C0(n159_adj_5507), 
          .D0(n29_adj_4842), .A1(d_tmp[45]), .B1(cout_adj_5551), .C1(n156_adj_5506), 
          .D1(n28_adj_4843), .CIN(n15765), .COUT(n15766), .S0(d6_71__N_1459[44]), 
          .S1(d6_71__N_1459[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_9 (.A0(d_tmp[42]), .B0(cout_adj_5551), .C0(n165_adj_5509), 
          .D0(n31_adj_4840), .A1(d_tmp[43]), .B1(cout_adj_5551), .C1(n162_adj_5508), 
          .D1(n30_adj_4841), .CIN(n15764), .COUT(n15765), .S0(d6_71__N_1459[42]), 
          .S1(d6_71__N_1459[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_7 (.A0(d_tmp[40]), .B0(cout_adj_5551), .C0(n171_adj_5511), 
          .D0(n33_adj_4838), .A1(d_tmp[41]), .B1(cout_adj_5551), .C1(n168_adj_5510), 
          .D1(n32_adj_4839), .CIN(n15763), .COUT(n15764), .S0(d6_71__N_1459[40]), 
          .S1(d6_71__N_1459[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_5 (.A0(d_tmp[38]), .B0(cout_adj_5551), .C0(n177_adj_5513), 
          .D0(n35_adj_4836), .A1(d_tmp[39]), .B1(cout_adj_5551), .C1(n174_adj_5512), 
          .D1(n34_adj_4837), .CIN(n15762), .COUT(n15763), .S0(d6_71__N_1459[38]), 
          .S1(d6_71__N_1459[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_3 (.A0(d_tmp[36]), .B0(cout_adj_5551), .C0(n183_adj_5515), 
          .D0(n37_adj_4854), .A1(d_tmp[37]), .B1(cout_adj_5551), .C1(n180_adj_5514), 
          .D1(n36_adj_4853), .CIN(n15761), .COUT(n15762), .S0(d6_71__N_1459[36]), 
          .S1(d6_71__N_1459[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1447_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1447_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1447_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5551), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15761));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1447_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1447_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1447_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1447_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_38 (.A0(d_d8_adj_5750[35]), .B0(d8_adj_5749[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15757), .S0(d9_71__N_1675_adj_5775[35]), 
          .S1(cout_adj_5517));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1606_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_36 (.A0(d_d8_adj_5750[33]), .B0(d8_adj_5749[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[34]), .B1(d8_adj_5749[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15756), .COUT(n15757), .S0(d9_71__N_1675_adj_5775[33]), 
          .S1(d9_71__N_1675_adj_5775[34]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_34 (.A0(d_d8_adj_5750[31]), .B0(d8_adj_5749[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[32]), .B1(d8_adj_5749[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15755), .COUT(n15756), .S0(d9_71__N_1675_adj_5775[31]), 
          .S1(d9_71__N_1675_adj_5775[32]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_32 (.A0(d_d8_adj_5750[29]), .B0(d8_adj_5749[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[30]), .B1(d8_adj_5749[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15754), .COUT(n15755), .S0(d9_71__N_1675_adj_5775[29]), 
          .S1(d9_71__N_1675_adj_5775[30]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_30 (.A0(d_d8_adj_5750[27]), .B0(d8_adj_5749[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[28]), .B1(d8_adj_5749[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15753), .COUT(n15754), .S0(d9_71__N_1675_adj_5775[27]), 
          .S1(d9_71__N_1675_adj_5775[28]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_28 (.A0(d_d8_adj_5750[25]), .B0(d8_adj_5749[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[26]), .B1(d8_adj_5749[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15752), .COUT(n15753), .S0(d9_71__N_1675_adj_5775[25]), 
          .S1(d9_71__N_1675_adj_5775[26]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_26 (.A0(d_d8_adj_5750[23]), .B0(d8_adj_5749[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[24]), .B1(d8_adj_5749[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15751), .COUT(n15752), .S0(d9_71__N_1675_adj_5775[23]), 
          .S1(d9_71__N_1675_adj_5775[24]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_24 (.A0(d_d8_adj_5750[21]), .B0(d8_adj_5749[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[22]), .B1(d8_adj_5749[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15750), .COUT(n15751), .S0(d9_71__N_1675_adj_5775[21]), 
          .S1(d9_71__N_1675_adj_5775[22]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_22 (.A0(d_d8_adj_5750[19]), .B0(d8_adj_5749[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[20]), .B1(d8_adj_5749[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15749), .COUT(n15750), .S0(d9_71__N_1675_adj_5775[19]), 
          .S1(d9_71__N_1675_adj_5775[20]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_20 (.A0(d_d8_adj_5750[17]), .B0(d8_adj_5749[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[18]), .B1(d8_adj_5749[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15748), .COUT(n15749), .S0(d9_71__N_1675_adj_5775[17]), 
          .S1(d9_71__N_1675_adj_5775[18]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_18 (.A0(d_d8_adj_5750[15]), .B0(d8_adj_5749[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[16]), .B1(d8_adj_5749[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15747), .COUT(n15748), .S0(d9_71__N_1675_adj_5775[15]), 
          .S1(d9_71__N_1675_adj_5775[16]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_16 (.A0(d_d8_adj_5750[13]), .B0(d8_adj_5749[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[14]), .B1(d8_adj_5749[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15746), .COUT(n15747), .S0(d9_71__N_1675_adj_5775[13]), 
          .S1(d9_71__N_1675_adj_5775[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_14 (.A0(d_d8_adj_5750[11]), .B0(d8_adj_5749[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[12]), .B1(d8_adj_5749[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15745), .COUT(n15746), .S0(d9_71__N_1675_adj_5775[11]), 
          .S1(d9_71__N_1675_adj_5775[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_12 (.A0(d_d8_adj_5750[9]), .B0(d8_adj_5749[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[10]), .B1(d8_adj_5749[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15744), .COUT(n15745), .S0(d9_71__N_1675_adj_5775[9]), 
          .S1(d9_71__N_1675_adj_5775[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_10 (.A0(d_d8_adj_5750[7]), .B0(d8_adj_5749[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[8]), .B1(d8_adj_5749[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15743), .COUT(n15744), .S0(d9_71__N_1675_adj_5775[7]), 
          .S1(d9_71__N_1675_adj_5775[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_8 (.A0(d_d8_adj_5750[5]), .B0(d8_adj_5749[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[6]), .B1(d8_adj_5749[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15742), .COUT(n15743), .S0(d9_71__N_1675_adj_5775[5]), 
          .S1(d9_71__N_1675_adj_5775[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_6 (.A0(d_d8_adj_5750[3]), .B0(d8_adj_5749[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[4]), .B1(d8_adj_5749[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15741), .COUT(n15742), .S0(d9_71__N_1675_adj_5775[3]), 
          .S1(d9_71__N_1675_adj_5775[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_4 (.A0(d_d8_adj_5750[1]), .B0(d8_adj_5749[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[2]), .B1(d8_adj_5749[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15740), .COUT(n15741), .S0(d9_71__N_1675_adj_5775[1]), 
          .S1(d9_71__N_1675_adj_5775[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1606_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1606_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8_adj_5750[0]), .B1(d8_adj_5749[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15740), .S1(d9_71__N_1675_adj_5775[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1606_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1606_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1606_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1606_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_63 (.A0(phase_inc_carrGen[62]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[63]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15738), .S0(n133_adj_5416), 
          .S1(n130));
    defparam _add_1_1483_add_4_63.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_63.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_63.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_63.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_61 (.A0(phase_inc_carrGen[60]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[61]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15737), .COUT(n15738), .S0(n139), 
          .S1(n136_adj_5417));
    defparam _add_1_1483_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_61.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_61.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_59 (.A0(phase_inc_carrGen[58]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[59]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15736), .COUT(n15737), .S0(n145), 
          .S1(n142));
    defparam _add_1_1483_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_57 (.A0(phase_inc_carrGen[56]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[57]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15735), .COUT(n15736), .S0(n151), 
          .S1(n148));
    defparam _add_1_1483_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_55 (.A0(phase_inc_carrGen[54]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[55]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15734), .COUT(n15735), .S0(n157), 
          .S1(n154));
    defparam _add_1_1483_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_53 (.A0(phase_inc_carrGen[52]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[53]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15733), .COUT(n15734), .S0(n163), 
          .S1(n160));
    defparam _add_1_1483_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_51 (.A0(phase_inc_carrGen[50]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[51]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15732), .COUT(n15733), .S0(n169), 
          .S1(n166));
    defparam _add_1_1483_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_49 (.A0(phase_inc_carrGen[48]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[49]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15731), .COUT(n15732), .S0(n175), 
          .S1(n172));
    defparam _add_1_1483_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_47 (.A0(phase_inc_carrGen[46]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[47]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15730), .COUT(n15731), .S0(n181), 
          .S1(n178));
    defparam _add_1_1483_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_1483_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_45 (.A0(phase_inc_carrGen[44]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[45]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15729), .COUT(n15730), .S0(n187), 
          .S1(n184));
    defparam _add_1_1483_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_45.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_43 (.A0(phase_inc_carrGen[42]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[43]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15728), .COUT(n15729), .S0(n193), 
          .S1(n190));
    defparam _add_1_1483_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_43.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_41 (.A0(phase_inc_carrGen[40]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[41]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15727), .COUT(n15728), .S0(n199), 
          .S1(n196));
    defparam _add_1_1483_add_4_41.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_39 (.A0(phase_inc_carrGen[38]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[39]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15726), .COUT(n15727), .S0(n205), 
          .S1(n202));
    defparam _add_1_1483_add_4_39.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_37 (.A0(phase_inc_carrGen[36]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[37]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15725), .COUT(n15726), .S0(n211), 
          .S1(n208));
    defparam _add_1_1483_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_35 (.A0(phase_inc_carrGen[34]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[35]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15724), .COUT(n15725), .S0(n217), 
          .S1(n214));
    defparam _add_1_1483_add_4_35.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_33 (.A0(phase_inc_carrGen[32]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[33]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15723), .COUT(n15724), .S0(n223), 
          .S1(n220));
    defparam _add_1_1483_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_31 (.A0(phase_inc_carrGen[30]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[31]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15722), .COUT(n15723), .S0(n229), 
          .S1(n226));
    defparam _add_1_1483_add_4_31.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_29 (.A0(phase_inc_carrGen[28]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[29]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15721), .COUT(n15722), .S0(n235), 
          .S1(n232));
    defparam _add_1_1483_add_4_29.INIT0 = 16'haaa0;
    defparam _add_1_1483_add_4_29.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_27 (.A0(phase_inc_carrGen[26]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[27]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15720), .COUT(n15721), .S0(n241), 
          .S1(n238));
    defparam _add_1_1483_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_25 (.A0(phase_inc_carrGen[24]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[25]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15719), .COUT(n15720), .S0(n247), 
          .S1(n244));
    defparam _add_1_1483_add_4_25.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_25.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_23 (.A0(phase_inc_carrGen[22]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[23]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15718), .COUT(n15719), .S0(n253), 
          .S1(n250));
    defparam _add_1_1483_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_21 (.A0(phase_inc_carrGen[20]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[21]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15717), .COUT(n15718), .S0(n259), 
          .S1(n256));
    defparam _add_1_1483_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_19 (.A0(phase_inc_carrGen[18]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[19]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15716), .COUT(n15717), .S0(n265), 
          .S1(n262));
    defparam _add_1_1483_add_4_19.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_17 (.A0(phase_inc_carrGen[16]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[17]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15715), .COUT(n15716), .S0(n271), 
          .S1(n268));
    defparam _add_1_1483_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1483_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_15 (.A0(phase_inc_carrGen[14]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[15]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15714), .COUT(n15715), .S0(n277), 
          .S1(n274));
    defparam _add_1_1483_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_13 (.A0(phase_inc_carrGen[12]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[13]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15713), .COUT(n15714), .S0(n283), 
          .S1(n280));
    defparam _add_1_1483_add_4_13.INIT0 = 16'h555f;
    defparam _add_1_1483_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_11 (.A0(phase_inc_carrGen[10]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[11]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15712), .COUT(n15713), .S0(n289), 
          .S1(n286));
    defparam _add_1_1483_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1483_add_4_11.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_9 (.A0(phase_inc_carrGen[8]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[9]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15711), .COUT(n15712), .S0(n295), 
          .S1(n292));
    defparam _add_1_1483_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1483_add_4_9.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_7 (.A0(phase_inc_carrGen[6]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[7]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15710), .COUT(n15711), .S0(n301), 
          .S1(n298));
    defparam _add_1_1483_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1483_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_5 (.A0(phase_inc_carrGen[4]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[5]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15709), .COUT(n15710), .S0(n307), 
          .S1(n304));
    defparam _add_1_1483_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1483_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_3 (.A0(phase_inc_carrGen[2]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen[3]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15708), .COUT(n15709), .S0(n313), 
          .S1(n310));
    defparam _add_1_1483_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1483_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1483_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1483_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_carrGen[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15708), .S1(n316));
    defparam _add_1_1483_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1483_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1483_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1483_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_37 (.A0(d1[70]), .B0(cout_adj_2824), .C0(n81_adj_5445), 
          .D0(d2[70]), .A1(d1[71]), .B1(cout_adj_2824), .C1(n78_adj_5444), 
          .D1(d2[71]), .CIN(n15706), .S0(d2_71__N_490[70]), .S1(d2_71__N_490[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_35 (.A0(d1[68]), .B0(cout_adj_2824), .C0(n87_adj_5447), 
          .D0(d2[68]), .A1(d1[69]), .B1(cout_adj_2824), .C1(n84_adj_5446), 
          .D1(d2[69]), .CIN(n15705), .COUT(n15706), .S0(d2_71__N_490[68]), 
          .S1(d2_71__N_490[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_33 (.A0(d1[66]), .B0(cout_adj_2824), .C0(n93_adj_5449), 
          .D0(d2[66]), .A1(d1[67]), .B1(cout_adj_2824), .C1(n90_adj_5448), 
          .D1(d2[67]), .CIN(n15704), .COUT(n15705), .S0(d2_71__N_490[66]), 
          .S1(d2_71__N_490[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_31 (.A0(d1[64]), .B0(cout_adj_2824), .C0(n99_adj_5451), 
          .D0(d2[64]), .A1(d1[65]), .B1(cout_adj_2824), .C1(n96_adj_5450), 
          .D1(d2[65]), .CIN(n15703), .COUT(n15704), .S0(d2_71__N_490[64]), 
          .S1(d2_71__N_490[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_29 (.A0(d1[62]), .B0(cout_adj_2824), .C0(n105_adj_5453), 
          .D0(d2[62]), .A1(d1[63]), .B1(cout_adj_2824), .C1(n102_adj_5452), 
          .D1(d2[63]), .CIN(n15702), .COUT(n15703), .S0(d2_71__N_490[62]), 
          .S1(d2_71__N_490[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_27 (.A0(d1[60]), .B0(cout_adj_2824), .C0(n111_adj_5455), 
          .D0(d2[60]), .A1(d1[61]), .B1(cout_adj_2824), .C1(n108_adj_5454), 
          .D1(d2[61]), .CIN(n15701), .COUT(n15702), .S0(d2_71__N_490[60]), 
          .S1(d2_71__N_490[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_25 (.A0(d1[58]), .B0(cout_adj_2824), .C0(n117_adj_5457), 
          .D0(d2[58]), .A1(d1[59]), .B1(cout_adj_2824), .C1(n114_adj_5456), 
          .D1(d2[59]), .CIN(n15700), .COUT(n15701), .S0(d2_71__N_490[58]), 
          .S1(d2_71__N_490[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_23 (.A0(d1[56]), .B0(cout_adj_2824), .C0(n123_adj_5459), 
          .D0(d2[56]), .A1(d1[57]), .B1(cout_adj_2824), .C1(n120_adj_5458), 
          .D1(d2[57]), .CIN(n15699), .COUT(n15700), .S0(d2_71__N_490[56]), 
          .S1(d2_71__N_490[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_21 (.A0(d1[54]), .B0(cout_adj_2824), .C0(n129_adj_5461), 
          .D0(d2[54]), .A1(d1[55]), .B1(cout_adj_2824), .C1(n126_adj_5460), 
          .D1(d2[55]), .CIN(n15698), .COUT(n15699), .S0(d2_71__N_490[54]), 
          .S1(d2_71__N_490[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_19 (.A0(d1[52]), .B0(cout_adj_2824), .C0(n135_adj_5463), 
          .D0(d2[52]), .A1(d1[53]), .B1(cout_adj_2824), .C1(n132_adj_5462), 
          .D1(d2[53]), .CIN(n15697), .COUT(n15698), .S0(d2_71__N_490[52]), 
          .S1(d2_71__N_490[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_17 (.A0(d1[50]), .B0(cout_adj_2824), .C0(n141_adj_5465), 
          .D0(d2[50]), .A1(d1[51]), .B1(cout_adj_2824), .C1(n138_adj_5464), 
          .D1(d2[51]), .CIN(n15696), .COUT(n15697), .S0(d2_71__N_490[50]), 
          .S1(d2_71__N_490[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_15 (.A0(d1[48]), .B0(cout_adj_2824), .C0(n147_adj_5467), 
          .D0(d2[48]), .A1(d1[49]), .B1(cout_adj_2824), .C1(n144_adj_5466), 
          .D1(d2[49]), .CIN(n15695), .COUT(n15696), .S0(d2_71__N_490[48]), 
          .S1(d2_71__N_490[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_13 (.A0(d1[46]), .B0(cout_adj_2824), .C0(n153_adj_5469), 
          .D0(d2[46]), .A1(d1[47]), .B1(cout_adj_2824), .C1(n150_adj_5468), 
          .D1(d2[47]), .CIN(n15694), .COUT(n15695), .S0(d2_71__N_490[46]), 
          .S1(d2_71__N_490[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_11 (.A0(d1[44]), .B0(cout_adj_2824), .C0(n159_adj_5471), 
          .D0(d2[44]), .A1(d1[45]), .B1(cout_adj_2824), .C1(n156_adj_5470), 
          .D1(d2[45]), .CIN(n15693), .COUT(n15694), .S0(d2_71__N_490[44]), 
          .S1(d2_71__N_490[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_9 (.A0(d1[42]), .B0(cout_adj_2824), .C0(n165_adj_5473), 
          .D0(d2[42]), .A1(d1[43]), .B1(cout_adj_2824), .C1(n162_adj_5472), 
          .D1(d2[43]), .CIN(n15692), .COUT(n15693), .S0(d2_71__N_490[42]), 
          .S1(d2_71__N_490[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_7 (.A0(d1[40]), .B0(cout_adj_2824), .C0(n171_adj_5475), 
          .D0(d2[40]), .A1(d1[41]), .B1(cout_adj_2824), .C1(n168_adj_5474), 
          .D1(d2[41]), .CIN(n15691), .COUT(n15692), .S0(d2_71__N_490[40]), 
          .S1(d2_71__N_490[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_5 (.A0(d1[38]), .B0(cout_adj_2824), .C0(n177_adj_5477), 
          .D0(d2[38]), .A1(d1[39]), .B1(cout_adj_2824), .C1(n174_adj_5476), 
          .D1(d2[39]), .CIN(n15690), .COUT(n15691), .S0(d2_71__N_490[38]), 
          .S1(d2_71__N_490[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_3 (.A0(d1[36]), .B0(cout_adj_2824), .C0(n183_adj_5479), 
          .D0(d2[36]), .A1(d1[37]), .B1(cout_adj_2824), .C1(n180_adj_5478), 
          .D1(d2[37]), .CIN(n15689), .COUT(n15690), .S0(d2_71__N_490[36]), 
          .S1(d2_71__N_490[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1516_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1516_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1516_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_2824), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15689));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1516_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1516_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1516_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1516_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_38 (.A0(d1_adj_5740[71]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15685), .S0(n78_adj_2860));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1570_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_36 (.A0(d1_adj_5740[69]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[70]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15684), .COUT(n15685), .S0(n84_adj_2858), 
          .S1(n81_adj_2859));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_34 (.A0(d1_adj_5740[67]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[68]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15683), .COUT(n15684), .S0(n90_adj_2856), 
          .S1(n87_adj_2857));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_32 (.A0(d1_adj_5740[65]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[66]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15682), .COUT(n15683), .S0(n96_adj_2854), 
          .S1(n93_adj_2855));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_30 (.A0(d1_adj_5740[63]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[64]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15681), .COUT(n15682), .S0(n102_adj_2852), 
          .S1(n99_adj_2853));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_28 (.A0(d1_adj_5740[61]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[62]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15680), .COUT(n15681), .S0(n108_adj_2850), 
          .S1(n105_adj_2851));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_26 (.A0(d1_adj_5740[59]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[60]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15679), .COUT(n15680), .S0(n114_adj_2848), 
          .S1(n111_adj_2849));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_24 (.A0(d1_adj_5740[57]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[58]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15678), .COUT(n15679), .S0(n120_adj_2846), 
          .S1(n117_adj_2847));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_22 (.A0(d1_adj_5740[55]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[56]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15677), .COUT(n15678), .S0(n126_adj_2844), 
          .S1(n123_adj_2845));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_20 (.A0(d1_adj_5740[53]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[54]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15676), .COUT(n15677), .S0(n132_adj_2842), 
          .S1(n129_adj_2843));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_18 (.A0(d1_adj_5740[51]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[52]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15675), .COUT(n15676), .S0(n138_adj_2840), 
          .S1(n135_adj_2841));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_16 (.A0(d1_adj_5740[49]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[50]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15674), .COUT(n15675), .S0(n144_adj_2838), 
          .S1(n141_adj_2839));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_14 (.A0(d1_adj_5740[47]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[48]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15673), .COUT(n15674), .S0(n150_adj_2836), 
          .S1(n147_adj_2837));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_12 (.A0(d1_adj_5740[45]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[46]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15672), .COUT(n15673), .S0(n156_adj_2834), 
          .S1(n153_adj_2835));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_10 (.A0(d1_adj_5740[43]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[44]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15671), .COUT(n15672), .S0(n162_adj_2832), 
          .S1(n159_adj_2833));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_8 (.A0(d1_adj_5740[41]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[42]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15670), .COUT(n15671), .S0(n168_adj_2830), 
          .S1(n165_adj_2831));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_6 (.A0(d1_adj_5740[39]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[40]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15669), .COUT(n15670), .S0(n174_adj_2828), 
          .S1(n171_adj_2829));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_4 (.A0(d1_adj_5740[37]), .B0(MixerOutCos[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d1_adj_5740[38]), .B1(MixerOutCos[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15668), .COUT(n15669), .S0(n180_adj_2826), 
          .S1(n177_adj_2827));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1570_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1570_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d1_adj_5740[36]), .B1(MixerOutCos[11]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15668), .S1(n183_adj_2825));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1570_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1570_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1570_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1570_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_37 (.A0(d4[70]), .B0(cout_adj_5326), .C0(n81_adj_5365), 
          .D0(d5[70]), .A1(d4[71]), .B1(cout_adj_5326), .C1(n78_adj_5364), 
          .D1(d5[71]), .CIN(n15666), .S0(d5_71__N_706[70]), .S1(d5_71__N_706[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_35 (.A0(d4[68]), .B0(cout_adj_5326), .C0(n87_adj_5367), 
          .D0(d5[68]), .A1(d4[69]), .B1(cout_adj_5326), .C1(n84_adj_5366), 
          .D1(d5[69]), .CIN(n15665), .COUT(n15666), .S0(d5_71__N_706[68]), 
          .S1(d5_71__N_706[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_33 (.A0(d4[66]), .B0(cout_adj_5326), .C0(n93_adj_5369), 
          .D0(d5[66]), .A1(d4[67]), .B1(cout_adj_5326), .C1(n90_adj_5368), 
          .D1(d5[67]), .CIN(n15664), .COUT(n15665), .S0(d5_71__N_706[66]), 
          .S1(d5_71__N_706[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_31 (.A0(d4[64]), .B0(cout_adj_5326), .C0(n99_adj_5371), 
          .D0(d5[64]), .A1(d4[65]), .B1(cout_adj_5326), .C1(n96_adj_5370), 
          .D1(d5[65]), .CIN(n15663), .COUT(n15664), .S0(d5_71__N_706[64]), 
          .S1(d5_71__N_706[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_29 (.A0(d4[62]), .B0(cout_adj_5326), .C0(n105_adj_5373), 
          .D0(d5[62]), .A1(d4[63]), .B1(cout_adj_5326), .C1(n102_adj_5372), 
          .D1(d5[63]), .CIN(n15662), .COUT(n15663), .S0(d5_71__N_706[62]), 
          .S1(d5_71__N_706[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_27 (.A0(d4[60]), .B0(cout_adj_5326), .C0(n111_adj_5375), 
          .D0(d5[60]), .A1(d4[61]), .B1(cout_adj_5326), .C1(n108_adj_5374), 
          .D1(d5[61]), .CIN(n15661), .COUT(n15662), .S0(d5_71__N_706[60]), 
          .S1(d5_71__N_706[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_25 (.A0(d4[58]), .B0(cout_adj_5326), .C0(n117_adj_5377), 
          .D0(d5[58]), .A1(d4[59]), .B1(cout_adj_5326), .C1(n114_adj_5376), 
          .D1(d5[59]), .CIN(n15660), .COUT(n15661), .S0(d5_71__N_706[58]), 
          .S1(d5_71__N_706[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_23 (.A0(d4[56]), .B0(cout_adj_5326), .C0(n123_adj_5379), 
          .D0(d5[56]), .A1(d4[57]), .B1(cout_adj_5326), .C1(n120_adj_5378), 
          .D1(d5[57]), .CIN(n15659), .COUT(n15660), .S0(d5_71__N_706[56]), 
          .S1(d5_71__N_706[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_21 (.A0(d4[54]), .B0(cout_adj_5326), .C0(n129_adj_5381), 
          .D0(d5[54]), .A1(d4[55]), .B1(cout_adj_5326), .C1(n126_adj_5380), 
          .D1(d5[55]), .CIN(n15658), .COUT(n15659), .S0(d5_71__N_706[54]), 
          .S1(d5_71__N_706[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_19 (.A0(d4[52]), .B0(cout_adj_5326), .C0(n135_adj_5383), 
          .D0(d5[52]), .A1(d4[53]), .B1(cout_adj_5326), .C1(n132_adj_5382), 
          .D1(d5[53]), .CIN(n15657), .COUT(n15658), .S0(d5_71__N_706[52]), 
          .S1(d5_71__N_706[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_17 (.A0(d4[50]), .B0(cout_adj_5326), .C0(n141_adj_5385), 
          .D0(d5[50]), .A1(d4[51]), .B1(cout_adj_5326), .C1(n138_adj_5384), 
          .D1(d5[51]), .CIN(n15656), .COUT(n15657), .S0(d5_71__N_706[50]), 
          .S1(d5_71__N_706[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_15 (.A0(d4[48]), .B0(cout_adj_5326), .C0(n147_adj_5387), 
          .D0(d5[48]), .A1(d4[49]), .B1(cout_adj_5326), .C1(n144_adj_5386), 
          .D1(d5[49]), .CIN(n15655), .COUT(n15656), .S0(d5_71__N_706[48]), 
          .S1(d5_71__N_706[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_13 (.A0(d4[46]), .B0(cout_adj_5326), .C0(n153_adj_5389), 
          .D0(d5[46]), .A1(d4[47]), .B1(cout_adj_5326), .C1(n150_adj_5388), 
          .D1(d5[47]), .CIN(n15654), .COUT(n15655), .S0(d5_71__N_706[46]), 
          .S1(d5_71__N_706[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_36 (.A0(d_d8_adj_5750[69]), .B0(d8_adj_5749[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[70]), .B1(d8_adj_5749[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16007), .COUT(n16008), .S0(n84_adj_4990), 
          .S1(n81_adj_4989));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_34 (.A0(d_d8_adj_5750[67]), .B0(d8_adj_5749[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[68]), .B1(d8_adj_5749[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16006), .COUT(n16007), .S0(n90_adj_4992), 
          .S1(n87_adj_4991));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_32 (.A0(d_d8_adj_5750[65]), .B0(d8_adj_5749[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[66]), .B1(d8_adj_5749[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16005), .COUT(n16006), .S0(n96_adj_4994), 
          .S1(n93_adj_4993));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_30 (.A0(d_d8_adj_5750[63]), .B0(d8_adj_5749[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[64]), .B1(d8_adj_5749[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16004), .COUT(n16005), .S0(n102_adj_4996), 
          .S1(n99_adj_4995));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_28 (.A0(d_d8_adj_5750[61]), .B0(d8_adj_5749[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[62]), .B1(d8_adj_5749[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16003), .COUT(n16004), .S0(n108_adj_4998), 
          .S1(n105_adj_4997));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_26 (.A0(d_d8_adj_5750[59]), .B0(d8_adj_5749[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[60]), .B1(d8_adj_5749[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16002), .COUT(n16003), .S0(n114_adj_5000), 
          .S1(n111_adj_4999));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_24 (.A0(d_d8_adj_5750[57]), .B0(d8_adj_5749[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[58]), .B1(d8_adj_5749[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16001), .COUT(n16002), .S0(n120_adj_5002), 
          .S1(n117_adj_5001));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_22 (.A0(d_d8_adj_5750[55]), .B0(d8_adj_5749[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[56]), .B1(d8_adj_5749[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16000), .COUT(n16001), .S0(n126_adj_5004), 
          .S1(n123_adj_5003));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_20 (.A0(d_d8_adj_5750[53]), .B0(d8_adj_5749[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[54]), .B1(d8_adj_5749[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15999), .COUT(n16000), .S0(n132_adj_5006), 
          .S1(n129_adj_5005));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_18 (.A0(d_d8_adj_5750[51]), .B0(d8_adj_5749[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[52]), .B1(d8_adj_5749[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15998), .COUT(n15999), .S0(n138_adj_5008), 
          .S1(n135_adj_5007));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_16 (.A0(d_d8_adj_5750[49]), .B0(d8_adj_5749[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[50]), .B1(d8_adj_5749[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15997), .COUT(n15998), .S0(n144_adj_5010), 
          .S1(n141_adj_5009));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_14 (.A0(d_d8_adj_5750[47]), .B0(d8_adj_5749[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[48]), .B1(d8_adj_5749[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15996), .COUT(n15997), .S0(n150_adj_5012), 
          .S1(n147_adj_5011));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_12 (.A0(d_d8_adj_5750[45]), .B0(d8_adj_5749[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[46]), .B1(d8_adj_5749[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15995), .COUT(n15996), .S0(n156_adj_5014), 
          .S1(n153_adj_5013));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_10 (.A0(d_d8_adj_5750[43]), .B0(d8_adj_5749[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[44]), .B1(d8_adj_5749[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15994), .COUT(n15995), .S0(n162_adj_5016), 
          .S1(n159_adj_5015));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_8 (.A0(d_d8_adj_5750[41]), .B0(d8_adj_5749[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[42]), .B1(d8_adj_5749[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15993), .COUT(n15994), .S0(n168_adj_5018), 
          .S1(n165_adj_5017));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_6 (.A0(d_d8_adj_5750[39]), .B0(d8_adj_5749[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[40]), .B1(d8_adj_5749[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15992), .COUT(n15993), .S0(n174_adj_5020), 
          .S1(n171_adj_5019));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_4 (.A0(d_d8_adj_5750[37]), .B0(d8_adj_5749[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d8_adj_5750[38]), .B1(d8_adj_5749[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15991), .COUT(n15992), .S0(n180_adj_5022), 
          .S1(n177_adj_5021));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1639_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1639_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8_adj_5750[36]), .B1(d8_adj_5749[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15991), .S1(n183_adj_5023));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1639_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1639_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1639_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1639_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_38 (.A0(d_d9_adj_5752[71]), .B0(d9_adj_5751[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15990), .S0(n78_adj_5024));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1642_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_36 (.A0(d_d9_adj_5752[69]), .B0(d9_adj_5751[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[70]), .B1(d9_adj_5751[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15989), .COUT(n15990), .S0(n84_adj_5026), 
          .S1(n81_adj_5025));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_34 (.A0(d_d9_adj_5752[67]), .B0(d9_adj_5751[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[68]), .B1(d9_adj_5751[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15988), .COUT(n15989), .S0(n90_adj_5028), 
          .S1(n87_adj_5027));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_32 (.A0(d_d9_adj_5752[65]), .B0(d9_adj_5751[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[66]), .B1(d9_adj_5751[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15987), .COUT(n15988), .S0(n96_adj_5030), 
          .S1(n93_adj_5029));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_30 (.A0(d_d9_adj_5752[63]), .B0(d9_adj_5751[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[64]), .B1(d9_adj_5751[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15986), .COUT(n15987), .S0(n102_adj_5032), 
          .S1(n99_adj_5031));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_28 (.A0(d_d9_adj_5752[61]), .B0(d9_adj_5751[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[62]), .B1(d9_adj_5751[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15985), .COUT(n15986), .S0(n108_adj_5034), 
          .S1(n105_adj_5033));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_26 (.A0(d_d9_adj_5752[59]), .B0(d9_adj_5751[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[60]), .B1(d9_adj_5751[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15984), .COUT(n15985), .S0(n114_adj_5036), 
          .S1(n111_adj_5035));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_24 (.A0(d_d9_adj_5752[57]), .B0(d9_adj_5751[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[58]), .B1(d9_adj_5751[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15983), .COUT(n15984), .S0(n120_adj_5038), 
          .S1(n117_adj_5037));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_22 (.A0(d_d9_adj_5752[55]), .B0(d9_adj_5751[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[56]), .B1(d9_adj_5751[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15982), .COUT(n15983));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_20 (.A0(d_d9_adj_5752[53]), .B0(d9_adj_5751[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[54]), .B1(d9_adj_5751[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15981), .COUT(n15982));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_18 (.A0(d_d9_adj_5752[51]), .B0(d9_adj_5751[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[52]), .B1(d9_adj_5751[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15980), .COUT(n15981));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_16 (.A0(d_d9_adj_5752[49]), .B0(d9_adj_5751[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[50]), .B1(d9_adj_5751[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15979), .COUT(n15980));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_14 (.A0(d_d9_adj_5752[47]), .B0(d9_adj_5751[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[48]), .B1(d9_adj_5751[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15978), .COUT(n15979));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_12 (.A0(d_d9_adj_5752[45]), .B0(d9_adj_5751[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[46]), .B1(d9_adj_5751[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15977), .COUT(n15978));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_10 (.A0(d_d9_adj_5752[43]), .B0(d9_adj_5751[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[44]), .B1(d9_adj_5751[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15976), .COUT(n15977));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_8 (.A0(d_d9_adj_5752[41]), .B0(d9_adj_5751[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[42]), .B1(d9_adj_5751[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15975), .COUT(n15976));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_6 (.A0(d_d9_adj_5752[39]), .B0(d9_adj_5751[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[40]), .B1(d9_adj_5751[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15974), .COUT(n15975));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_4 (.A0(d_d9_adj_5752[37]), .B0(d9_adj_5751[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[38]), .B1(d9_adj_5751[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15973), .COUT(n15974));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1642_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1642_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9_adj_5752[36]), .B1(d9_adj_5751[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15973));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1642_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1642_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1642_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1642_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_38 (.A0(d_d7[71]), .B0(d7[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15972), .S0(n78_adj_5039));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1645_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_36 (.A0(d_d7[69]), .B0(d7[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[70]), .B1(d7[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15971), .COUT(n15972), .S0(n84_adj_5041), .S1(n81_adj_5040));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_34 (.A0(d_d7[67]), .B0(d7[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[68]), .B1(d7[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15970), .COUT(n15971), .S0(n90_adj_5043), .S1(n87_adj_5042));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_32 (.A0(d_d7[65]), .B0(d7[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[66]), .B1(d7[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15969), .COUT(n15970), .S0(n96_adj_5045), .S1(n93_adj_5044));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_30 (.A0(d_d7[63]), .B0(d7[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[64]), .B1(d7[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15968), .COUT(n15969), .S0(n102_adj_5047), .S1(n99_adj_5046));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_28 (.A0(d_d7[61]), .B0(d7[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[62]), .B1(d7[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15967), .COUT(n15968), .S0(n108_adj_5049), .S1(n105_adj_5048));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_26 (.A0(d_d7[59]), .B0(d7[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[60]), .B1(d7[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15966), .COUT(n15967), .S0(n114_adj_5051), .S1(n111_adj_5050));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_24 (.A0(d_d7[57]), .B0(d7[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[58]), .B1(d7[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15965), .COUT(n15966), .S0(n120_adj_5053), .S1(n117_adj_5052));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_22 (.A0(d_d7[55]), .B0(d7[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[56]), .B1(d7[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15964), .COUT(n15965), .S0(n126_adj_5055), .S1(n123_adj_5054));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_20 (.A0(d_d7[53]), .B0(d7[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[54]), .B1(d7[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15963), .COUT(n15964), .S0(n132_adj_5057), .S1(n129_adj_5056));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_18 (.A0(d_d7[51]), .B0(d7[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[52]), .B1(d7[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15962), .COUT(n15963), .S0(n138_adj_5059), .S1(n135_adj_5058));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_16 (.A0(d_d7[49]), .B0(d7[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[50]), .B1(d7[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15961), .COUT(n15962), .S0(n144_adj_5061), .S1(n141_adj_5060));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_14 (.A0(d_d7[47]), .B0(d7[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[48]), .B1(d7[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15960), .COUT(n15961), .S0(n150_adj_5063), .S1(n147_adj_5062));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_12 (.A0(d_d7[45]), .B0(d7[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[46]), .B1(d7[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15959), .COUT(n15960), .S0(n156_adj_5065), .S1(n153_adj_5064));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_10 (.A0(d_d7[43]), .B0(d7[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[44]), .B1(d7[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15958), .COUT(n15959), .S0(n162_adj_5067), .S1(n159_adj_5066));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_8 (.A0(d_d7[41]), .B0(d7[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[42]), .B1(d7[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15957), .COUT(n15958), .S0(n168_adj_5069), .S1(n165_adj_5068));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_6 (.A0(d_d7[39]), .B0(d7[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[40]), .B1(d7[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15956), .COUT(n15957), .S0(n174_adj_5071), .S1(n171_adj_5070));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_4 (.A0(d_d7[37]), .B0(d7[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[38]), .B1(d7[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15955), .COUT(n15956), .S0(n180_adj_5073), .S1(n177_adj_5072));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1645_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1645_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7[36]), .B1(d7[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15955), .S1(n183_adj_5074));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1645_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1645_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1645_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1645_add_4_2.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_64 (.A0(phase_inc_carrGen1[62]), .B0(phase_accum[62]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[63]), .B1(phase_accum[63]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15953), .S0(n135_adj_4623), 
          .S1(n132_adj_4624));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_64.INIT0 = 16'h666a;
    defparam phase_accum_add_4_64.INIT1 = 16'h666a;
    defparam phase_accum_add_4_64.INJECT1_0 = "NO";
    defparam phase_accum_add_4_64.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_62 (.A0(phase_inc_carrGen1[60]), .B0(phase_accum[60]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[61]), .B1(phase_accum[61]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15952), .COUT(n15953), .S0(n141_adj_4621), 
          .S1(n138_adj_4622));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_62.INIT0 = 16'h666a;
    defparam phase_accum_add_4_62.INIT1 = 16'h666a;
    defparam phase_accum_add_4_62.INJECT1_0 = "NO";
    defparam phase_accum_add_4_62.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_60 (.A0(phase_inc_carrGen1[58]), .B0(phase_accum[58]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[59]), .B1(phase_accum[59]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15951), .COUT(n15952), .S0(n147_adj_4619), 
          .S1(n144_adj_4620));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_60.INIT0 = 16'h666a;
    defparam phase_accum_add_4_60.INIT1 = 16'h666a;
    defparam phase_accum_add_4_60.INJECT1_0 = "NO";
    defparam phase_accum_add_4_60.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_58 (.A0(phase_inc_carrGen1[56]), .B0(phase_accum[56]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[57]), .B1(phase_accum[57]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15950), .COUT(n15951), .S0(n153_adj_4617), 
          .S1(n150_adj_4618));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_58.INIT0 = 16'h666a;
    defparam phase_accum_add_4_58.INIT1 = 16'h666a;
    defparam phase_accum_add_4_58.INJECT1_0 = "NO";
    defparam phase_accum_add_4_58.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_56 (.A0(phase_inc_carrGen1[54]), .B0(phase_accum_adj_5732[54]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[55]), .B1(phase_accum_adj_5732[55]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15949), .COUT(n15950), .S0(n159_adj_4615), 
          .S1(n156_adj_4616));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_56.INIT0 = 16'h666a;
    defparam phase_accum_add_4_56.INIT1 = 16'h666a;
    defparam phase_accum_add_4_56.INJECT1_0 = "NO";
    defparam phase_accum_add_4_56.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_54 (.A0(phase_inc_carrGen1[52]), .B0(phase_accum_adj_5732[52]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[53]), .B1(phase_accum_adj_5732[53]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15948), .COUT(n15949), .S0(n165_adj_4613), 
          .S1(n162_adj_4614));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_54.INIT0 = 16'h666a;
    defparam phase_accum_add_4_54.INIT1 = 16'h666a;
    defparam phase_accum_add_4_54.INJECT1_0 = "NO";
    defparam phase_accum_add_4_54.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_52 (.A0(phase_inc_carrGen1[50]), .B0(phase_accum_adj_5732[50]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[51]), .B1(phase_accum_adj_5732[51]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15947), .COUT(n15948), .S0(n171_adj_4611), 
          .S1(n168_adj_4612));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_52.INIT0 = 16'h666a;
    defparam phase_accum_add_4_52.INIT1 = 16'h666a;
    defparam phase_accum_add_4_52.INJECT1_0 = "NO";
    defparam phase_accum_add_4_52.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_50 (.A0(phase_inc_carrGen1[48]), .B0(phase_accum_adj_5732[48]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[49]), .B1(phase_accum_adj_5732[49]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15946), .COUT(n15947), .S0(n177_adj_4609), 
          .S1(n174_adj_4610));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_50.INIT0 = 16'h666a;
    defparam phase_accum_add_4_50.INIT1 = 16'h666a;
    defparam phase_accum_add_4_50.INJECT1_0 = "NO";
    defparam phase_accum_add_4_50.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_48 (.A0(phase_inc_carrGen1[46]), .B0(phase_accum_adj_5732[46]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[47]), .B1(phase_accum_adj_5732[47]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15945), .COUT(n15946), .S0(n183_adj_4607), 
          .S1(n180_adj_4608));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_48.INIT0 = 16'h666a;
    defparam phase_accum_add_4_48.INIT1 = 16'h666a;
    defparam phase_accum_add_4_48.INJECT1_0 = "NO";
    defparam phase_accum_add_4_48.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_46 (.A0(phase_inc_carrGen1[44]), .B0(phase_accum_adj_5732[44]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[45]), .B1(phase_accum_adj_5732[45]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15944), .COUT(n15945), .S0(n189), 
          .S1(n186));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_46.INIT0 = 16'h666a;
    defparam phase_accum_add_4_46.INIT1 = 16'h666a;
    defparam phase_accum_add_4_46.INJECT1_0 = "NO";
    defparam phase_accum_add_4_46.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_44 (.A0(phase_inc_carrGen1[42]), .B0(phase_accum_adj_5732[42]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[43]), .B1(phase_accum_adj_5732[43]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15943), .COUT(n15944), .S0(n195), 
          .S1(n192));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_44.INIT0 = 16'h666a;
    defparam phase_accum_add_4_44.INIT1 = 16'h666a;
    defparam phase_accum_add_4_44.INJECT1_0 = "NO";
    defparam phase_accum_add_4_44.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_42 (.A0(phase_inc_carrGen1[40]), .B0(phase_accum_adj_5732[40]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[41]), .B1(phase_accum_adj_5732[41]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15942), .COUT(n15943), .S0(n201), 
          .S1(n198));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_42.INIT0 = 16'h666a;
    defparam phase_accum_add_4_42.INIT1 = 16'h666a;
    defparam phase_accum_add_4_42.INJECT1_0 = "NO";
    defparam phase_accum_add_4_42.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_40 (.A0(phase_inc_carrGen1[38]), .B0(phase_accum_adj_5732[38]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[39]), .B1(phase_accum_adj_5732[39]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15941), .COUT(n15942), .S0(n207), 
          .S1(n204));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_40.INIT0 = 16'h666a;
    defparam phase_accum_add_4_40.INIT1 = 16'h666a;
    defparam phase_accum_add_4_40.INJECT1_0 = "NO";
    defparam phase_accum_add_4_40.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_38 (.A0(phase_inc_carrGen1[36]), .B0(phase_accum_adj_5732[36]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[37]), .B1(phase_accum_adj_5732[37]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15940), .COUT(n15941), .S0(n213), 
          .S1(n210));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_38.INIT0 = 16'h666a;
    defparam phase_accum_add_4_38.INIT1 = 16'h666a;
    defparam phase_accum_add_4_38.INJECT1_0 = "NO";
    defparam phase_accum_add_4_38.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_36 (.A0(phase_inc_carrGen1[34]), .B0(phase_accum_adj_5732[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[35]), .B1(phase_accum_adj_5732[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15939), .COUT(n15940), .S0(n219), 
          .S1(n216));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_36.INIT0 = 16'h666a;
    defparam phase_accum_add_4_36.INIT1 = 16'h666a;
    defparam phase_accum_add_4_36.INJECT1_0 = "NO";
    defparam phase_accum_add_4_36.INJECT1_1 = "NO";
    FD1S3AX phase_accum_e3_i0_i1 (.D(n318), .CK(clk_80mhz), .Q(phase_accum_adj_5732[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i1.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i2 (.D(n315), .CK(clk_80mhz), .Q(phase_accum_adj_5732[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i2.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i3 (.D(n312), .CK(clk_80mhz), .Q(phase_accum_adj_5732[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i3.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i4 (.D(n309), .CK(clk_80mhz), .Q(phase_accum_adj_5732[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i4.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i5 (.D(n306), .CK(clk_80mhz), .Q(phase_accum_adj_5732[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i5.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i6 (.D(n303), .CK(clk_80mhz), .Q(phase_accum_adj_5732[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i6.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i7 (.D(n300), .CK(clk_80mhz), .Q(phase_accum_adj_5732[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i7.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i8 (.D(n297), .CK(clk_80mhz), .Q(phase_accum_adj_5732[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i8.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i9 (.D(n294), .CK(clk_80mhz), .Q(phase_accum_adj_5732[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i9.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i10 (.D(n291), .CK(clk_80mhz), .Q(phase_accum_adj_5732[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i10.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i11 (.D(n288), .CK(clk_80mhz), .Q(phase_accum_adj_5732[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i11.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i12 (.D(n285), .CK(clk_80mhz), .Q(phase_accum_adj_5732[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i12.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i13 (.D(n282), .CK(clk_80mhz), .Q(phase_accum_adj_5732[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i13.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i14 (.D(n279), .CK(clk_80mhz), .Q(phase_accum_adj_5732[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i14.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i15 (.D(n276), .CK(clk_80mhz), .Q(phase_accum_adj_5732[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i15.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i16 (.D(n273), .CK(clk_80mhz), .Q(phase_accum_adj_5732[16]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i16.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i17 (.D(n270), .CK(clk_80mhz), .Q(phase_accum_adj_5732[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i17.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i18 (.D(n267), .CK(clk_80mhz), .Q(phase_accum_adj_5732[18]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i18.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i19 (.D(n264), .CK(clk_80mhz), .Q(phase_accum_adj_5732[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i19.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i20 (.D(n261), .CK(clk_80mhz), .Q(phase_accum_adj_5732[20]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i20.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i21 (.D(n258), .CK(clk_80mhz), .Q(phase_accum_adj_5732[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i21.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i22 (.D(n255), .CK(clk_80mhz), .Q(phase_accum_adj_5732[22]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i22.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i23 (.D(n252), .CK(clk_80mhz), .Q(phase_accum_adj_5732[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i23.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i24 (.D(n249), .CK(clk_80mhz), .Q(phase_accum_adj_5732[24]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i24.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i25 (.D(n246), .CK(clk_80mhz), .Q(phase_accum_adj_5732[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i25.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i26 (.D(n243), .CK(clk_80mhz), .Q(phase_accum_adj_5732[26]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i26.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i27 (.D(n240), .CK(clk_80mhz), .Q(phase_accum_adj_5732[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i27.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i28 (.D(n237), .CK(clk_80mhz), .Q(phase_accum_adj_5732[28]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i28.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i29 (.D(n234), .CK(clk_80mhz), .Q(phase_accum_adj_5732[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i29.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i30 (.D(n231), .CK(clk_80mhz), .Q(phase_accum_adj_5732[30]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i30.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i31 (.D(n228), .CK(clk_80mhz), .Q(phase_accum_adj_5732[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i31.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i32 (.D(n225), .CK(clk_80mhz), .Q(phase_accum_adj_5732[32]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i32.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i33 (.D(n222), .CK(clk_80mhz), .Q(phase_accum_adj_5732[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i33.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i34 (.D(n219), .CK(clk_80mhz), .Q(phase_accum_adj_5732[34]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i34.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i35 (.D(n216), .CK(clk_80mhz), .Q(phase_accum_adj_5732[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i35.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i36 (.D(n213), .CK(clk_80mhz), .Q(phase_accum_adj_5732[36]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i36.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i37 (.D(n210), .CK(clk_80mhz), .Q(phase_accum_adj_5732[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i37.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i38 (.D(n207), .CK(clk_80mhz), .Q(phase_accum_adj_5732[38]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i38.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i39 (.D(n204), .CK(clk_80mhz), .Q(phase_accum_adj_5732[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i39.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i40 (.D(n201), .CK(clk_80mhz), .Q(phase_accum_adj_5732[40]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i40.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i41 (.D(n198), .CK(clk_80mhz), .Q(phase_accum_adj_5732[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i41.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i42 (.D(n195), .CK(clk_80mhz), .Q(phase_accum_adj_5732[42]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i42.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i43 (.D(n192), .CK(clk_80mhz), .Q(phase_accum_adj_5732[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i43.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i44 (.D(n189), .CK(clk_80mhz), .Q(phase_accum_adj_5732[44]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i44.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i45 (.D(n186), .CK(clk_80mhz), .Q(phase_accum_adj_5732[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i45.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i46 (.D(n183_adj_4607), .CK(clk_80mhz), .Q(phase_accum_adj_5732[46]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i46.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i47 (.D(n180_adj_4608), .CK(clk_80mhz), .Q(phase_accum_adj_5732[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i47.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i48 (.D(n177_adj_4609), .CK(clk_80mhz), .Q(phase_accum_adj_5732[48]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i48.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i49 (.D(n174_adj_4610), .CK(clk_80mhz), .Q(phase_accum_adj_5732[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i49.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i50 (.D(n171_adj_4611), .CK(clk_80mhz), .Q(phase_accum_adj_5732[50]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i50.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i51 (.D(n168_adj_4612), .CK(clk_80mhz), .Q(phase_accum_adj_5732[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i51.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i52 (.D(n165_adj_4613), .CK(clk_80mhz), .Q(phase_accum_adj_5732[52]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i52.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i53 (.D(n162_adj_4614), .CK(clk_80mhz), .Q(phase_accum_adj_5732[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i53.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i54 (.D(n159_adj_4615), .CK(clk_80mhz), .Q(phase_accum_adj_5732[54]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i54.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i55 (.D(n156_adj_4616), .CK(clk_80mhz), .Q(phase_accum_adj_5732[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i55.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i56 (.D(n153_adj_4617), .CK(clk_80mhz), .Q(phase_accum[56]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i56.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i57 (.D(n150_adj_4618), .CK(clk_80mhz), .Q(phase_accum[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i57.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i58 (.D(n147_adj_4619), .CK(clk_80mhz), .Q(phase_accum[58]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i58.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i59 (.D(n144_adj_4620), .CK(clk_80mhz), .Q(phase_accum[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i59.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i60 (.D(n141_adj_4621), .CK(clk_80mhz), .Q(phase_accum[60]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i60.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i61 (.D(n138_adj_4622), .CK(clk_80mhz), .Q(phase_accum[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i61.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i62 (.D(n135_adj_4623), .CK(clk_80mhz), .Q(phase_accum[62]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i62.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i63 (.D(n132_adj_4624), .CK(clk_80mhz), .Q(phase_accum[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_e3_i0_i63.GSR = "ENABLED";
    CCU2C _add_1_1507_add_4_11 (.A0(d4[44]), .B0(cout_adj_5326), .C0(n159_adj_5391), 
          .D0(d5[44]), .A1(d4[45]), .B1(cout_adj_5326), .C1(n156_adj_5390), 
          .D1(d5[45]), .CIN(n15653), .COUT(n15654), .S0(d5_71__N_706[44]), 
          .S1(d5_71__N_706[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_9 (.A0(d4[42]), .B0(cout_adj_5326), .C0(n165_adj_5393), 
          .D0(d5[42]), .A1(d4[43]), .B1(cout_adj_5326), .C1(n162_adj_5392), 
          .D1(d5[43]), .CIN(n15652), .COUT(n15653), .S0(d5_71__N_706[42]), 
          .S1(d5_71__N_706[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_7 (.A0(d4[40]), .B0(cout_adj_5326), .C0(n171_adj_5395), 
          .D0(d5[40]), .A1(d4[41]), .B1(cout_adj_5326), .C1(n168_adj_5394), 
          .D1(d5[41]), .CIN(n15651), .COUT(n15652), .S0(d5_71__N_706[40]), 
          .S1(d5_71__N_706[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_5 (.A0(d4[38]), .B0(cout_adj_5326), .C0(n177_adj_5397), 
          .D0(d5[38]), .A1(d4[39]), .B1(cout_adj_5326), .C1(n174_adj_5396), 
          .D1(d5[39]), .CIN(n15650), .COUT(n15651), .S0(d5_71__N_706[38]), 
          .S1(d5_71__N_706[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_3 (.A0(d4[36]), .B0(cout_adj_5326), .C0(n183_adj_5399), 
          .D0(d5[36]), .A1(d4[37]), .B1(cout_adj_5326), .C1(n180_adj_5398), 
          .D1(d5[37]), .CIN(n15649), .COUT(n15650), .S0(d5_71__N_706[36]), 
          .S1(d5_71__N_706[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1507_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1507_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1507_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5326), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15649));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1507_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1507_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1507_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1507_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_37 (.A0(d_d9[71]), .B0(d9[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15645), .S0(n76));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_37.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_37.INIT1 = 16'h0000;
    defparam _add_1_1486_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_35 (.A0(d_d9[69]), .B0(d9[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[70]), .B1(d9[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15644), .COUT(n15645), .S0(n82), .S1(n79));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_35.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_35.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_33 (.A0(d_d9[67]), .B0(d9[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[68]), .B1(d9[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15643), .COUT(n15644), .S0(n88), .S1(n85));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_33.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_33.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_31 (.A0(d_d9[65]), .B0(d9[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[66]), .B1(d9[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15642), .COUT(n15643), .S0(n94), .S1(n91));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_31.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_31.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_29 (.A0(d_d9[63]), .B0(d9[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[64]), .B1(d9[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15641), .COUT(n15642), .S0(n100), .S1(n97));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_29.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_29.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_27 (.A0(d_d9[61]), .B0(d9[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[62]), .B1(d9[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15640), .COUT(n15641), .S0(n106), .S1(n103));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_27.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_27.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_25 (.A0(d_d9[59]), .B0(d9[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[60]), .B1(d9[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15639), .COUT(n15640), .S0(n112), .S1(n109));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_25.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_25.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_23 (.A0(d_d9[57]), .B0(d9[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[58]), .B1(d9[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15638), .COUT(n15639), .S0(n118), .S1(n115));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_23.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_23.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_21 (.A0(d_d9[55]), .B0(d9[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[56]), .B1(d9[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15637), .COUT(n15638));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_21.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_21.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_19 (.A0(d_d9[53]), .B0(d9[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[54]), .B1(d9[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15636), .COUT(n15637));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_19.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_19.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_17 (.A0(d_d9[51]), .B0(d9[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[52]), .B1(d9[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15635), .COUT(n15636));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_17.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_17.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_15 (.A0(d_d9[49]), .B0(d9[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[50]), .B1(d9[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15634), .COUT(n15635));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_15.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_15.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_13 (.A0(d_d9[47]), .B0(d9[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[48]), .B1(d9[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15633), .COUT(n15634));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_13.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_13.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_11 (.A0(d_d9[45]), .B0(d9[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[46]), .B1(d9[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15632), .COUT(n15633));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_9 (.A0(d_d9[43]), .B0(d9[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[44]), .B1(d9[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15631), .COUT(n15632));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_7 (.A0(d_d9[41]), .B0(d9[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[42]), .B1(d9[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15630), .COUT(n15631));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_5 (.A0(d_d9[39]), .B0(d9[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[40]), .B1(d9[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15629), .COUT(n15630));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_3 (.A0(d_d9[37]), .B0(d9[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[38]), .B1(d9[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15628), .COUT(n15629));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_1486_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1486_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[36]), .B1(d9[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15628));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1486_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1486_add_4_1.INIT1 = 16'h9995;
    defparam _add_1_1486_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1486_add_4_1.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_26 (.A0(MultResult2[23]), .B0(MultResult1[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15627), .S0(n54_adj_5418));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_26.INIT0 = 16'h666a;
    defparam ISquare_add_4_26.INIT1 = 16'h0000;
    defparam ISquare_add_4_26.INJECT1_0 = "NO";
    defparam ISquare_add_4_26.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_24 (.A0(MultResult2[22]), .B0(MultResult1[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[23]), .B1(MultResult1[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15626), .COUT(n15627), .S0(n60_adj_5420), 
          .S1(n57_adj_5419));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_24.INIT0 = 16'h666a;
    defparam ISquare_add_4_24.INIT1 = 16'h666a;
    defparam ISquare_add_4_24.INJECT1_0 = "NO";
    defparam ISquare_add_4_24.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_22 (.A0(MultResult2[20]), .B0(MultResult1[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[21]), .B1(MultResult1[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15625), .COUT(n15626), .S0(n66_adj_5422), 
          .S1(n63_adj_5421));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_22.INIT0 = 16'h666a;
    defparam ISquare_add_4_22.INIT1 = 16'h666a;
    defparam ISquare_add_4_22.INJECT1_0 = "NO";
    defparam ISquare_add_4_22.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_20 (.A0(MultResult2[18]), .B0(MultResult1[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[19]), .B1(MultResult1[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15624), .COUT(n15625), .S0(n72_adj_5424), 
          .S1(n69_adj_5423));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_20.INIT0 = 16'h666a;
    defparam ISquare_add_4_20.INIT1 = 16'h666a;
    defparam ISquare_add_4_20.INJECT1_0 = "NO";
    defparam ISquare_add_4_20.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_18 (.A0(MultResult2[16]), .B0(MultResult1[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[17]), .B1(MultResult1[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15623), .COUT(n15624), .S0(n78_adj_5426), 
          .S1(n75_adj_5425));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_18.INIT0 = 16'h666a;
    defparam ISquare_add_4_18.INIT1 = 16'h666a;
    defparam ISquare_add_4_18.INJECT1_0 = "NO";
    defparam ISquare_add_4_18.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_16 (.A0(MultResult2[14]), .B0(MultResult1[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[15]), .B1(MultResult1[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15622), .COUT(n15623), .S0(n84_adj_5428), 
          .S1(n81_adj_5427));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_16.INIT0 = 16'h666a;
    defparam ISquare_add_4_16.INIT1 = 16'h666a;
    defparam ISquare_add_4_16.INJECT1_0 = "NO";
    defparam ISquare_add_4_16.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_14 (.A0(MultResult2[12]), .B0(MultResult1[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[13]), .B1(MultResult1[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15621), .COUT(n15622), .S0(n90_adj_5430), 
          .S1(n87_adj_5429));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_14.INIT0 = 16'h666a;
    defparam ISquare_add_4_14.INIT1 = 16'h666a;
    defparam ISquare_add_4_14.INJECT1_0 = "NO";
    defparam ISquare_add_4_14.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_12 (.A0(MultResult2[10]), .B0(MultResult1[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(MultResult2[11]), .B1(MultResult1[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15620), .COUT(n15621), .S0(n96_adj_5432), 
          .S1(n93_adj_5431));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_12.INIT0 = 16'h666a;
    defparam ISquare_add_4_12.INIT1 = 16'h666a;
    defparam ISquare_add_4_12.INJECT1_0 = "NO";
    defparam ISquare_add_4_12.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_10 (.A0(MultResult2[8]), .B0(MultResult1[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[9]), .B1(MultResult1[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15619), .COUT(n15620), .S0(n102_adj_5434), 
          .S1(n99_adj_5433));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_10.INIT0 = 16'h666a;
    defparam ISquare_add_4_10.INIT1 = 16'h666a;
    defparam ISquare_add_4_10.INJECT1_0 = "NO";
    defparam ISquare_add_4_10.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_8 (.A0(MultResult2[6]), .B0(MultResult1[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[7]), .B1(MultResult1[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15618), .COUT(n15619), .S0(n108_adj_5436), 
          .S1(n105_adj_5435));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_8.INIT0 = 16'h666a;
    defparam ISquare_add_4_8.INIT1 = 16'h666a;
    defparam ISquare_add_4_8.INJECT1_0 = "NO";
    defparam ISquare_add_4_8.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_6 (.A0(MultResult2[4]), .B0(MultResult1[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[5]), .B1(MultResult1[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15617), .COUT(n15618), .S0(n114_adj_5438), 
          .S1(n111_adj_5437));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_6.INIT0 = 16'h666a;
    defparam ISquare_add_4_6.INIT1 = 16'h666a;
    defparam ISquare_add_4_6.INJECT1_0 = "NO";
    defparam ISquare_add_4_6.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_4 (.A0(MultResult2[2]), .B0(MultResult1[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[3]), .B1(MultResult1[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15616), .COUT(n15617), .S0(n120_adj_5440), 
          .S1(n117_adj_5439));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_4.INIT0 = 16'h666a;
    defparam ISquare_add_4_4.INIT1 = 16'h666a;
    defparam ISquare_add_4_4.INJECT1_0 = "NO";
    defparam ISquare_add_4_4.INJECT1_1 = "NO";
    CCU2C ISquare_add_4_2 (.A0(MultResult2[0]), .B0(MultResult1[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(MultResult2[1]), .B1(MultResult1[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15616), .S1(n123_adj_5441));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(90[20:45])
    defparam ISquare_add_4_2.INIT0 = 16'h0008;
    defparam ISquare_add_4_2.INIT1 = 16'h666a;
    defparam ISquare_add_4_2.INJECT1_0 = "NO";
    defparam ISquare_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_37 (.A0(d8[70]), .B0(cout_adj_5113), .C0(n81_adj_5225), 
          .D0(n3_adj_4877), .A1(d8[71]), .B1(cout_adj_5113), .C1(n78_adj_5224), 
          .D1(n2_adj_4878), .CIN(n15613), .S0(d9_71__N_1675[70]), .S1(d9_71__N_1675[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_35 (.A0(d8[68]), .B0(cout_adj_5113), .C0(n87_adj_5227), 
          .D0(n5_adj_4875), .A1(d8[69]), .B1(cout_adj_5113), .C1(n84_adj_5226), 
          .D1(n4_adj_4876), .CIN(n15612), .COUT(n15613), .S0(d9_71__N_1675[68]), 
          .S1(d9_71__N_1675[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_33 (.A0(d8[66]), .B0(cout_adj_5113), .C0(n93_adj_5229), 
          .D0(n7_adj_4873), .A1(d8[67]), .B1(cout_adj_5113), .C1(n90_adj_5228), 
          .D1(n6_adj_4874), .CIN(n15611), .COUT(n15612), .S0(d9_71__N_1675[66]), 
          .S1(d9_71__N_1675[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_31 (.A0(d8[64]), .B0(cout_adj_5113), .C0(n99_adj_5231), 
          .D0(n9_adj_4871), .A1(d8[65]), .B1(cout_adj_5113), .C1(n96_adj_5230), 
          .D1(n8_adj_4872), .CIN(n15610), .COUT(n15611), .S0(d9_71__N_1675[64]), 
          .S1(d9_71__N_1675[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_29 (.A0(d8[62]), .B0(cout_adj_5113), .C0(n105_adj_5233), 
          .D0(n11_adj_4869), .A1(d8[63]), .B1(cout_adj_5113), .C1(n102_adj_5232), 
          .D1(n10_adj_4870), .CIN(n15609), .COUT(n15610), .S0(d9_71__N_1675[62]), 
          .S1(d9_71__N_1675[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_27 (.A0(d8[60]), .B0(cout_adj_5113), .C0(n111_adj_5235), 
          .D0(n13_adj_4867), .A1(d8[61]), .B1(cout_adj_5113), .C1(n108_adj_5234), 
          .D1(n12_adj_4868), .CIN(n15608), .COUT(n15609), .S0(d9_71__N_1675[60]), 
          .S1(d9_71__N_1675[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_25 (.A0(d8[58]), .B0(cout_adj_5113), .C0(n117_adj_5237), 
          .D0(n15_adj_4865), .A1(d8[59]), .B1(cout_adj_5113), .C1(n114_adj_5236), 
          .D1(n14_adj_4866), .CIN(n15607), .COUT(n15608), .S0(d9_71__N_1675[58]), 
          .S1(d9_71__N_1675[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_23 (.A0(d8[56]), .B0(cout_adj_5113), .C0(n123_adj_5239), 
          .D0(n17_adj_4863), .A1(d8[57]), .B1(cout_adj_5113), .C1(n120_adj_5238), 
          .D1(n16_adj_4864), .CIN(n15606), .COUT(n15607), .S0(d9_71__N_1675[56]), 
          .S1(d9_71__N_1675[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_21 (.A0(d8[54]), .B0(cout_adj_5113), .C0(n129_adj_5241), 
          .D0(n19_adj_4861), .A1(d8[55]), .B1(cout_adj_5113), .C1(n126_adj_5240), 
          .D1(n18_adj_4862), .CIN(n15605), .COUT(n15606), .S0(d9_71__N_1675[54]), 
          .S1(d9_71__N_1675[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_19 (.A0(d8[52]), .B0(cout_adj_5113), .C0(n135_adj_5243), 
          .D0(n21_adj_4859), .A1(d8[53]), .B1(cout_adj_5113), .C1(n132_adj_5242), 
          .D1(n20_adj_4860), .CIN(n15604), .COUT(n15605), .S0(d9_71__N_1675[52]), 
          .S1(d9_71__N_1675[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_17 (.A0(d8[50]), .B0(cout_adj_5113), .C0(n141_adj_5245), 
          .D0(n23_adj_4857), .A1(d8[51]), .B1(cout_adj_5113), .C1(n138_adj_5244), 
          .D1(n22_adj_4858), .CIN(n15603), .COUT(n15604), .S0(d9_71__N_1675[50]), 
          .S1(d9_71__N_1675[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_15 (.A0(d8[48]), .B0(cout_adj_5113), .C0(n147_adj_5247), 
          .D0(n25_adj_4831), .A1(d8[49]), .B1(cout_adj_5113), .C1(n144_adj_5246), 
          .D1(n24_adj_4832), .CIN(n15602), .COUT(n15603), .S0(d9_71__N_1675[48]), 
          .S1(d9_71__N_1675[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_13 (.A0(d8[46]), .B0(cout_adj_5113), .C0(n153_adj_5249), 
          .D0(n27_adj_4829), .A1(d8[47]), .B1(cout_adj_5113), .C1(n150_adj_5248), 
          .D1(n26_adj_4830), .CIN(n15601), .COUT(n15602), .S0(d9_71__N_1675[46]), 
          .S1(d9_71__N_1675[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_11 (.A0(d8[44]), .B0(cout_adj_5113), .C0(n159_adj_5251), 
          .D0(n29_adj_4827), .A1(d8[45]), .B1(cout_adj_5113), .C1(n156_adj_5250), 
          .D1(n28_adj_4828), .CIN(n15600), .COUT(n15601), .S0(d9_71__N_1675[44]), 
          .S1(d9_71__N_1675[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_9 (.A0(d8[42]), .B0(cout_adj_5113), .C0(n165_adj_5253), 
          .D0(n31_adj_4825), .A1(d8[43]), .B1(cout_adj_5113), .C1(n162_adj_5252), 
          .D1(n30_adj_4826), .CIN(n15599), .COUT(n15600), .S0(d9_71__N_1675[42]), 
          .S1(d9_71__N_1675[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_7 (.A0(d8[40]), .B0(cout_adj_5113), .C0(n171_adj_5255), 
          .D0(n33_adj_4823), .A1(d8[41]), .B1(cout_adj_5113), .C1(n168_adj_5254), 
          .D1(n32_adj_4824), .CIN(n15598), .COUT(n15599), .S0(d9_71__N_1675[40]), 
          .S1(d9_71__N_1675[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_5 (.A0(d8[38]), .B0(cout_adj_5113), .C0(n177_adj_5257), 
          .D0(n35_adj_4821), .A1(d8[39]), .B1(cout_adj_5113), .C1(n174_adj_5256), 
          .D1(n34_adj_4822), .CIN(n15597), .COUT(n15598), .S0(d9_71__N_1675[38]), 
          .S1(d9_71__N_1675[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_3 (.A0(d8[36]), .B0(cout_adj_5113), .C0(n183_adj_5259), 
          .D0(n37_adj_4819), .A1(d8[37]), .B1(cout_adj_5113), .C1(n180_adj_5258), 
          .D1(n36_adj_4820), .CIN(n15596), .COUT(n15597), .S0(d9_71__N_1675[36]), 
          .S1(d9_71__N_1675[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1489_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1489_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1489_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5113), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15596));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1489_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1489_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1489_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1489_add_4_1.INJECT1_1 = "NO";
    LUT4 i6351_3_lut_4_lut (.A(n17934), .B(n12563), .C(n18121), .D(led_c_3), 
         .Z(clk_80mhz_enable_1471)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam i6351_3_lut_4_lut.init = 16'h80f0;
    LUT4 i5418_4_lut_rep_226 (.A(n17401), .B(n17940), .C(n17906), .D(n17777), 
         .Z(n18121)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C))) */ ;
    defparam i5418_4_lut_rep_226.init = 16'hc0c8;
    LUT4 i1_2_lut (.A(led_c_3), .B(n18075), .Z(n17094)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut.init = 16'hbbbb;
    CCU2C _add_1_1621_add_4_38 (.A0(d_d_tmp_adj_5739[35]), .B0(d_tmp_adj_5738[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15592), .S0(d6_71__N_1459_adj_5772[35]), 
          .S1(cout_adj_5605));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1621_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_36 (.A0(d_d_tmp_adj_5739[33]), .B0(d_tmp_adj_5738[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[34]), .B1(d_tmp_adj_5738[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15591), .COUT(n15592), .S0(d6_71__N_1459_adj_5772[33]), 
          .S1(d6_71__N_1459_adj_5772[34]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_34 (.A0(d_d_tmp_adj_5739[31]), .B0(d_tmp_adj_5738[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[32]), .B1(d_tmp_adj_5738[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15590), .COUT(n15591), .S0(d6_71__N_1459_adj_5772[31]), 
          .S1(d6_71__N_1459_adj_5772[32]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_32 (.A0(d_d_tmp_adj_5739[29]), .B0(d_tmp_adj_5738[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[30]), .B1(d_tmp_adj_5738[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15589), .COUT(n15590), .S0(d6_71__N_1459_adj_5772[29]), 
          .S1(d6_71__N_1459_adj_5772[30]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_30 (.A0(d_d_tmp_adj_5739[27]), .B0(d_tmp_adj_5738[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[28]), .B1(d_tmp_adj_5738[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15588), .COUT(n15589), .S0(d6_71__N_1459_adj_5772[27]), 
          .S1(d6_71__N_1459_adj_5772[28]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_28 (.A0(d_d_tmp_adj_5739[25]), .B0(d_tmp_adj_5738[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[26]), .B1(d_tmp_adj_5738[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15587), .COUT(n15588), .S0(d6_71__N_1459_adj_5772[25]), 
          .S1(d6_71__N_1459_adj_5772[26]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_26 (.A0(d_d_tmp_adj_5739[23]), .B0(d_tmp_adj_5738[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[24]), .B1(d_tmp_adj_5738[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15586), .COUT(n15587), .S0(d6_71__N_1459_adj_5772[23]), 
          .S1(d6_71__N_1459_adj_5772[24]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_24 (.A0(d_d_tmp_adj_5739[21]), .B0(d_tmp_adj_5738[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[22]), .B1(d_tmp_adj_5738[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15585), .COUT(n15586), .S0(d6_71__N_1459_adj_5772[21]), 
          .S1(d6_71__N_1459_adj_5772[22]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_22 (.A0(d_d_tmp_adj_5739[19]), .B0(d_tmp_adj_5738[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[20]), .B1(d_tmp_adj_5738[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15584), .COUT(n15585), .S0(d6_71__N_1459_adj_5772[19]), 
          .S1(d6_71__N_1459_adj_5772[20]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_20 (.A0(d_d_tmp_adj_5739[17]), .B0(d_tmp_adj_5738[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[18]), .B1(d_tmp_adj_5738[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15583), .COUT(n15584), .S0(d6_71__N_1459_adj_5772[17]), 
          .S1(d6_71__N_1459_adj_5772[18]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_18 (.A0(d_d_tmp_adj_5739[15]), .B0(d_tmp_adj_5738[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[16]), .B1(d_tmp_adj_5738[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15582), .COUT(n15583), .S0(d6_71__N_1459_adj_5772[15]), 
          .S1(d6_71__N_1459_adj_5772[16]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_16 (.A0(d_d_tmp_adj_5739[13]), .B0(d_tmp_adj_5738[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[14]), .B1(d_tmp_adj_5738[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15581), .COUT(n15582), .S0(d6_71__N_1459_adj_5772[13]), 
          .S1(d6_71__N_1459_adj_5772[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_14 (.A0(d_d_tmp_adj_5739[11]), .B0(d_tmp_adj_5738[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[12]), .B1(d_tmp_adj_5738[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15580), .COUT(n15581), .S0(d6_71__N_1459_adj_5772[11]), 
          .S1(d6_71__N_1459_adj_5772[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_12 (.A0(d_d_tmp_adj_5739[9]), .B0(d_tmp_adj_5738[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[10]), .B1(d_tmp_adj_5738[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15579), .COUT(n15580), .S0(d6_71__N_1459_adj_5772[9]), 
          .S1(d6_71__N_1459_adj_5772[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_10 (.A0(d_d_tmp_adj_5739[7]), .B0(d_tmp_adj_5738[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[8]), .B1(d_tmp_adj_5738[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15578), .COUT(n15579), .S0(d6_71__N_1459_adj_5772[7]), 
          .S1(d6_71__N_1459_adj_5772[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_8 (.A0(d_d_tmp_adj_5739[5]), .B0(d_tmp_adj_5738[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[6]), .B1(d_tmp_adj_5738[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15577), .COUT(n15578), .S0(d6_71__N_1459_adj_5772[5]), 
          .S1(d6_71__N_1459_adj_5772[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_6 (.A0(d_d_tmp_adj_5739[3]), .B0(d_tmp_adj_5738[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[4]), .B1(d_tmp_adj_5738[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15576), .COUT(n15577), .S0(d6_71__N_1459_adj_5772[3]), 
          .S1(d6_71__N_1459_adj_5772[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_4 (.A0(d_d_tmp_adj_5739[1]), .B0(d_tmp_adj_5738[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[2]), .B1(d_tmp_adj_5738[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15575), .COUT(n15576), .S0(d6_71__N_1459_adj_5772[1]), 
          .S1(d6_71__N_1459_adj_5772[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1621_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1621_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp_adj_5739[0]), .B1(d_tmp_adj_5738[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15575), .S1(d6_71__N_1459_adj_5772[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1621_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1621_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1621_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1621_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_37 (.A0(d4_adj_5743[70]), .B0(cout_adj_5363), 
          .C0(n81_adj_5189), .D0(d5_adj_5744[70]), .A1(d4_adj_5743[71]), 
          .B1(cout_adj_5363), .C1(n78_adj_5188), .D1(d5_adj_5744[71]), 
          .CIN(n15573), .S0(d5_71__N_706_adj_5760[70]), .S1(d5_71__N_706_adj_5760[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_35 (.A0(d4_adj_5743[68]), .B0(cout_adj_5363), 
          .C0(n87_adj_5191), .D0(d5_adj_5744[68]), .A1(d4_adj_5743[69]), 
          .B1(cout_adj_5363), .C1(n84_adj_5190), .D1(d5_adj_5744[69]), 
          .CIN(n15572), .COUT(n15573), .S0(d5_71__N_706_adj_5760[68]), 
          .S1(d5_71__N_706_adj_5760[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_33 (.A0(d4_adj_5743[66]), .B0(cout_adj_5363), 
          .C0(n93_adj_5193), .D0(d5_adj_5744[66]), .A1(d4_adj_5743[67]), 
          .B1(cout_adj_5363), .C1(n90_adj_5192), .D1(d5_adj_5744[67]), 
          .CIN(n15571), .COUT(n15572), .S0(d5_71__N_706_adj_5760[66]), 
          .S1(d5_71__N_706_adj_5760[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_31 (.A0(d4_adj_5743[64]), .B0(cout_adj_5363), 
          .C0(n99_adj_5195), .D0(d5_adj_5744[64]), .A1(d4_adj_5743[65]), 
          .B1(cout_adj_5363), .C1(n96_adj_5194), .D1(d5_adj_5744[65]), 
          .CIN(n15570), .COUT(n15571), .S0(d5_71__N_706_adj_5760[64]), 
          .S1(d5_71__N_706_adj_5760[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_29 (.A0(d4_adj_5743[62]), .B0(cout_adj_5363), 
          .C0(n105_adj_5197), .D0(d5_adj_5744[62]), .A1(d4_adj_5743[63]), 
          .B1(cout_adj_5363), .C1(n102_adj_5196), .D1(d5_adj_5744[63]), 
          .CIN(n15569), .COUT(n15570), .S0(d5_71__N_706_adj_5760[62]), 
          .S1(d5_71__N_706_adj_5760[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_27 (.A0(d4_adj_5743[60]), .B0(cout_adj_5363), 
          .C0(n111_adj_5199), .D0(d5_adj_5744[60]), .A1(d4_adj_5743[61]), 
          .B1(cout_adj_5363), .C1(n108_adj_5198), .D1(d5_adj_5744[61]), 
          .CIN(n15568), .COUT(n15569), .S0(d5_71__N_706_adj_5760[60]), 
          .S1(d5_71__N_706_adj_5760[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_25 (.A0(d4_adj_5743[58]), .B0(cout_adj_5363), 
          .C0(n117_adj_5201), .D0(d5_adj_5744[58]), .A1(d4_adj_5743[59]), 
          .B1(cout_adj_5363), .C1(n114_adj_5200), .D1(d5_adj_5744[59]), 
          .CIN(n15567), .COUT(n15568), .S0(d5_71__N_706_adj_5760[58]), 
          .S1(d5_71__N_706_adj_5760[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_23 (.A0(d4_adj_5743[56]), .B0(cout_adj_5363), 
          .C0(n123_adj_5203), .D0(d5_adj_5744[56]), .A1(d4_adj_5743[57]), 
          .B1(cout_adj_5363), .C1(n120_adj_5202), .D1(d5_adj_5744[57]), 
          .CIN(n15566), .COUT(n15567), .S0(d5_71__N_706_adj_5760[56]), 
          .S1(d5_71__N_706_adj_5760[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_21 (.A0(d4_adj_5743[54]), .B0(cout_adj_5363), 
          .C0(n129_adj_5205), .D0(d5_adj_5744[54]), .A1(d4_adj_5743[55]), 
          .B1(cout_adj_5363), .C1(n126_adj_5204), .D1(d5_adj_5744[55]), 
          .CIN(n15565), .COUT(n15566), .S0(d5_71__N_706_adj_5760[54]), 
          .S1(d5_71__N_706_adj_5760[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_19 (.A0(d4_adj_5743[52]), .B0(cout_adj_5363), 
          .C0(n135_adj_5207), .D0(d5_adj_5744[52]), .A1(d4_adj_5743[53]), 
          .B1(cout_adj_5363), .C1(n132_adj_5206), .D1(d5_adj_5744[53]), 
          .CIN(n15564), .COUT(n15565), .S0(d5_71__N_706_adj_5760[52]), 
          .S1(d5_71__N_706_adj_5760[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_17 (.A0(d4_adj_5743[50]), .B0(cout_adj_5363), 
          .C0(n141_adj_5209), .D0(d5_adj_5744[50]), .A1(d4_adj_5743[51]), 
          .B1(cout_adj_5363), .C1(n138_adj_5208), .D1(d5_adj_5744[51]), 
          .CIN(n15563), .COUT(n15564), .S0(d5_71__N_706_adj_5760[50]), 
          .S1(d5_71__N_706_adj_5760[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_15 (.A0(d4_adj_5743[48]), .B0(cout_adj_5363), 
          .C0(n147_adj_5211), .D0(d5_adj_5744[48]), .A1(d4_adj_5743[49]), 
          .B1(cout_adj_5363), .C1(n144_adj_5210), .D1(d5_adj_5744[49]), 
          .CIN(n15562), .COUT(n15563), .S0(d5_71__N_706_adj_5760[48]), 
          .S1(d5_71__N_706_adj_5760[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_13 (.A0(d4_adj_5743[46]), .B0(cout_adj_5363), 
          .C0(n153_adj_5213), .D0(d5_adj_5744[46]), .A1(d4_adj_5743[47]), 
          .B1(cout_adj_5363), .C1(n150_adj_5212), .D1(d5_adj_5744[47]), 
          .CIN(n15561), .COUT(n15562), .S0(d5_71__N_706_adj_5760[46]), 
          .S1(d5_71__N_706_adj_5760[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_11 (.A0(d4_adj_5743[44]), .B0(cout_adj_5363), 
          .C0(n159_adj_5215), .D0(d5_adj_5744[44]), .A1(d4_adj_5743[45]), 
          .B1(cout_adj_5363), .C1(n156_adj_5214), .D1(d5_adj_5744[45]), 
          .CIN(n15560), .COUT(n15561), .S0(d5_71__N_706_adj_5760[44]), 
          .S1(d5_71__N_706_adj_5760[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_9 (.A0(d4_adj_5743[42]), .B0(cout_adj_5363), 
          .C0(n165_adj_5217), .D0(d5_adj_5744[42]), .A1(d4_adj_5743[43]), 
          .B1(cout_adj_5363), .C1(n162_adj_5216), .D1(d5_adj_5744[43]), 
          .CIN(n15559), .COUT(n15560), .S0(d5_71__N_706_adj_5760[42]), 
          .S1(d5_71__N_706_adj_5760[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_7 (.A0(d4_adj_5743[40]), .B0(cout_adj_5363), 
          .C0(n171_adj_5219), .D0(d5_adj_5744[40]), .A1(d4_adj_5743[41]), 
          .B1(cout_adj_5363), .C1(n168_adj_5218), .D1(d5_adj_5744[41]), 
          .CIN(n15558), .COUT(n15559), .S0(d5_71__N_706_adj_5760[40]), 
          .S1(d5_71__N_706_adj_5760[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_5 (.A0(d4_adj_5743[38]), .B0(cout_adj_5363), 
          .C0(n177_adj_5221), .D0(d5_adj_5744[38]), .A1(d4_adj_5743[39]), 
          .B1(cout_adj_5363), .C1(n174_adj_5220), .D1(d5_adj_5744[39]), 
          .CIN(n15557), .COUT(n15558), .S0(d5_71__N_706_adj_5760[38]), 
          .S1(d5_71__N_706_adj_5760[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_3 (.A0(d4_adj_5743[36]), .B0(cout_adj_5363), 
          .C0(n183_adj_5223), .D0(d5_adj_5744[36]), .A1(d4_adj_5743[37]), 
          .B1(cout_adj_5363), .C1(n180_adj_5222), .D1(d5_adj_5744[37]), 
          .CIN(n15556), .COUT(n15557), .S0(d5_71__N_706_adj_5760[36]), 
          .S1(d5_71__N_706_adj_5760[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1492_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1492_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1492_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5363), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15556));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1492_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1492_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1492_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1492_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1453_add_4_13 (.A0(LOSine[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15552), .S0(MixerOutSin_11__N_236[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1453_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_1453_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_1453_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1453_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1453_add_4_11 (.A0(LOSine[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15551), .COUT(n15552), .S0(MixerOutSin_11__N_236[9]), 
          .S1(MixerOutSin_11__N_236[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1453_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_1453_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_1453_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1453_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1453_add_4_9 (.A0(LOSine[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15550), .COUT(n15551), .S0(MixerOutSin_11__N_236[7]), 
          .S1(MixerOutSin_11__N_236[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1453_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_1453_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_1453_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1453_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1453_add_4_7 (.A0(LOSine[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15549), .COUT(n15550), .S0(MixerOutSin_11__N_236[5]), 
          .S1(MixerOutSin_11__N_236[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1453_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_1453_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_1453_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1453_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1453_add_4_5 (.A0(LOSine[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15548), .COUT(n15549), .S0(MixerOutSin_11__N_236[3]), 
          .S1(MixerOutSin_11__N_236[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1453_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_1453_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_1453_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1453_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1453_add_4_3 (.A0(LOSine[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15547), .COUT(n15548), .S0(MixerOutSin_11__N_236[1]), 
          .S1(MixerOutSin_11__N_236[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1453_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_1453_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_1453_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1453_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1453_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(LOSine[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15547), .S1(MixerOutSin_11__N_236[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(48[22:29])
    defparam _add_1_1453_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1453_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_1453_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1453_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_38 (.A0(d2_adj_5741[71]), .B0(d1_adj_5740[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15546), .S0(n78));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1573_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_36 (.A0(d2_adj_5741[69]), .B0(d1_adj_5740[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[70]), .B1(d1_adj_5740[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15545), .COUT(n15546), .S0(n84), 
          .S1(n81));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_34 (.A0(d2_adj_5741[67]), .B0(d1_adj_5740[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[68]), .B1(d1_adj_5740[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15544), .COUT(n15545), .S0(n90), 
          .S1(n87));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_32 (.A0(d2_adj_5741[65]), .B0(d1_adj_5740[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[66]), .B1(d1_adj_5740[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15543), .COUT(n15544), .S0(n96), 
          .S1(n93));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_30 (.A0(d2_adj_5741[63]), .B0(d1_adj_5740[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[64]), .B1(d1_adj_5740[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15542), .COUT(n15543), .S0(n102), 
          .S1(n99));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_28 (.A0(d2_adj_5741[61]), .B0(d1_adj_5740[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[62]), .B1(d1_adj_5740[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15541), .COUT(n15542), .S0(n108), 
          .S1(n105));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_26 (.A0(d2_adj_5741[59]), .B0(d1_adj_5740[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[60]), .B1(d1_adj_5740[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15540), .COUT(n15541), .S0(n114), 
          .S1(n111));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_24 (.A0(d2_adj_5741[57]), .B0(d1_adj_5740[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[58]), .B1(d1_adj_5740[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15539), .COUT(n15540), .S0(n120), 
          .S1(n117));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_22 (.A0(d2_adj_5741[55]), .B0(d1_adj_5740[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[56]), .B1(d1_adj_5740[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15538), .COUT(n15539), .S0(n126), 
          .S1(n123));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_20 (.A0(d2_adj_5741[53]), .B0(d1_adj_5740[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[54]), .B1(d1_adj_5740[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15537), .COUT(n15538), .S0(n132), 
          .S1(n129));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_18 (.A0(d2_adj_5741[51]), .B0(d1_adj_5740[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[52]), .B1(d1_adj_5740[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15536), .COUT(n15537), .S0(n138), 
          .S1(n135));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_16 (.A0(d2_adj_5741[49]), .B0(d1_adj_5740[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[50]), .B1(d1_adj_5740[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15535), .COUT(n15536), .S0(n144), 
          .S1(n141));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_14 (.A0(d2_adj_5741[47]), .B0(d1_adj_5740[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[48]), .B1(d1_adj_5740[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15534), .COUT(n15535), .S0(n150), 
          .S1(n147));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_12 (.A0(d2_adj_5741[45]), .B0(d1_adj_5740[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[46]), .B1(d1_adj_5740[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15533), .COUT(n15534), .S0(n156), 
          .S1(n153));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_10 (.A0(d2_adj_5741[43]), .B0(d1_adj_5740[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[44]), .B1(d1_adj_5740[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15532), .COUT(n15533), .S0(n162), 
          .S1(n159));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_8 (.A0(d2_adj_5741[41]), .B0(d1_adj_5740[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[42]), .B1(d1_adj_5740[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15531), .COUT(n15532), .S0(n168), 
          .S1(n165));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_6 (.A0(d2_adj_5741[39]), .B0(d1_adj_5740[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[40]), .B1(d1_adj_5740[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15530), .COUT(n15531), .S0(n174), 
          .S1(n171));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_4 (.A0(d2_adj_5741[37]), .B0(d1_adj_5740[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d2_adj_5741[38]), .B1(d1_adj_5740[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15529), .COUT(n15530), .S0(n180), 
          .S1(n177));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1573_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1573_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d2_adj_5741[36]), .B1(d1_adj_5740[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15529), .S1(n183));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1573_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1573_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1573_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1573_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_37 (.A0(d3[70]), .B0(cout_adj_5288), .C0(n81_adj_5690), 
          .D0(d4[70]), .A1(d3[71]), .B1(cout_adj_5288), .C1(n78_adj_5689), 
          .D1(d4[71]), .CIN(n15527), .S0(d4_71__N_634[70]), .S1(d4_71__N_634[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_35 (.A0(d3[68]), .B0(cout_adj_5288), .C0(n87_adj_5692), 
          .D0(d4[68]), .A1(d3[69]), .B1(cout_adj_5288), .C1(n84_adj_5691), 
          .D1(d4[69]), .CIN(n15526), .COUT(n15527), .S0(d4_71__N_634[68]), 
          .S1(d4_71__N_634[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_33 (.A0(d3[66]), .B0(cout_adj_5288), .C0(n93_adj_5694), 
          .D0(d4[66]), .A1(d3[67]), .B1(cout_adj_5288), .C1(n90_adj_5693), 
          .D1(d4[67]), .CIN(n15525), .COUT(n15526), .S0(d4_71__N_634[66]), 
          .S1(d4_71__N_634[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_31 (.A0(d3[64]), .B0(cout_adj_5288), .C0(n99_adj_5696), 
          .D0(d4[64]), .A1(d3[65]), .B1(cout_adj_5288), .C1(n96_adj_5695), 
          .D1(d4[65]), .CIN(n15524), .COUT(n15525), .S0(d4_71__N_634[64]), 
          .S1(d4_71__N_634[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_29 (.A0(d3[62]), .B0(cout_adj_5288), .C0(n105_adj_5698), 
          .D0(d4[62]), .A1(d3[63]), .B1(cout_adj_5288), .C1(n102_adj_5697), 
          .D1(d4[63]), .CIN(n15523), .COUT(n15524), .S0(d4_71__N_634[62]), 
          .S1(d4_71__N_634[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_27 (.A0(d3[60]), .B0(cout_adj_5288), .C0(n111_adj_5700), 
          .D0(d4[60]), .A1(d3[61]), .B1(cout_adj_5288), .C1(n108_adj_5699), 
          .D1(d4[61]), .CIN(n15522), .COUT(n15523), .S0(d4_71__N_634[60]), 
          .S1(d4_71__N_634[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_25 (.A0(d3[58]), .B0(cout_adj_5288), .C0(n117_adj_5702), 
          .D0(d4[58]), .A1(d3[59]), .B1(cout_adj_5288), .C1(n114_adj_5701), 
          .D1(d4[59]), .CIN(n15521), .COUT(n15522), .S0(d4_71__N_634[58]), 
          .S1(d4_71__N_634[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_23 (.A0(d3[56]), .B0(cout_adj_5288), .C0(n123_adj_5704), 
          .D0(d4[56]), .A1(d3[57]), .B1(cout_adj_5288), .C1(n120_adj_5703), 
          .D1(d4[57]), .CIN(n15520), .COUT(n15521), .S0(d4_71__N_634[56]), 
          .S1(d4_71__N_634[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_21 (.A0(d3[54]), .B0(cout_adj_5288), .C0(n129_adj_5706), 
          .D0(d4[54]), .A1(d3[55]), .B1(cout_adj_5288), .C1(n126_adj_5705), 
          .D1(d4[55]), .CIN(n15519), .COUT(n15520), .S0(d4_71__N_634[54]), 
          .S1(d4_71__N_634[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_19 (.A0(d3[52]), .B0(cout_adj_5288), .C0(n135_adj_5708), 
          .D0(d4[52]), .A1(d3[53]), .B1(cout_adj_5288), .C1(n132_adj_5707), 
          .D1(d4[53]), .CIN(n15518), .COUT(n15519), .S0(d4_71__N_634[52]), 
          .S1(d4_71__N_634[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_17 (.A0(d3[50]), .B0(cout_adj_5288), .C0(n141_adj_5710), 
          .D0(d4[50]), .A1(d3[51]), .B1(cout_adj_5288), .C1(n138_adj_5709), 
          .D1(d4[51]), .CIN(n15517), .COUT(n15518), .S0(d4_71__N_634[50]), 
          .S1(d4_71__N_634[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_15 (.A0(d3[48]), .B0(cout_adj_5288), .C0(n147_adj_5712), 
          .D0(d4[48]), .A1(d3[49]), .B1(cout_adj_5288), .C1(n144_adj_5711), 
          .D1(d4[49]), .CIN(n15516), .COUT(n15517), .S0(d4_71__N_634[48]), 
          .S1(d4_71__N_634[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_13 (.A0(d3[46]), .B0(cout_adj_5288), .C0(n153_adj_5714), 
          .D0(d4[46]), .A1(d3[47]), .B1(cout_adj_5288), .C1(n150_adj_5713), 
          .D1(d4[47]), .CIN(n15515), .COUT(n15516), .S0(d4_71__N_634[46]), 
          .S1(d4_71__N_634[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_11 (.A0(d3[44]), .B0(cout_adj_5288), .C0(n159_adj_5716), 
          .D0(d4[44]), .A1(d3[45]), .B1(cout_adj_5288), .C1(n156_adj_5715), 
          .D1(d4[45]), .CIN(n15514), .COUT(n15515), .S0(d4_71__N_634[44]), 
          .S1(d4_71__N_634[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_9 (.A0(d3[42]), .B0(cout_adj_5288), .C0(n165_adj_5718), 
          .D0(d4[42]), .A1(d3[43]), .B1(cout_adj_5288), .C1(n162_adj_5717), 
          .D1(d4[43]), .CIN(n15513), .COUT(n15514), .S0(d4_71__N_634[42]), 
          .S1(d4_71__N_634[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_7 (.A0(d3[40]), .B0(cout_adj_5288), .C0(n171_adj_5720), 
          .D0(d4[40]), .A1(d3[41]), .B1(cout_adj_5288), .C1(n168_adj_5719), 
          .D1(d4[41]), .CIN(n15512), .COUT(n15513), .S0(d4_71__N_634[40]), 
          .S1(d4_71__N_634[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_5 (.A0(d3[38]), .B0(cout_adj_5288), .C0(n177_adj_5722), 
          .D0(d4[38]), .A1(d3[39]), .B1(cout_adj_5288), .C1(n174_adj_5721), 
          .D1(d4[39]), .CIN(n15511), .COUT(n15512), .S0(d4_71__N_634[38]), 
          .S1(d4_71__N_634[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_3 (.A0(d3[36]), .B0(cout_adj_5288), .C0(n183_adj_5724), 
          .D0(d4[36]), .A1(d3[37]), .B1(cout_adj_5288), .C1(n180_adj_5723), 
          .D1(d4[37]), .CIN(n15510), .COUT(n15511), .S0(d4_71__N_634[36]), 
          .S1(d4_71__N_634[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1510_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1510_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1510_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5288), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15510));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1510_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1510_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1510_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1510_add_4_1.INJECT1_1 = "NO";
    CCU2C add_3837_19 (.A0(d_out_d_11__N_1882[17]), .B0(n48_adj_5347), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n45_adj_5346), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15505), .S0(n45_adj_5518), 
          .S1(d_out_d_11__N_1884[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3837_19.INIT0 = 16'h9995;
    defparam add_3837_19.INIT1 = 16'h9995;
    defparam add_3837_19.INJECT1_0 = "NO";
    defparam add_3837_19.INJECT1_1 = "NO";
    CCU2C add_3837_17 (.A0(d_out_d_11__N_1882[17]), .B0(n54_adj_5349), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n51_adj_5348), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15504), .COUT(n15505), .S0(n51_adj_5520), 
          .S1(n48_adj_5519));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3837_17.INIT0 = 16'h9995;
    defparam add_3837_17.INIT1 = 16'h9995;
    defparam add_3837_17.INJECT1_0 = "NO";
    defparam add_3837_17.INJECT1_1 = "NO";
    CCU2C add_3837_15 (.A0(d_out_d_11__N_1882[17]), .B0(n60_adj_5351), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n57_adj_5350), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15503), .COUT(n15504), .S0(n57_adj_5522), 
          .S1(n54_adj_5521));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3837_15.INIT0 = 16'h9995;
    defparam add_3837_15.INIT1 = 16'h9995;
    defparam add_3837_15.INJECT1_0 = "NO";
    defparam add_3837_15.INJECT1_1 = "NO";
    CCU2C add_3837_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1882[17]), .C0(n66_adj_5353), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1882[17]), 
          .C1(n63_adj_5352), .D1(VCC_net), .CIN(n15502), .COUT(n15503), 
          .S0(n63_adj_5524), .S1(n60_adj_5523));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3837_13.INIT0 = 16'h6969;
    defparam add_3837_13.INIT1 = 16'h6969;
    defparam add_3837_13.INJECT1_0 = "NO";
    defparam add_3837_13.INJECT1_1 = "NO";
    CCU2C add_3837_11 (.A0(d_out_d_11__N_1882[17]), .B0(n72_adj_5355), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1882[17]), 
          .C1(n69_adj_5354), .D1(VCC_net), .CIN(n15501), .COUT(n15502), 
          .S0(n69_adj_5526), .S1(n66_adj_5525));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3837_11.INIT0 = 16'h9995;
    defparam add_3837_11.INIT1 = 16'h6969;
    defparam add_3837_11.INJECT1_0 = "NO";
    defparam add_3837_11.INJECT1_1 = "NO";
    CCU2C add_3837_9 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1882[17]), 
          .C0(n78_adj_5357), .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), 
          .B1(n17938), .C1(n75_adj_5356), .D1(VCC_net), .CIN(n15500), 
          .COUT(n15501), .S0(n75_adj_5528), .S1(n72_adj_5527));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3837_9.INIT0 = 16'h9696;
    defparam add_3837_9.INIT1 = 16'h6969;
    defparam add_3837_9.INJECT1_0 = "NO";
    defparam add_3837_9.INJECT1_1 = "NO";
    CCU2C add_3837_7 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1882[17]), 
          .C0(n84_adj_5359), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1882[17]), .C1(n81_adj_5358), .D1(VCC_net), 
          .CIN(n15499), .COUT(n15500), .S0(n81_adj_5530), .S1(n78_adj_5529));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3837_7.INIT0 = 16'h9696;
    defparam add_3837_7.INIT1 = 16'h9696;
    defparam add_3837_7.INJECT1_0 = "NO";
    defparam add_3837_7.INJECT1_1 = "NO";
    CCU2C add_3837_5 (.A0(n90_adj_5361), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1880[17]), .B1(d_out_d_11__N_1882[17]), .C1(n87_adj_5360), 
          .D1(VCC_net), .CIN(n15498), .COUT(n15499), .S0(n87_adj_5532), 
          .S1(n84_adj_5531));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3837_5.INIT0 = 16'haaa0;
    defparam add_3837_5.INIT1 = 16'h9696;
    defparam add_3837_5.INJECT1_0 = "NO";
    defparam add_3837_5.INJECT1_1 = "NO";
    CCU2C add_3837_3 (.A0(d_out_d_11__N_1882[17]), .B0(ISquare[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15497), .COUT(n15498), .S1(n90_adj_5533));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3837_3.INIT0 = 16'h666a;
    defparam add_3837_3.INIT1 = 16'h555f;
    defparam add_3837_3.INJECT1_0 = "NO";
    defparam add_3837_3.INJECT1_1 = "NO";
    CCU2C add_3837_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1882[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15497));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3837_1.INIT0 = 16'h0000;
    defparam add_3837_1.INIT1 = 16'haaaf;
    defparam add_3837_1.INJECT1_0 = "NO";
    defparam add_3837_1.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_38 (.A0(d_d6[35]), .B0(d6[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15492), .S0(d7_71__N_1531[35]), .S1(cout_adj_5443));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1522_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_36 (.A0(d_d6[33]), .B0(d6[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[34]), .B1(d6[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15491), .COUT(n15492), .S0(d7_71__N_1531[33]), .S1(d7_71__N_1531[34]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_34 (.A0(d_d6[31]), .B0(d6[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[32]), .B1(d6[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15490), .COUT(n15491), .S0(d7_71__N_1531[31]), .S1(d7_71__N_1531[32]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_32 (.A0(d_d6[29]), .B0(d6[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[30]), .B1(d6[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15489), .COUT(n15490), .S0(d7_71__N_1531[29]), .S1(d7_71__N_1531[30]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_30 (.A0(d_d6[27]), .B0(d6[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[28]), .B1(d6[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15488), .COUT(n15489), .S0(d7_71__N_1531[27]), .S1(d7_71__N_1531[28]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_28 (.A0(d_d6[25]), .B0(d6[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[26]), .B1(d6[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15487), .COUT(n15488), .S0(d7_71__N_1531[25]), .S1(d7_71__N_1531[26]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_26 (.A0(d_d6[23]), .B0(d6[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[24]), .B1(d6[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15486), .COUT(n15487), .S0(d7_71__N_1531[23]), .S1(d7_71__N_1531[24]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_24 (.A0(d_d6[21]), .B0(d6[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[22]), .B1(d6[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15485), .COUT(n15486), .S0(d7_71__N_1531[21]), .S1(d7_71__N_1531[22]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_22 (.A0(d_d6[19]), .B0(d6[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[20]), .B1(d6[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15484), .COUT(n15485), .S0(d7_71__N_1531[19]), .S1(d7_71__N_1531[20]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_20 (.A0(d_d6[17]), .B0(d6[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[18]), .B1(d6[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15483), .COUT(n15484), .S0(d7_71__N_1531[17]), .S1(d7_71__N_1531[18]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_18 (.A0(d_d6[15]), .B0(d6[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[16]), .B1(d6[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15482), .COUT(n15483), .S0(d7_71__N_1531[15]), .S1(d7_71__N_1531[16]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_16 (.A0(d_d6[13]), .B0(d6[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[14]), .B1(d6[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15481), .COUT(n15482), .S0(d7_71__N_1531[13]), .S1(d7_71__N_1531[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_14 (.A0(d_d6[11]), .B0(d6[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[12]), .B1(d6[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15480), .COUT(n15481), .S0(d7_71__N_1531[11]), .S1(d7_71__N_1531[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_12 (.A0(d_d6[9]), .B0(d6[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[10]), .B1(d6[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15479), .COUT(n15480), .S0(d7_71__N_1531[9]), .S1(d7_71__N_1531[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_10 (.A0(d_d6[7]), .B0(d6[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[8]), .B1(d6[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15478), .COUT(n15479), .S0(d7_71__N_1531[7]), .S1(d7_71__N_1531[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_8 (.A0(d_d6[5]), .B0(d6[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[6]), .B1(d6[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15477), .COUT(n15478), .S0(d7_71__N_1531[5]), .S1(d7_71__N_1531[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_6 (.A0(d_d6[3]), .B0(d6[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[4]), .B1(d6[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15476), .COUT(n15477), .S0(d7_71__N_1531[3]), .S1(d7_71__N_1531[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_4 (.A0(d_d6[1]), .B0(d6[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[2]), .B1(d6[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15475), .COUT(n15476), .S0(d7_71__N_1531[1]), .S1(d7_71__N_1531[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1522_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1522_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[0]), .B1(d6[0]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15475), .S1(d7_71__N_1531[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1522_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1522_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1522_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1522_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_38 (.A0(d2[71]), .B0(d1[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15474), .S0(n78_adj_5444));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1558_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_36 (.A0(d2[69]), .B0(d1[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[70]), .B1(d1[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15473), .COUT(n15474), .S0(n84_adj_5446), .S1(n81_adj_5445));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_34 (.A0(d2[67]), .B0(d1[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[68]), .B1(d1[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15472), .COUT(n15473), .S0(n90_adj_5448), .S1(n87_adj_5447));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_32 (.A0(d2[65]), .B0(d1[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[66]), .B1(d1[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15471), .COUT(n15472), .S0(n96_adj_5450), .S1(n93_adj_5449));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_30 (.A0(d2[63]), .B0(d1[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[64]), .B1(d1[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15470), .COUT(n15471), .S0(n102_adj_5452), .S1(n99_adj_5451));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_28 (.A0(d2[61]), .B0(d1[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[62]), .B1(d1[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15469), .COUT(n15470), .S0(n108_adj_5454), .S1(n105_adj_5453));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_26 (.A0(d2[59]), .B0(d1[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[60]), .B1(d1[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15468), .COUT(n15469), .S0(n114_adj_5456), .S1(n111_adj_5455));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_24 (.A0(d2[57]), .B0(d1[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[58]), .B1(d1[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15467), .COUT(n15468), .S0(n120_adj_5458), .S1(n117_adj_5457));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_22 (.A0(d2[55]), .B0(d1[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[56]), .B1(d1[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15466), .COUT(n15467), .S0(n126_adj_5460), .S1(n123_adj_5459));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_20 (.A0(d2[53]), .B0(d1[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[54]), .B1(d1[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15465), .COUT(n15466), .S0(n132_adj_5462), .S1(n129_adj_5461));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_18 (.A0(d2[51]), .B0(d1[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[52]), .B1(d1[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15464), .COUT(n15465), .S0(n138_adj_5464), .S1(n135_adj_5463));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_16 (.A0(d2[49]), .B0(d1[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[50]), .B1(d1[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15463), .COUT(n15464), .S0(n144_adj_5466), .S1(n141_adj_5465));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_14 (.A0(d2[47]), .B0(d1[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[48]), .B1(d1[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15462), .COUT(n15463), .S0(n150_adj_5468), .S1(n147_adj_5467));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_12 (.A0(d2[45]), .B0(d1[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[46]), .B1(d1[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15461), .COUT(n15462), .S0(n156_adj_5470), .S1(n153_adj_5469));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_10 (.A0(d2[43]), .B0(d1[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[44]), .B1(d1[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15460), .COUT(n15461), .S0(n162_adj_5472), .S1(n159_adj_5471));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_8 (.A0(d2[41]), .B0(d1[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[42]), .B1(d1[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15459), .COUT(n15460), .S0(n168_adj_5474), .S1(n165_adj_5473));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_6 (.A0(d2[39]), .B0(d1[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[40]), .B1(d1[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15458), .COUT(n15459), .S0(n174_adj_5476), .S1(n171_adj_5475));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_4 (.A0(d2[37]), .B0(d1[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[38]), .B1(d1[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15457), .COUT(n15458), .S0(n180_adj_5478), .S1(n177_adj_5477));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1558_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1558_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[36]), .B1(d1[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15457), .S1(n183_adj_5479));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1558_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1558_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1558_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1558_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_38 (.A0(d_d8[71]), .B0(d8[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15456), .S0(n78_adj_5224));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1585_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_36 (.A0(d_d8[69]), .B0(d8[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[70]), .B1(d8[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15455), .COUT(n15456), .S0(n84_adj_5226), .S1(n81_adj_5225));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_34 (.A0(d_d8[67]), .B0(d8[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[68]), .B1(d8[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15454), .COUT(n15455), .S0(n90_adj_5228), .S1(n87_adj_5227));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_32 (.A0(d_d8[65]), .B0(d8[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[66]), .B1(d8[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15453), .COUT(n15454), .S0(n96_adj_5230), .S1(n93_adj_5229));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_30 (.A0(d_d8[63]), .B0(d8[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[64]), .B1(d8[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15452), .COUT(n15453), .S0(n102_adj_5232), .S1(n99_adj_5231));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_28 (.A0(d_d8[61]), .B0(d8[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[62]), .B1(d8[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15451), .COUT(n15452), .S0(n108_adj_5234), .S1(n105_adj_5233));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_26 (.A0(d_d8[59]), .B0(d8[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[60]), .B1(d8[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15450), .COUT(n15451), .S0(n114_adj_5236), .S1(n111_adj_5235));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_24 (.A0(d_d8[57]), .B0(d8[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[58]), .B1(d8[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15449), .COUT(n15450), .S0(n120_adj_5238), .S1(n117_adj_5237));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_22 (.A0(d_d8[55]), .B0(d8[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[56]), .B1(d8[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15448), .COUT(n15449), .S0(n126_adj_5240), .S1(n123_adj_5239));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_20 (.A0(d_d8[53]), .B0(d8[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[54]), .B1(d8[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15447), .COUT(n15448), .S0(n132_adj_5242), .S1(n129_adj_5241));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_18 (.A0(d_d8[51]), .B0(d8[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[52]), .B1(d8[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15446), .COUT(n15447), .S0(n138_adj_5244), .S1(n135_adj_5243));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_16 (.A0(d_d8[49]), .B0(d8[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[50]), .B1(d8[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15445), .COUT(n15446), .S0(n144_adj_5246), .S1(n141_adj_5245));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_14 (.A0(d_d8[47]), .B0(d8[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[48]), .B1(d8[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15444), .COUT(n15445), .S0(n150_adj_5248), .S1(n147_adj_5247));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_12 (.A0(d_d8[45]), .B0(d8[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[46]), .B1(d8[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15443), .COUT(n15444), .S0(n156_adj_5250), .S1(n153_adj_5249));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_10 (.A0(d_d8[43]), .B0(d8[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[44]), .B1(d8[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15442), .COUT(n15443), .S0(n162_adj_5252), .S1(n159_adj_5251));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_8 (.A0(d_d8[41]), .B0(d8[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[42]), .B1(d8[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15441), .COUT(n15442), .S0(n168_adj_5254), .S1(n165_adj_5253));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_6 (.A0(d_d8[39]), .B0(d8[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[40]), .B1(d8[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15440), .COUT(n15441), .S0(n174_adj_5256), .S1(n171_adj_5255));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_4 (.A0(d_d8[37]), .B0(d8[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[38]), .B1(d8[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15439), .COUT(n15440), .S0(n180_adj_5258), .S1(n177_adj_5257));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1585_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1585_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d8[36]), .B1(d8[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15439), .S1(n183_adj_5259));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1585_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1585_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1585_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1585_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_38 (.A0(d_d9[71]), .B0(d9[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15438), .S0(n78_adj_5260));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1588_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_36 (.A0(d_d9[69]), .B0(d9[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[70]), .B1(d9[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15437), .COUT(n15438), .S0(n84_adj_5262), .S1(n81_adj_5261));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_34 (.A0(d_d9[67]), .B0(d9[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[68]), .B1(d9[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15436), .COUT(n15437), .S0(n90_adj_5264), .S1(n87_adj_5263));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_32 (.A0(d_d9[65]), .B0(d9[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[66]), .B1(d9[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15435), .COUT(n15436), .S0(n96_adj_5266), .S1(n93_adj_5265));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_30 (.A0(d_d9[63]), .B0(d9[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[64]), .B1(d9[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15434), .COUT(n15435), .S0(n102_adj_5268), .S1(n99_adj_5267));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_28 (.A0(d_d9[61]), .B0(d9[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[62]), .B1(d9[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15433), .COUT(n15434), .S0(n108_adj_5270), .S1(n105_adj_5269));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_26 (.A0(d_d9[59]), .B0(d9[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[60]), .B1(d9[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15432), .COUT(n15433), .S0(n114_adj_5272), .S1(n111_adj_5271));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_24 (.A0(d_d9[57]), .B0(d9[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[58]), .B1(d9[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15431), .COUT(n15432), .S0(n120_adj_5274), .S1(n117_adj_5273));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_22 (.A0(d_d9[55]), .B0(d9[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[56]), .B1(d9[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15430), .COUT(n15431));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_20 (.A0(d_d9[53]), .B0(d9[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[54]), .B1(d9[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15429), .COUT(n15430));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_18 (.A0(d_d9[51]), .B0(d9[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[52]), .B1(d9[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15428), .COUT(n15429));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_16 (.A0(d_d9[49]), .B0(d9[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[50]), .B1(d9[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15427), .COUT(n15428));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_14 (.A0(d_d9[47]), .B0(d9[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[48]), .B1(d9[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15426), .COUT(n15427));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_12 (.A0(d_d9[45]), .B0(d9[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[46]), .B1(d9[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15425), .COUT(n15426));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_10 (.A0(d_d9[43]), .B0(d9[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[44]), .B1(d9[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15424), .COUT(n15425));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_8 (.A0(d_d9[41]), .B0(d9[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[42]), .B1(d9[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15423), .COUT(n15424));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_6 (.A0(d_d9[39]), .B0(d9[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[40]), .B1(d9[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15422), .COUT(n15423));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_4 (.A0(d_d9[37]), .B0(d9[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[38]), .B1(d9[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15421), .COUT(n15422));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1588_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1588_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[36]), .B1(d9[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15421));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1588_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1588_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1588_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1588_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1591_add_4_20 (.A0(n916), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15420), .S0(d_out_d_11__N_2383[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1591_add_4_20.INIT0 = 16'h555f;
    defparam _add_1_1591_add_4_20.INIT1 = 16'h0000;
    defparam _add_1_1591_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1591_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1591_add_4_18 (.A0(ISquare[31]), .B0(n918), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(n917), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15419), .COUT(n15420));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1591_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1591_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1591_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1591_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1591_add_4_16 (.A0(n920), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(n919), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15418), .COUT(n15419));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1591_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1591_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1591_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1591_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1591_add_4_14 (.A0(d_out_d_11__N_1874[17]), .B0(n922), 
          .C0(GND_net), .D0(VCC_net), .A1(ISquare[31]), .B1(n17942), 
          .C1(n921), .D1(VCC_net), .CIN(n15417), .COUT(n15418));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1591_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1591_add_4_14.INIT1 = 16'he1e1;
    defparam _add_1_1591_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1591_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1591_add_4_12 (.A0(d_out_d_11__N_1878[17]), .B0(n924), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n923), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15416), .COUT(n15417));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1591_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1591_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1591_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1591_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1591_add_4_10 (.A0(d_out_d_11__N_1882[17]), .B0(n926), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n925), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15415), .COUT(n15416));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1591_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1591_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1591_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1591_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1591_add_4_8 (.A0(d_out_d_11__N_1886[17]), .B0(n928), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), .B1(n927), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15414), .COUT(n15415));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1591_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1591_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1591_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1591_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1591_add_4_6 (.A0(d_out_d_11__N_1890[17]), .B0(n930), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n929), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15413), .COUT(n15414));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1591_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1591_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1591_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1591_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1591_add_4_4 (.A0(d_out_d_11__N_1892[17]), .B0(ISquare[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1892[17]), .B1(n931), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15412), .COUT(n15413));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1591_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1591_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1591_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1591_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1591_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15412));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[15:27])
    defparam _add_1_1591_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1591_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1591_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1591_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15411), .S0(cout_adj_5288));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1418_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1418_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_36 (.A0(d4[34]), .B0(d3[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[35]), .B1(d3[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15410), .COUT(n15411), .S0(d4_71__N_634[34]), .S1(d4_71__N_634[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_34 (.A0(d4[32]), .B0(d3[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[33]), .B1(d3[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15409), .COUT(n15410), .S0(d4_71__N_634[32]), .S1(d4_71__N_634[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_32 (.A0(d4[30]), .B0(d3[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[31]), .B1(d3[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15408), .COUT(n15409), .S0(d4_71__N_634[30]), .S1(d4_71__N_634[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_30 (.A0(d4[28]), .B0(d3[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[29]), .B1(d3[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15407), .COUT(n15408), .S0(d4_71__N_634[28]), .S1(d4_71__N_634[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_28 (.A0(d4[26]), .B0(d3[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[27]), .B1(d3[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15406), .COUT(n15407), .S0(d4_71__N_634[26]), .S1(d4_71__N_634[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_26 (.A0(d4[24]), .B0(d3[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[25]), .B1(d3[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15405), .COUT(n15406), .S0(d4_71__N_634[24]), .S1(d4_71__N_634[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_24 (.A0(d4[22]), .B0(d3[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[23]), .B1(d3[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15404), .COUT(n15405), .S0(d4_71__N_634[22]), .S1(d4_71__N_634[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_22 (.A0(d4[20]), .B0(d3[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[21]), .B1(d3[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15403), .COUT(n15404), .S0(d4_71__N_634[20]), .S1(d4_71__N_634[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_20 (.A0(d4[18]), .B0(d3[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[19]), .B1(d3[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15402), .COUT(n15403), .S0(d4_71__N_634[18]), .S1(d4_71__N_634[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_18 (.A0(d4[16]), .B0(d3[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[17]), .B1(d3[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15401), .COUT(n15402), .S0(d4_71__N_634[16]), .S1(d4_71__N_634[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_16 (.A0(d4[14]), .B0(d3[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[15]), .B1(d3[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15400), .COUT(n15401), .S0(d4_71__N_634[14]), .S1(d4_71__N_634[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_14 (.A0(d4[12]), .B0(d3[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[13]), .B1(d3[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15399), .COUT(n15400), .S0(d4_71__N_634[12]), .S1(d4_71__N_634[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_12 (.A0(d4[10]), .B0(d3[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[11]), .B1(d3[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15398), .COUT(n15399), .S0(d4_71__N_634[10]), .S1(d4_71__N_634[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_10 (.A0(d4[8]), .B0(d3[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d4[9]), .B1(d3[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15397), .COUT(n15398), .S0(d4_71__N_634[8]), .S1(d4_71__N_634[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_8 (.A0(d4[6]), .B0(d3[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[7]), .B1(d3[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15396), 
          .COUT(n15397), .S0(d4_71__N_634[6]), .S1(d4_71__N_634[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_6 (.A0(d4[4]), .B0(d3[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[5]), .B1(d3[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15395), 
          .COUT(n15396), .S0(d4_71__N_634[4]), .S1(d4_71__N_634[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_4 (.A0(d4[2]), .B0(d3[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[3]), .B1(d3[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15394), 
          .COUT(n15395), .S0(d4_71__N_634[2]), .S1(d4_71__N_634[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1418_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1418_add_4_2 (.A0(d4[0]), .B0(d3[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d4[1]), .B1(d3[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15394), 
          .S1(d4_71__N_634[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1418_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1418_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1418_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1418_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_38 (.A0(d1[71]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15392), .S0(n78_adj_5289));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1555_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_36 (.A0(d1[69]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[70]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15391), .COUT(n15392), .S0(n84_adj_5291), 
          .S1(n81_adj_5290));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_34 (.A0(d1[67]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[68]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15390), .COUT(n15391), .S0(n90_adj_5293), 
          .S1(n87_adj_5292));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_32 (.A0(d1[65]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[66]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15389), .COUT(n15390), .S0(n96_adj_5295), 
          .S1(n93_adj_5294));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_30 (.A0(d1[63]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[64]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15388), .COUT(n15389), .S0(n102_adj_5297), 
          .S1(n99_adj_5296));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_28 (.A0(d1[61]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[62]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15387), .COUT(n15388), .S0(n108_adj_5299), 
          .S1(n105_adj_5298));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_26 (.A0(d1[59]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[60]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15386), .COUT(n15387), .S0(n114_adj_5301), 
          .S1(n111_adj_5300));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_24 (.A0(d1[57]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[58]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15385), .COUT(n15386), .S0(n120_adj_5303), 
          .S1(n117_adj_5302));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_22 (.A0(d1[55]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[56]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15384), .COUT(n15385), .S0(n126_adj_5305), 
          .S1(n123_adj_5304));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_20 (.A0(d1[53]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[54]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15383), .COUT(n15384), .S0(n132_adj_5307), 
          .S1(n129_adj_5306));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_18 (.A0(d1[51]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[52]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15382), .COUT(n15383), .S0(n138_adj_5309), 
          .S1(n135_adj_5308));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_16 (.A0(d1[49]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[50]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15381), .COUT(n15382), .S0(n144_adj_5311), 
          .S1(n141_adj_5310));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_14 (.A0(d1[47]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[48]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15380), .COUT(n15381), .S0(n150_adj_5313), 
          .S1(n147_adj_5312));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_12 (.A0(d1[45]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[46]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15379), .COUT(n15380), .S0(n156_adj_5315), 
          .S1(n153_adj_5314));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_10 (.A0(d1[43]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[44]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15378), .COUT(n15379), .S0(n162_adj_5317), 
          .S1(n159_adj_5316));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_8 (.A0(d1[41]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[42]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15377), .COUT(n15378), .S0(n168_adj_5319), 
          .S1(n165_adj_5318));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_6 (.A0(d1[39]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[40]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15376), .COUT(n15377), .S0(n174_adj_5321), 
          .S1(n171_adj_5320));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_4 (.A0(d1[37]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[38]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15375), .COUT(n15376), .S0(n180_adj_5323), 
          .S1(n177_adj_5322));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1555_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1555_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[36]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15375), .S1(n183_adj_5324));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1555_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1555_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1555_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1555_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15374), .S0(cout_adj_2824));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1412_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1412_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_36 (.A0(d2[34]), .B0(d1[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[35]), .B1(d1[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15373), .COUT(n15374), .S0(d2_71__N_490[34]), .S1(d2_71__N_490[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_34 (.A0(d2[32]), .B0(d1[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[33]), .B1(d1[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15372), .COUT(n15373), .S0(d2_71__N_490[32]), .S1(d2_71__N_490[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_32 (.A0(d2[30]), .B0(d1[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[31]), .B1(d1[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15371), .COUT(n15372), .S0(d2_71__N_490[30]), .S1(d2_71__N_490[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_30 (.A0(d2[28]), .B0(d1[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[29]), .B1(d1[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15370), .COUT(n15371), .S0(d2_71__N_490[28]), .S1(d2_71__N_490[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_28 (.A0(d2[26]), .B0(d1[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[27]), .B1(d1[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15369), .COUT(n15370), .S0(d2_71__N_490[26]), .S1(d2_71__N_490[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_26 (.A0(d2[24]), .B0(d1[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[25]), .B1(d1[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15368), .COUT(n15369), .S0(d2_71__N_490[24]), .S1(d2_71__N_490[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_24 (.A0(d2[22]), .B0(d1[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[23]), .B1(d1[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15367), .COUT(n15368), .S0(d2_71__N_490[22]), .S1(d2_71__N_490[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_22 (.A0(d2[20]), .B0(d1[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[21]), .B1(d1[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15366), .COUT(n15367), .S0(d2_71__N_490[20]), .S1(d2_71__N_490[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_20 (.A0(d2[18]), .B0(d1[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[19]), .B1(d1[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15365), .COUT(n15366), .S0(d2_71__N_490[18]), .S1(d2_71__N_490[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_18 (.A0(d2[16]), .B0(d1[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[17]), .B1(d1[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15364), .COUT(n15365), .S0(d2_71__N_490[16]), .S1(d2_71__N_490[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_16 (.A0(d2[14]), .B0(d1[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[15]), .B1(d1[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15363), .COUT(n15364), .S0(d2_71__N_490[14]), .S1(d2_71__N_490[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_14 (.A0(d2[12]), .B0(d1[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[13]), .B1(d1[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15362), .COUT(n15363), .S0(d2_71__N_490[12]), .S1(d2_71__N_490[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_12 (.A0(d2[10]), .B0(d1[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[11]), .B1(d1[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15361), .COUT(n15362), .S0(d2_71__N_490[10]), .S1(d2_71__N_490[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_10 (.A0(d2[8]), .B0(d1[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d2[9]), .B1(d1[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15360), .COUT(n15361), .S0(d2_71__N_490[8]), .S1(d2_71__N_490[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_8 (.A0(d2[6]), .B0(d1[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[7]), .B1(d1[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15359), 
          .COUT(n15360), .S0(d2_71__N_490[6]), .S1(d2_71__N_490[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_6 (.A0(d2[4]), .B0(d1[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[5]), .B1(d1[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15358), 
          .COUT(n15359), .S0(d2_71__N_490[4]), .S1(d2_71__N_490[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_4 (.A0(d2[2]), .B0(d1[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[3]), .B1(d1[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15357), 
          .COUT(n15358), .S0(d2_71__N_490[2]), .S1(d2_71__N_490[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1412_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1412_add_4_2 (.A0(d2[0]), .B0(d1[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d2[1]), .B1(d1[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15357), 
          .S1(d2_71__N_490[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1412_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1412_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1412_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1412_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_37 (.A0(d2[70]), .B0(cout), .C0(n81_adj_5553), 
          .D0(d3[70]), .A1(d2[71]), .B1(cout), .C1(n78_adj_5552), .D1(d3[71]), 
          .CIN(n15354), .S0(d3_71__N_562[70]), .S1(d3_71__N_562[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_35 (.A0(d2[68]), .B0(cout), .C0(n87_adj_5555), 
          .D0(d3[68]), .A1(d2[69]), .B1(cout), .C1(n84_adj_5554), .D1(d3[69]), 
          .CIN(n15353), .COUT(n15354), .S0(d3_71__N_562[68]), .S1(d3_71__N_562[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_33 (.A0(d2[66]), .B0(cout), .C0(n93_adj_5557), 
          .D0(d3[66]), .A1(d2[67]), .B1(cout), .C1(n90_adj_5556), .D1(d3[67]), 
          .CIN(n15352), .COUT(n15353), .S0(d3_71__N_562[66]), .S1(d3_71__N_562[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_31 (.A0(d2[64]), .B0(cout), .C0(n99_adj_5559), 
          .D0(d3[64]), .A1(d2[65]), .B1(cout), .C1(n96_adj_5558), .D1(d3[65]), 
          .CIN(n15351), .COUT(n15352), .S0(d3_71__N_562[64]), .S1(d3_71__N_562[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_29 (.A0(d2[62]), .B0(cout), .C0(n105_adj_5561), 
          .D0(d3[62]), .A1(d2[63]), .B1(cout), .C1(n102_adj_5560), .D1(d3[63]), 
          .CIN(n15350), .COUT(n15351), .S0(d3_71__N_562[62]), .S1(d3_71__N_562[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_27 (.A0(d2[60]), .B0(cout), .C0(n111_adj_5563), 
          .D0(d3[60]), .A1(d2[61]), .B1(cout), .C1(n108_adj_5562), .D1(d3[61]), 
          .CIN(n15349), .COUT(n15350), .S0(d3_71__N_562[60]), .S1(d3_71__N_562[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_25 (.A0(d2[58]), .B0(cout), .C0(n117_adj_5565), 
          .D0(d3[58]), .A1(d2[59]), .B1(cout), .C1(n114_adj_5564), .D1(d3[59]), 
          .CIN(n15348), .COUT(n15349), .S0(d3_71__N_562[58]), .S1(d3_71__N_562[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_23 (.A0(d2[56]), .B0(cout), .C0(n123_adj_5567), 
          .D0(d3[56]), .A1(d2[57]), .B1(cout), .C1(n120_adj_5566), .D1(d3[57]), 
          .CIN(n15347), .COUT(n15348), .S0(d3_71__N_562[56]), .S1(d3_71__N_562[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_21 (.A0(d2[54]), .B0(cout), .C0(n129_adj_5569), 
          .D0(d3[54]), .A1(d2[55]), .B1(cout), .C1(n126_adj_5568), .D1(d3[55]), 
          .CIN(n15346), .COUT(n15347), .S0(d3_71__N_562[54]), .S1(d3_71__N_562[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_19 (.A0(d2[52]), .B0(cout), .C0(n135_adj_5571), 
          .D0(d3[52]), .A1(d2[53]), .B1(cout), .C1(n132_adj_5570), .D1(d3[53]), 
          .CIN(n15345), .COUT(n15346), .S0(d3_71__N_562[52]), .S1(d3_71__N_562[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_17 (.A0(d2[50]), .B0(cout), .C0(n141_adj_5573), 
          .D0(d3[50]), .A1(d2[51]), .B1(cout), .C1(n138_adj_5572), .D1(d3[51]), 
          .CIN(n15344), .COUT(n15345), .S0(d3_71__N_562[50]), .S1(d3_71__N_562[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_15 (.A0(d2[48]), .B0(cout), .C0(n147_adj_5575), 
          .D0(d3[48]), .A1(d2[49]), .B1(cout), .C1(n144_adj_5574), .D1(d3[49]), 
          .CIN(n15343), .COUT(n15344), .S0(d3_71__N_562[48]), .S1(d3_71__N_562[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_13 (.A0(d2[46]), .B0(cout), .C0(n153_adj_5577), 
          .D0(d3[46]), .A1(d2[47]), .B1(cout), .C1(n150_adj_5576), .D1(d3[47]), 
          .CIN(n15342), .COUT(n15343), .S0(d3_71__N_562[46]), .S1(d3_71__N_562[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_11 (.A0(d2[44]), .B0(cout), .C0(n159_adj_5579), 
          .D0(d3[44]), .A1(d2[45]), .B1(cout), .C1(n156_adj_5578), .D1(d3[45]), 
          .CIN(n15341), .COUT(n15342), .S0(d3_71__N_562[44]), .S1(d3_71__N_562[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_9 (.A0(d2[42]), .B0(cout), .C0(n165_adj_5581), 
          .D0(d3[42]), .A1(d2[43]), .B1(cout), .C1(n162_adj_5580), .D1(d3[43]), 
          .CIN(n15340), .COUT(n15341), .S0(d3_71__N_562[42]), .S1(d3_71__N_562[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_7 (.A0(d2[40]), .B0(cout), .C0(n171_adj_5583), 
          .D0(d3[40]), .A1(d2[41]), .B1(cout), .C1(n168_adj_5582), .D1(d3[41]), 
          .CIN(n15339), .COUT(n15340), .S0(d3_71__N_562[40]), .S1(d3_71__N_562[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_5 (.A0(d2[38]), .B0(cout), .C0(n177_adj_5585), 
          .D0(d3[38]), .A1(d2[39]), .B1(cout), .C1(n174_adj_5584), .D1(d3[39]), 
          .CIN(n15338), .COUT(n15339), .S0(d3_71__N_562[38]), .S1(d3_71__N_562[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_3 (.A0(d2[36]), .B0(cout), .C0(n183_adj_5587), 
          .D0(d3[36]), .A1(d2[37]), .B1(cout), .C1(n180_adj_5586), .D1(d3[37]), 
          .CIN(n15337), .COUT(n15338), .S0(d3_71__N_562[36]), .S1(d3_71__N_562[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1513_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1513_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1513_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15337));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1513_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1513_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1513_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1513_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_37 (.A0(d3_adj_5742[70]), .B0(cout_adj_5362), 
          .C0(n81_adj_5151), .D0(d4_adj_5743[70]), .A1(d3_adj_5742[71]), 
          .B1(cout_adj_5362), .C1(n78_adj_5150), .D1(d4_adj_5743[71]), 
          .CIN(n15332), .S0(d4_71__N_634_adj_5759[70]), .S1(d4_71__N_634_adj_5759[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_35 (.A0(d3_adj_5742[68]), .B0(cout_adj_5362), 
          .C0(n87_adj_5153), .D0(d4_adj_5743[68]), .A1(d3_adj_5742[69]), 
          .B1(cout_adj_5362), .C1(n84_adj_5152), .D1(d4_adj_5743[69]), 
          .CIN(n15331), .COUT(n15332), .S0(d4_71__N_634_adj_5759[68]), 
          .S1(d4_71__N_634_adj_5759[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_33 (.A0(d3_adj_5742[66]), .B0(cout_adj_5362), 
          .C0(n93_adj_5155), .D0(d4_adj_5743[66]), .A1(d3_adj_5742[67]), 
          .B1(cout_adj_5362), .C1(n90_adj_5154), .D1(d4_adj_5743[67]), 
          .CIN(n15330), .COUT(n15331), .S0(d4_71__N_634_adj_5759[66]), 
          .S1(d4_71__N_634_adj_5759[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_31 (.A0(d3_adj_5742[64]), .B0(cout_adj_5362), 
          .C0(n99_adj_5157), .D0(d4_adj_5743[64]), .A1(d3_adj_5742[65]), 
          .B1(cout_adj_5362), .C1(n96_adj_5156), .D1(d4_adj_5743[65]), 
          .CIN(n15329), .COUT(n15330), .S0(d4_71__N_634_adj_5759[64]), 
          .S1(d4_71__N_634_adj_5759[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_29 (.A0(d3_adj_5742[62]), .B0(cout_adj_5362), 
          .C0(n105_adj_5159), .D0(d4_adj_5743[62]), .A1(d3_adj_5742[63]), 
          .B1(cout_adj_5362), .C1(n102_adj_5158), .D1(d4_adj_5743[63]), 
          .CIN(n15328), .COUT(n15329), .S0(d4_71__N_634_adj_5759[62]), 
          .S1(d4_71__N_634_adj_5759[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_27 (.A0(d3_adj_5742[60]), .B0(cout_adj_5362), 
          .C0(n111_adj_5161), .D0(d4_adj_5743[60]), .A1(d3_adj_5742[61]), 
          .B1(cout_adj_5362), .C1(n108_adj_5160), .D1(d4_adj_5743[61]), 
          .CIN(n15327), .COUT(n15328), .S0(d4_71__N_634_adj_5759[60]), 
          .S1(d4_71__N_634_adj_5759[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_25 (.A0(d3_adj_5742[58]), .B0(cout_adj_5362), 
          .C0(n117_adj_5163), .D0(d4_adj_5743[58]), .A1(d3_adj_5742[59]), 
          .B1(cout_adj_5362), .C1(n114_adj_5162), .D1(d4_adj_5743[59]), 
          .CIN(n15326), .COUT(n15327), .S0(d4_71__N_634_adj_5759[58]), 
          .S1(d4_71__N_634_adj_5759[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_23 (.A0(d3_adj_5742[56]), .B0(cout_adj_5362), 
          .C0(n123_adj_5165), .D0(d4_adj_5743[56]), .A1(d3_adj_5742[57]), 
          .B1(cout_adj_5362), .C1(n120_adj_5164), .D1(d4_adj_5743[57]), 
          .CIN(n15325), .COUT(n15326), .S0(d4_71__N_634_adj_5759[56]), 
          .S1(d4_71__N_634_adj_5759[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_21 (.A0(d3_adj_5742[54]), .B0(cout_adj_5362), 
          .C0(n129_adj_5167), .D0(d4_adj_5743[54]), .A1(d3_adj_5742[55]), 
          .B1(cout_adj_5362), .C1(n126_adj_5166), .D1(d4_adj_5743[55]), 
          .CIN(n15324), .COUT(n15325), .S0(d4_71__N_634_adj_5759[54]), 
          .S1(d4_71__N_634_adj_5759[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_19 (.A0(d3_adj_5742[52]), .B0(cout_adj_5362), 
          .C0(n135_adj_5169), .D0(d4_adj_5743[52]), .A1(d3_adj_5742[53]), 
          .B1(cout_adj_5362), .C1(n132_adj_5168), .D1(d4_adj_5743[53]), 
          .CIN(n15323), .COUT(n15324), .S0(d4_71__N_634_adj_5759[52]), 
          .S1(d4_71__N_634_adj_5759[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_17 (.A0(d3_adj_5742[50]), .B0(cout_adj_5362), 
          .C0(n141_adj_5171), .D0(d4_adj_5743[50]), .A1(d3_adj_5742[51]), 
          .B1(cout_adj_5362), .C1(n138_adj_5170), .D1(d4_adj_5743[51]), 
          .CIN(n15322), .COUT(n15323), .S0(d4_71__N_634_adj_5759[50]), 
          .S1(d4_71__N_634_adj_5759[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_15 (.A0(d3_adj_5742[48]), .B0(cout_adj_5362), 
          .C0(n147_adj_5173), .D0(d4_adj_5743[48]), .A1(d3_adj_5742[49]), 
          .B1(cout_adj_5362), .C1(n144_adj_5172), .D1(d4_adj_5743[49]), 
          .CIN(n15321), .COUT(n15322), .S0(d4_71__N_634_adj_5759[48]), 
          .S1(d4_71__N_634_adj_5759[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_13 (.A0(d3_adj_5742[46]), .B0(cout_adj_5362), 
          .C0(n153_adj_5175), .D0(d4_adj_5743[46]), .A1(d3_adj_5742[47]), 
          .B1(cout_adj_5362), .C1(n150_adj_5174), .D1(d4_adj_5743[47]), 
          .CIN(n15320), .COUT(n15321), .S0(d4_71__N_634_adj_5759[46]), 
          .S1(d4_71__N_634_adj_5759[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_11 (.A0(d3_adj_5742[44]), .B0(cout_adj_5362), 
          .C0(n159_adj_5177), .D0(d4_adj_5743[44]), .A1(d3_adj_5742[45]), 
          .B1(cout_adj_5362), .C1(n156_adj_5176), .D1(d4_adj_5743[45]), 
          .CIN(n15319), .COUT(n15320), .S0(d4_71__N_634_adj_5759[44]), 
          .S1(d4_71__N_634_adj_5759[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_9 (.A0(d3_adj_5742[42]), .B0(cout_adj_5362), 
          .C0(n165_adj_5179), .D0(d4_adj_5743[42]), .A1(d3_adj_5742[43]), 
          .B1(cout_adj_5362), .C1(n162_adj_5178), .D1(d4_adj_5743[43]), 
          .CIN(n15318), .COUT(n15319), .S0(d4_71__N_634_adj_5759[42]), 
          .S1(d4_71__N_634_adj_5759[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_7 (.A0(d3_adj_5742[40]), .B0(cout_adj_5362), 
          .C0(n171_adj_5181), .D0(d4_adj_5743[40]), .A1(d3_adj_5742[41]), 
          .B1(cout_adj_5362), .C1(n168_adj_5180), .D1(d4_adj_5743[41]), 
          .CIN(n15317), .COUT(n15318), .S0(d4_71__N_634_adj_5759[40]), 
          .S1(d4_71__N_634_adj_5759[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_5 (.A0(d3_adj_5742[38]), .B0(cout_adj_5362), 
          .C0(n177_adj_5183), .D0(d4_adj_5743[38]), .A1(d3_adj_5742[39]), 
          .B1(cout_adj_5362), .C1(n174_adj_5182), .D1(d4_adj_5743[39]), 
          .CIN(n15316), .COUT(n15317), .S0(d4_71__N_634_adj_5759[38]), 
          .S1(d4_71__N_634_adj_5759[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_3 (.A0(d3_adj_5742[36]), .B0(cout_adj_5362), 
          .C0(n183_adj_5185), .D0(d4_adj_5743[36]), .A1(d3_adj_5742[37]), 
          .B1(cout_adj_5362), .C1(n180_adj_5184), .D1(d4_adj_5743[37]), 
          .CIN(n15315), .COUT(n15316), .S0(d4_71__N_634_adj_5759[36]), 
          .S1(d4_71__N_634_adj_5759[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1495_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1495_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1495_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5362), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15315));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(65[15:24])
    defparam _add_1_1495_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1495_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1495_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1495_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15311), .S0(cout));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1415_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1415_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_36 (.A0(d3[34]), .B0(d2[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[35]), .B1(d2[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15310), .COUT(n15311), .S0(d3_71__N_562[34]), .S1(d3_71__N_562[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_34 (.A0(d3[32]), .B0(d2[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[33]), .B1(d2[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15309), .COUT(n15310), .S0(d3_71__N_562[32]), .S1(d3_71__N_562[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_32 (.A0(d3[30]), .B0(d2[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[31]), .B1(d2[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15308), .COUT(n15309), .S0(d3_71__N_562[30]), .S1(d3_71__N_562[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_30 (.A0(d3[28]), .B0(d2[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[29]), .B1(d2[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15307), .COUT(n15308), .S0(d3_71__N_562[28]), .S1(d3_71__N_562[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_28 (.A0(d3[26]), .B0(d2[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[27]), .B1(d2[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15306), .COUT(n15307), .S0(d3_71__N_562[26]), .S1(d3_71__N_562[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_26 (.A0(d3[24]), .B0(d2[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[25]), .B1(d2[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15305), .COUT(n15306), .S0(d3_71__N_562[24]), .S1(d3_71__N_562[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_24 (.A0(d3[22]), .B0(d2[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[23]), .B1(d2[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15304), .COUT(n15305), .S0(d3_71__N_562[22]), .S1(d3_71__N_562[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_22 (.A0(d3[20]), .B0(d2[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[21]), .B1(d2[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15303), .COUT(n15304), .S0(d3_71__N_562[20]), .S1(d3_71__N_562[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_20 (.A0(d3[18]), .B0(d2[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[19]), .B1(d2[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15302), .COUT(n15303), .S0(d3_71__N_562[18]), .S1(d3_71__N_562[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_18 (.A0(d3[16]), .B0(d2[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[17]), .B1(d2[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15301), .COUT(n15302), .S0(d3_71__N_562[16]), .S1(d3_71__N_562[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_16 (.A0(d3[14]), .B0(d2[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[15]), .B1(d2[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15300), .COUT(n15301), .S0(d3_71__N_562[14]), .S1(d3_71__N_562[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_14 (.A0(d3[12]), .B0(d2[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[13]), .B1(d2[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15299), .COUT(n15300), .S0(d3_71__N_562[12]), .S1(d3_71__N_562[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_12 (.A0(d3[10]), .B0(d2[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[11]), .B1(d2[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15298), .COUT(n15299), .S0(d3_71__N_562[10]), .S1(d3_71__N_562[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_10 (.A0(d3[8]), .B0(d2[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[9]), .B1(d2[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15297), .COUT(n15298), .S0(d3_71__N_562[8]), .S1(d3_71__N_562[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_8 (.A0(d3[6]), .B0(d2[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[7]), .B1(d2[7]), .C1(GND_net), .D1(VCC_net), .CIN(n15296), 
          .COUT(n15297), .S0(d3_71__N_562[6]), .S1(d3_71__N_562[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_6 (.A0(d3[4]), .B0(d2[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[5]), .B1(d2[5]), .C1(GND_net), .D1(VCC_net), .CIN(n15295), 
          .COUT(n15296), .S0(d3_71__N_562[4]), .S1(d3_71__N_562[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_4 (.A0(d3[2]), .B0(d2[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[3]), .B1(d2[3]), .C1(GND_net), .D1(VCC_net), .CIN(n15294), 
          .COUT(n15295), .S0(d3_71__N_562[2]), .S1(d3_71__N_562[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1415_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1415_add_4_2 (.A0(d3[0]), .B0(d2[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d3[1]), .B1(d2[1]), .C1(GND_net), .D1(VCC_net), .COUT(n15294), 
          .S1(d3_71__N_562[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1415_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1415_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1415_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1415_add_4_2.INJECT1_1 = "NO";
    LUT4 i5418_4_lut_rep_227 (.A(n17401), .B(n17940), .C(n17906), .D(n17777), 
         .Z(clk_80mhz_enable_1459)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C))) */ ;
    defparam i5418_4_lut_rep_227.init = 16'hc0c8;
    CCU2C _add_1_1603_add_4_38 (.A0(d_d9_adj_5752[35]), .B0(d9_adj_5751[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15292), .S1(cout_adj_5516));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1603_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_36 (.A0(d_d9_adj_5752[33]), .B0(d9_adj_5751[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[34]), .B1(d9_adj_5751[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15291), .COUT(n15292));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_34 (.A0(d_d9_adj_5752[31]), .B0(d9_adj_5751[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[32]), .B1(d9_adj_5751[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15290), .COUT(n15291));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_32 (.A0(d_d9_adj_5752[29]), .B0(d9_adj_5751[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[30]), .B1(d9_adj_5751[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15289), .COUT(n15290));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_30 (.A0(d_d9_adj_5752[27]), .B0(d9_adj_5751[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[28]), .B1(d9_adj_5751[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15288), .COUT(n15289));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_28 (.A0(d_d9_adj_5752[25]), .B0(d9_adj_5751[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[26]), .B1(d9_adj_5751[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15287), .COUT(n15288));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_26 (.A0(d_d9_adj_5752[23]), .B0(d9_adj_5751[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[24]), .B1(d9_adj_5751[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15286), .COUT(n15287));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_24 (.A0(d_d9_adj_5752[21]), .B0(d9_adj_5751[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[22]), .B1(d9_adj_5751[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15285), .COUT(n15286));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_22 (.A0(d_d9_adj_5752[19]), .B0(d9_adj_5751[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[20]), .B1(d9_adj_5751[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15284), .COUT(n15285));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_20 (.A0(d_d9_adj_5752[17]), .B0(d9_adj_5751[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[18]), .B1(d9_adj_5751[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15283), .COUT(n15284));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_18 (.A0(d_d9_adj_5752[15]), .B0(d9_adj_5751[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[16]), .B1(d9_adj_5751[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15282), .COUT(n15283));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_16 (.A0(d_d9_adj_5752[13]), .B0(d9_adj_5751[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[14]), .B1(d9_adj_5751[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15281), .COUT(n15282));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_14 (.A0(d_d9_adj_5752[11]), .B0(d9_adj_5751[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[12]), .B1(d9_adj_5751[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15280), .COUT(n15281));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_12 (.A0(d_d9_adj_5752[9]), .B0(d9_adj_5751[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[10]), .B1(d9_adj_5751[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15279), .COUT(n15280));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_10 (.A0(d_d9_adj_5752[7]), .B0(d9_adj_5751[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[8]), .B1(d9_adj_5751[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15278), .COUT(n15279));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_8 (.A0(d_d9_adj_5752[5]), .B0(d9_adj_5751[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[6]), .B1(d9_adj_5751[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15277), .COUT(n15278));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_6 (.A0(d_d9_adj_5752[3]), .B0(d9_adj_5751[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[4]), .B1(d9_adj_5751[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15276), .COUT(n15277));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_4 (.A0(d_d9_adj_5752[1]), .B0(d9_adj_5751[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[2]), .B1(d9_adj_5751[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15275), .COUT(n15276));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1603_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1603_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9_adj_5752[0]), .B1(d9_adj_5751[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15275));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1603_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1603_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1603_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1603_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_38 (.A0(d_d7_adj_5748[35]), .B0(d7_adj_5747[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15274), .S0(d8_71__N_1603_adj_5774[35]), 
          .S1(cout_adj_5613));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1612_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_36 (.A0(d_d7_adj_5748[33]), .B0(d7_adj_5747[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[34]), .B1(d7_adj_5747[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15273), .COUT(n15274), .S0(d8_71__N_1603_adj_5774[33]), 
          .S1(d8_71__N_1603_adj_5774[34]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_34 (.A0(d_d7_adj_5748[31]), .B0(d7_adj_5747[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[32]), .B1(d7_adj_5747[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15272), .COUT(n15273), .S0(d8_71__N_1603_adj_5774[31]), 
          .S1(d8_71__N_1603_adj_5774[32]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_32 (.A0(d_d7_adj_5748[29]), .B0(d7_adj_5747[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[30]), .B1(d7_adj_5747[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15271), .COUT(n15272), .S0(d8_71__N_1603_adj_5774[29]), 
          .S1(d8_71__N_1603_adj_5774[30]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_30 (.A0(d_d7_adj_5748[27]), .B0(d7_adj_5747[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[28]), .B1(d7_adj_5747[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15270), .COUT(n15271), .S0(d8_71__N_1603_adj_5774[27]), 
          .S1(d8_71__N_1603_adj_5774[28]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_28 (.A0(d_d7_adj_5748[25]), .B0(d7_adj_5747[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[26]), .B1(d7_adj_5747[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15269), .COUT(n15270), .S0(d8_71__N_1603_adj_5774[25]), 
          .S1(d8_71__N_1603_adj_5774[26]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_26 (.A0(d_d7_adj_5748[23]), .B0(d7_adj_5747[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[24]), .B1(d7_adj_5747[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15268), .COUT(n15269), .S0(d8_71__N_1603_adj_5774[23]), 
          .S1(d8_71__N_1603_adj_5774[24]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_24 (.A0(d_d7_adj_5748[21]), .B0(d7_adj_5747[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[22]), .B1(d7_adj_5747[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15267), .COUT(n15268), .S0(d8_71__N_1603_adj_5774[21]), 
          .S1(d8_71__N_1603_adj_5774[22]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_22 (.A0(d_d7_adj_5748[19]), .B0(d7_adj_5747[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[20]), .B1(d7_adj_5747[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15266), .COUT(n15267), .S0(d8_71__N_1603_adj_5774[19]), 
          .S1(d8_71__N_1603_adj_5774[20]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_20 (.A0(d_d7_adj_5748[17]), .B0(d7_adj_5747[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[18]), .B1(d7_adj_5747[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15265), .COUT(n15266), .S0(d8_71__N_1603_adj_5774[17]), 
          .S1(d8_71__N_1603_adj_5774[18]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_18 (.A0(d_d7_adj_5748[15]), .B0(d7_adj_5747[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[16]), .B1(d7_adj_5747[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15264), .COUT(n15265), .S0(d8_71__N_1603_adj_5774[15]), 
          .S1(d8_71__N_1603_adj_5774[16]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_16 (.A0(d_d7_adj_5748[13]), .B0(d7_adj_5747[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[14]), .B1(d7_adj_5747[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15263), .COUT(n15264), .S0(d8_71__N_1603_adj_5774[13]), 
          .S1(d8_71__N_1603_adj_5774[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_14 (.A0(d_d7_adj_5748[11]), .B0(d7_adj_5747[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[12]), .B1(d7_adj_5747[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15262), .COUT(n15263), .S0(d8_71__N_1603_adj_5774[11]), 
          .S1(d8_71__N_1603_adj_5774[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_12 (.A0(d_d7_adj_5748[9]), .B0(d7_adj_5747[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[10]), .B1(d7_adj_5747[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15261), .COUT(n15262), .S0(d8_71__N_1603_adj_5774[9]), 
          .S1(d8_71__N_1603_adj_5774[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_10 (.A0(d_d7_adj_5748[7]), .B0(d7_adj_5747[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[8]), .B1(d7_adj_5747[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15260), .COUT(n15261), .S0(d8_71__N_1603_adj_5774[7]), 
          .S1(d8_71__N_1603_adj_5774[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_8 (.A0(d_d7_adj_5748[5]), .B0(d7_adj_5747[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[6]), .B1(d7_adj_5747[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15259), .COUT(n15260), .S0(d8_71__N_1603_adj_5774[5]), 
          .S1(d8_71__N_1603_adj_5774[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_6 (.A0(d_d7_adj_5748[3]), .B0(d7_adj_5747[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[4]), .B1(d7_adj_5747[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15258), .COUT(n15259), .S0(d8_71__N_1603_adj_5774[3]), 
          .S1(d8_71__N_1603_adj_5774[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_4 (.A0(d_d7_adj_5748[1]), .B0(d7_adj_5747[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[2]), .B1(d7_adj_5747[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15257), .COUT(n15258), .S0(d8_71__N_1603_adj_5774[1]), 
          .S1(d8_71__N_1603_adj_5774[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1612_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1612_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d7_adj_5748[0]), .B1(d7_adj_5747[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15257), .S1(d8_71__N_1603_adj_5774[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1612_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1612_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1612_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1612_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_38 (.A0(d_d_tmp_adj_5739[71]), .B0(d_tmp_adj_5738[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15256), .S0(n78_adj_4880));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1630_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_36 (.A0(d_d_tmp_adj_5739[69]), .B0(d_tmp_adj_5738[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[70]), .B1(d_tmp_adj_5738[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15255), .COUT(n15256), .S0(n84_adj_4882), 
          .S1(n81_adj_4881));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_34 (.A0(d_d_tmp_adj_5739[67]), .B0(d_tmp_adj_5738[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[68]), .B1(d_tmp_adj_5738[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15254), .COUT(n15255), .S0(n90_adj_4884), 
          .S1(n87_adj_4883));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_32 (.A0(d_d_tmp_adj_5739[65]), .B0(d_tmp_adj_5738[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[66]), .B1(d_tmp_adj_5738[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15253), .COUT(n15254), .S0(n96_adj_4886), 
          .S1(n93_adj_4885));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_30 (.A0(d_d_tmp_adj_5739[63]), .B0(d_tmp_adj_5738[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[64]), .B1(d_tmp_adj_5738[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15252), .COUT(n15253), .S0(n102_adj_4888), 
          .S1(n99_adj_4887));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_28 (.A0(d_d_tmp_adj_5739[61]), .B0(d_tmp_adj_5738[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[62]), .B1(d_tmp_adj_5738[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15251), .COUT(n15252), .S0(n108_adj_4890), 
          .S1(n105_adj_4889));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_26 (.A0(d_d_tmp_adj_5739[59]), .B0(d_tmp_adj_5738[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[60]), .B1(d_tmp_adj_5738[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15250), .COUT(n15251), .S0(n114_adj_4892), 
          .S1(n111_adj_4891));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_24 (.A0(d_d_tmp_adj_5739[57]), .B0(d_tmp_adj_5738[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[58]), .B1(d_tmp_adj_5738[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15249), .COUT(n15250), .S0(n120_adj_4894), 
          .S1(n117_adj_4893));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_22 (.A0(d_d_tmp_adj_5739[55]), .B0(d_tmp_adj_5738[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[56]), .B1(d_tmp_adj_5738[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15248), .COUT(n15249), .S0(n126_adj_4896), 
          .S1(n123_adj_4895));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_20 (.A0(d_d_tmp_adj_5739[53]), .B0(d_tmp_adj_5738[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[54]), .B1(d_tmp_adj_5738[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15247), .COUT(n15248), .S0(n132_adj_4898), 
          .S1(n129_adj_4897));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_18 (.A0(d_d_tmp_adj_5739[51]), .B0(d_tmp_adj_5738[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[52]), .B1(d_tmp_adj_5738[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15246), .COUT(n15247), .S0(n138_adj_4900), 
          .S1(n135_adj_4899));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_16 (.A0(d_d_tmp_adj_5739[49]), .B0(d_tmp_adj_5738[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[50]), .B1(d_tmp_adj_5738[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15245), .COUT(n15246), .S0(n144_adj_4902), 
          .S1(n141_adj_4901));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_14 (.A0(d_d_tmp_adj_5739[47]), .B0(d_tmp_adj_5738[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[48]), .B1(d_tmp_adj_5738[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15244), .COUT(n15245), .S0(n150_adj_4904), 
          .S1(n147_adj_4903));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_12 (.A0(d_d_tmp_adj_5739[45]), .B0(d_tmp_adj_5738[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[46]), .B1(d_tmp_adj_5738[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15243), .COUT(n15244), .S0(n156_adj_4906), 
          .S1(n153_adj_4905));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_10 (.A0(d_d_tmp_adj_5739[43]), .B0(d_tmp_adj_5738[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[44]), .B1(d_tmp_adj_5738[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15242), .COUT(n15243), .S0(n162_adj_4908), 
          .S1(n159_adj_4907));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_8 (.A0(d_d_tmp_adj_5739[41]), .B0(d_tmp_adj_5738[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[42]), .B1(d_tmp_adj_5738[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15241), .COUT(n15242), .S0(n168_adj_4910), 
          .S1(n165_adj_4909));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_6 (.A0(d_d_tmp_adj_5739[39]), .B0(d_tmp_adj_5738[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[40]), .B1(d_tmp_adj_5738[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15240), .COUT(n15241), .S0(n174_adj_4912), 
          .S1(n171_adj_4911));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_4 (.A0(d_d_tmp_adj_5739[37]), .B0(d_tmp_adj_5738[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d_tmp_adj_5739[38]), .B1(d_tmp_adj_5738[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15239), .COUT(n15240), .S0(n180_adj_4914), 
          .S1(n177_adj_4913));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1630_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1630_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp_adj_5739[36]), .B1(d_tmp_adj_5738[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15239), .S1(n183_adj_4915));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1630_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1630_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1630_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1630_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1654_add_4_12 (.A0(counter[9]), .B0(DataInReg[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15238), .S1(cout_adj_5112));
    defparam _add_1_1654_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1654_add_4_12.INIT1 = 16'h0000;
    defparam _add_1_1654_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1654_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1654_add_4_10 (.A0(counter[7]), .B0(DataInReg[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[8]), .B1(DataInReg[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15237), .COUT(n15238));
    defparam _add_1_1654_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1654_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1654_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1654_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1654_add_4_8 (.A0(counter[5]), .B0(DataInReg[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[6]), .B1(DataInReg[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15236), .COUT(n15237));
    defparam _add_1_1654_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1654_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1654_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1654_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1654_add_4_6 (.A0(counter[3]), .B0(DataInReg[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[4]), .B1(DataInReg[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15235), .COUT(n15236));
    defparam _add_1_1654_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1654_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1654_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1654_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1654_add_4_4 (.A0(counter[1]), .B0(DataInReg[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[2]), .B1(DataInReg[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15234), .COUT(n15235));
    defparam _add_1_1654_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1654_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1654_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1654_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1654_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[0]), .B1(DataInReg[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15234));
    defparam _add_1_1654_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1654_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1654_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1654_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_37 (.A0(d_d9_adj_5752[71]), .B0(d9_adj_5751[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15233), .S0(n76_adj_5616));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_37.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_37.INIT1 = 16'h0000;
    defparam _add_1_1468_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_35 (.A0(d_d9_adj_5752[69]), .B0(d9_adj_5751[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[70]), .B1(d9_adj_5751[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15232), .COUT(n15233), .S0(n82_adj_5618), 
          .S1(n79_adj_5617));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_35.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_35.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_33 (.A0(d_d9_adj_5752[67]), .B0(d9_adj_5751[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[68]), .B1(d9_adj_5751[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15231), .COUT(n15232), .S0(n88_adj_5620), 
          .S1(n85_adj_5619));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_33.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_33.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_31 (.A0(d_d9_adj_5752[65]), .B0(d9_adj_5751[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[66]), .B1(d9_adj_5751[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15230), .COUT(n15231), .S0(n94_adj_5622), 
          .S1(n91_adj_5621));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_31.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_31.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_29 (.A0(d_d9_adj_5752[63]), .B0(d9_adj_5751[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[64]), .B1(d9_adj_5751[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15229), .COUT(n15230), .S0(n100_adj_5624), 
          .S1(n97_adj_5623));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_29.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_29.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_27 (.A0(d_d9_adj_5752[61]), .B0(d9_adj_5751[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[62]), .B1(d9_adj_5751[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15228), .COUT(n15229), .S0(n106_adj_5626), 
          .S1(n103_adj_5625));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_27.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_27.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_25 (.A0(d_d9_adj_5752[59]), .B0(d9_adj_5751[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[60]), .B1(d9_adj_5751[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15227), .COUT(n15228), .S0(n112_adj_5628), 
          .S1(n109_adj_5627));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_25.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_25.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_23 (.A0(d_d9_adj_5752[57]), .B0(d9_adj_5751[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[58]), .B1(d9_adj_5751[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15226), .COUT(n15227), .S0(n118_adj_5630), 
          .S1(n115_adj_5629));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_23.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_23.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_21 (.A0(d_d9_adj_5752[55]), .B0(d9_adj_5751[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[56]), .B1(d9_adj_5751[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15225), .COUT(n15226));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_21.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_21.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_19 (.A0(d_d9_adj_5752[53]), .B0(d9_adj_5751[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[54]), .B1(d9_adj_5751[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15224), .COUT(n15225));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_19.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_19.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_17 (.A0(d_d9_adj_5752[51]), .B0(d9_adj_5751[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[52]), .B1(d9_adj_5751[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15223), .COUT(n15224));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_17.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_17.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_15 (.A0(d_d9_adj_5752[49]), .B0(d9_adj_5751[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[50]), .B1(d9_adj_5751[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15222), .COUT(n15223));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_15.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_15.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_13 (.A0(d_d9_adj_5752[47]), .B0(d9_adj_5751[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[48]), .B1(d9_adj_5751[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15221), .COUT(n15222));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_13.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_13.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_11 (.A0(d_d9_adj_5752[45]), .B0(d9_adj_5751[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[46]), .B1(d9_adj_5751[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15220), .COUT(n15221));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_9 (.A0(d_d9_adj_5752[43]), .B0(d9_adj_5751[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[44]), .B1(d9_adj_5751[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15219), .COUT(n15220));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_7 (.A0(d_d9_adj_5752[41]), .B0(d9_adj_5751[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[42]), .B1(d9_adj_5751[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15218), .COUT(n15219));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_5 (.A0(d_d9_adj_5752[39]), .B0(d9_adj_5751[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[40]), .B1(d9_adj_5751[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15217), .COUT(n15218));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_3 (.A0(d_d9_adj_5752[37]), .B0(d9_adj_5751[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d9_adj_5752[38]), .B1(d9_adj_5751[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15216), .COUT(n15217));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_1468_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1468_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9_adj_5752[36]), .B1(d9_adj_5751[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15216));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1468_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1468_add_4_1.INIT1 = 16'h9995;
    defparam _add_1_1468_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1468_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_38 (.A0(d_d8[35]), .B0(d8[35]), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15215), 
          .S0(d9_71__N_1675[35]), .S1(cout_adj_5113));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_36 (.A0(d_d8[33]), .B0(d8[33]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[34]), .B1(d8[34]), .C1(GND_net), .D1(VCC_net), .CIN(n15214), 
          .COUT(n15215), .S0(d9_71__N_1675[33]), .S1(d9_71__N_1675[34]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_34 (.A0(d_d8[31]), .B0(d8[31]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[32]), .B1(d8[32]), .C1(GND_net), .D1(VCC_net), .CIN(n15213), 
          .COUT(n15214), .S0(d9_71__N_1675[31]), .S1(d9_71__N_1675[32]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_32 (.A0(d_d8[29]), .B0(d8[29]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[30]), .B1(d8[30]), .C1(GND_net), .D1(VCC_net), .CIN(n15212), 
          .COUT(n15213), .S0(d9_71__N_1675[29]), .S1(d9_71__N_1675[30]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_30 (.A0(d_d8[27]), .B0(d8[27]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[28]), .B1(d8[28]), .C1(GND_net), .D1(VCC_net), .CIN(n15211), 
          .COUT(n15212), .S0(d9_71__N_1675[27]), .S1(d9_71__N_1675[28]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_28 (.A0(d_d8[25]), .B0(d8[25]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[26]), .B1(d8[26]), .C1(GND_net), .D1(VCC_net), .CIN(n15210), 
          .COUT(n15211), .S0(d9_71__N_1675[25]), .S1(d9_71__N_1675[26]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_26 (.A0(d_d8[23]), .B0(d8[23]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[24]), .B1(d8[24]), .C1(GND_net), .D1(VCC_net), .CIN(n15209), 
          .COUT(n15210), .S0(d9_71__N_1675[23]), .S1(d9_71__N_1675[24]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_24 (.A0(d_d8[21]), .B0(d8[21]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[22]), .B1(d8[22]), .C1(GND_net), .D1(VCC_net), .CIN(n15208), 
          .COUT(n15209), .S0(d9_71__N_1675[21]), .S1(d9_71__N_1675[22]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_22 (.A0(d_d8[19]), .B0(d8[19]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[20]), .B1(d8[20]), .C1(GND_net), .D1(VCC_net), .CIN(n15207), 
          .COUT(n15208), .S0(d9_71__N_1675[19]), .S1(d9_71__N_1675[20]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_14 (.A0(d_d8[11]), .B0(d8[11]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[12]), .B1(d8[12]), .C1(GND_net), .D1(VCC_net), .CIN(n15203), 
          .COUT(n15204), .S0(d9_71__N_1675[11]), .S1(d9_71__N_1675[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_20 (.A0(d_d8[17]), .B0(d8[17]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[18]), .B1(d8[18]), .C1(GND_net), .D1(VCC_net), .CIN(n15206), 
          .COUT(n15207), .S0(d9_71__N_1675[17]), .S1(d9_71__N_1675[18]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_10 (.A0(d_d8[7]), .B0(d8[7]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[8]), .B1(d8[8]), .C1(GND_net), .D1(VCC_net), .CIN(n15201), 
          .COUT(n15202), .S0(d9_71__N_1675[7]), .S1(d9_71__N_1675[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_18 (.A0(d_d8[15]), .B0(d8[15]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[16]), .B1(d8[16]), .C1(GND_net), .D1(VCC_net), .CIN(n15205), 
          .COUT(n15206), .S0(d9_71__N_1675[15]), .S1(d9_71__N_1675[16]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_8 (.A0(d_d8[5]), .B0(d8[5]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[6]), .B1(d8[6]), .C1(GND_net), .D1(VCC_net), .CIN(n15200), 
          .COUT(n15201), .S0(d9_71__N_1675[5]), .S1(d9_71__N_1675[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_6 (.A0(d_d8[3]), .B0(d8[3]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[4]), .B1(d8[4]), .C1(GND_net), .D1(VCC_net), .CIN(n15199), 
          .COUT(n15200), .S0(d9_71__N_1675[3]), .S1(d9_71__N_1675[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[0]), .B1(d8[0]), .C1(GND_net), .D1(VCC_net), .COUT(n15198), 
          .S1(d9_71__N_1675[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_12 (.A0(d_d8[9]), .B0(d8[9]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[10]), .B1(d8[10]), .C1(GND_net), .D1(VCC_net), .CIN(n15202), 
          .COUT(n15203), .S0(d9_71__N_1675[9]), .S1(d9_71__N_1675[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_16 (.A0(d_d8[13]), .B0(d8[13]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[14]), .B1(d8[14]), .C1(GND_net), .D1(VCC_net), .CIN(n15204), 
          .COUT(n15205), .S0(d9_71__N_1675[13]), .S1(d9_71__N_1675[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_add_4_16.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_34 (.A0(phase_inc_carrGen1[32]), .B0(phase_accum_adj_5732[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[33]), .B1(phase_accum_adj_5732[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15938), .COUT(n15939), .S0(n225), 
          .S1(n222));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_34.INIT0 = 16'h666a;
    defparam phase_accum_add_4_34.INIT1 = 16'h666a;
    defparam phase_accum_add_4_34.INJECT1_0 = "NO";
    defparam phase_accum_add_4_34.INJECT1_1 = "NO";
    CCU2C add_3830_19 (.A0(d_out_d_11__N_1886[17]), .B0(n48_adj_5536), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), .B1(n45_adj_5535), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16698), .S0(n45_adj_5275), 
          .S1(d_out_d_11__N_1888[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3830_19.INIT0 = 16'h9995;
    defparam add_3830_19.INIT1 = 16'h9995;
    defparam add_3830_19.INJECT1_0 = "NO";
    defparam add_3830_19.INJECT1_1 = "NO";
    CCU2C add_3830_17 (.A0(d_out_d_11__N_1886[17]), .B0(n54_adj_5538), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), .B1(n51_adj_5537), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16697), .COUT(n16698), .S0(n51_adj_5277), 
          .S1(n48_adj_5276));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3830_17.INIT0 = 16'h9995;
    defparam add_3830_17.INIT1 = 16'h9995;
    defparam add_3830_17.INJECT1_0 = "NO";
    defparam add_3830_17.INJECT1_1 = "NO";
    CCU2C add_3830_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1886[17]), .C0(n60_adj_5540), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1886[17]), 
          .C1(n57_adj_5539), .D1(VCC_net), .CIN(n16696), .COUT(n16697), 
          .S0(n57_adj_5279), .S1(n54_adj_5278));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3830_15.INIT0 = 16'h6969;
    defparam add_3830_15.INIT1 = 16'h6969;
    defparam add_3830_15.INJECT1_0 = "NO";
    defparam add_3830_15.INJECT1_1 = "NO";
    CCU2C add_3830_13 (.A0(d_out_d_11__N_1886[17]), .B0(n66_adj_5542), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1886[17]), 
          .C1(n63_adj_5541), .D1(VCC_net), .CIN(n16695), .COUT(n16696), 
          .S0(n63_adj_5281), .S1(n60_adj_5280));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3830_13.INIT0 = 16'h9995;
    defparam add_3830_13.INIT1 = 16'h6969;
    defparam add_3830_13.INJECT1_0 = "NO";
    defparam add_3830_13.INJECT1_1 = "NO";
    CCU2C add_3830_11 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(n72_adj_5544), .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), 
          .B1(n17938), .C1(n69_adj_5543), .D1(VCC_net), .CIN(n16694), 
          .COUT(n16695), .S0(n69), .S1(n66_adj_5282));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3830_11.INIT0 = 16'h9696;
    defparam add_3830_11.INIT1 = 16'h6969;
    defparam add_3830_11.INJECT1_0 = "NO";
    defparam add_3830_11.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_32 (.A0(phase_inc_carrGen1[30]), .B0(phase_accum_adj_5732[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[31]), .B1(phase_accum_adj_5732[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15937), .COUT(n15938), .S0(n231), 
          .S1(n228));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_32.INIT0 = 16'h666a;
    defparam phase_accum_add_4_32.INIT1 = 16'h666a;
    defparam phase_accum_add_4_32.INJECT1_0 = "NO";
    defparam phase_accum_add_4_32.INJECT1_1 = "NO";
    CCU2C add_3830_9 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(n78_adj_5546), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(n75_adj_5545), .D1(VCC_net), 
          .CIN(n16693), .COUT(n16694), .S0(n75), .S1(n72));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3830_9.INIT0 = 16'h9696;
    defparam add_3830_9.INIT1 = 16'h9696;
    defparam add_3830_9.INJECT1_0 = "NO";
    defparam add_3830_9.INJECT1_1 = "NO";
    CCU2C add_3830_7 (.A0(d_out_d_11__N_1882[17]), .B0(d_out_d_11__N_1886[17]), 
          .C0(n84_adj_5548), .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), 
          .B1(d_out_d_11__N_1886[17]), .C1(n81_adj_5547), .D1(VCC_net), 
          .CIN(n16692), .COUT(n16693), .S0(n81_adj_5284), .S1(n78_adj_5283));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3830_7.INIT0 = 16'h9696;
    defparam add_3830_7.INIT1 = 16'h9696;
    defparam add_3830_7.INJECT1_0 = "NO";
    defparam add_3830_7.INJECT1_1 = "NO";
    CCU2C add_3830_5 (.A0(n90_adj_5550), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1884[17]), .B1(d_out_d_11__N_1886[17]), .C1(n87_adj_5549), 
          .D1(VCC_net), .CIN(n16691), .COUT(n16692), .S0(n87_adj_5286), 
          .S1(n84_adj_5285));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3830_5.INIT0 = 16'haaa0;
    defparam add_3830_5.INIT1 = 16'h9696;
    defparam add_3830_5.INJECT1_0 = "NO";
    defparam add_3830_5.INJECT1_1 = "NO";
    CCU2C add_3830_3 (.A0(d_out_d_11__N_1886[17]), .B0(ISquare[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16690), .COUT(n16691), .S1(n90_adj_5287));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3830_3.INIT0 = 16'h666a;
    defparam add_3830_3.INIT1 = 16'h555f;
    defparam add_3830_3.INJECT1_0 = "NO";
    defparam add_3830_3.INJECT1_1 = "NO";
    FD1P3AX phase_inc_carrGen_i0_i2 (.D(n317), .SP(clk_80mhz_enable_1471), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i2.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i3 (.D(n314), .SP(clk_80mhz_enable_1471), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i3.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i4 (.D(n311), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i4.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i5 (.D(n308), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i5.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i6 (.D(n305), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i6.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i7 (.D(n302), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i7.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i8 (.D(n299), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i8.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i9 (.D(n296), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i9.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i10 (.D(n293), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i10.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i11 (.D(n290), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i11.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i12 (.D(n287), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i12.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i13 (.D(n284), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i13.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i14 (.D(n281), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i14.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i15 (.D(n278), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i15.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i16 (.D(n275), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[16]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i16.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i17 (.D(n272), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i17.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i18 (.D(n269), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[18]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i18.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i19 (.D(n266), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i19.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i20 (.D(n263), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[20]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i20.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i21 (.D(n260), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i21.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i22 (.D(n257), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[22]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i22.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i23 (.D(n254), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i23.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i24 (.D(n251), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[24]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i24.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i25 (.D(n248), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i25.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i26 (.D(n245), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[26]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i26.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i27 (.D(n242), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i27.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i28 (.D(n239), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[28]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i28.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i29 (.D(n236), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i29.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i30 (.D(n233), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[30]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i30.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i31 (.D(n230), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i31.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i32 (.D(n227), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[32]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i32.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i33 (.D(n224), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i33.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i34 (.D(n221), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[34]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i34.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i35 (.D(n218), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i35.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i36 (.D(n215), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[36]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i36.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i37 (.D(n212), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i37.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i38 (.D(n209), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[38]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i38.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i39 (.D(n206), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i39.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i40 (.D(n203), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[40]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i40.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i41 (.D(n200), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i41.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i42 (.D(n197), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[42]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i42.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i43 (.D(n194), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i43.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i44 (.D(n191), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[44]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i44.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i45 (.D(n188), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i45.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i46 (.D(n185), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[46]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i46.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i47 (.D(n182), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i47.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i48 (.D(n179), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[48]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i48.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i49 (.D(n176), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i49.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i50 (.D(n173), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[50]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i50.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i51 (.D(n170), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i51.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i52 (.D(n167), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[52]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i52.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i53 (.D(n164), .SP(clk_80mhz_enable_1459), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i53.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i54 (.D(n161), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[54]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i54.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i55 (.D(n158), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i55.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i56 (.D(n155), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[56]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i56.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i57 (.D(n152), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i57.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i58 (.D(n149), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[58]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i58.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i59 (.D(n146), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i59.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i60 (.D(n143), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[60]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i60.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i61 (.D(n140), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i61.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i62 (.D(n137), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[62]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i62.GSR = "ENABLED";
    FD1P3AX phase_inc_carrGen_i0_i63 (.D(n134_adj_5111), .SP(clk_80mhz_enable_1469), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i63.GSR = "ENABLED";
    CCU2C add_3830_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1886[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16690));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3830_1.INIT0 = 16'h0000;
    defparam add_3830_1.INIT1 = 16'haaaf;
    defparam add_3830_1.INJECT1_0 = "NO";
    defparam add_3830_1.INJECT1_1 = "NO";
    CCU2C _add_1_1439_add_4_30 (.A0(d5_adj_5744[28]), .B0(d4_adj_5743[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[29]), .B1(d4_adj_5743[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16113), .COUT(n16114), .S0(d5_71__N_706_adj_5760[28]), 
          .S1(d5_71__N_706_adj_5760[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_30.INJECT1_1 = "NO";
    LUT4 i2326_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(n18076), .D(n217_adj_5660), 
         .Z(n12124)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2326_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_325_i28_4_lut (.A(n12114), .B(n238), .C(n17925), .D(n2572), 
         .Z(n2344)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i28_4_lut.init = 16'hc0ca;
    LUT4 i2328_3_lut_4_lut (.A(n18075), .B(n17937), .C(led_c_3), .D(n214_adj_5659), 
         .Z(n12126)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2328_3_lut_4_lut.init = 16'hfb0b;
    CCU2C add_3831_19 (.A0(d_out_d_11__N_1890[17]), .B0(n48_adj_5589), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1890[17]), .B1(n45_adj_5588), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16684), .S0(n916), .S1(d_out_d_11__N_1892[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3831_19.INIT0 = 16'h9995;
    defparam add_3831_19.INIT1 = 16'h9995;
    defparam add_3831_19.INJECT1_0 = "NO";
    defparam add_3831_19.INJECT1_1 = "NO";
    LUT4 mux_325_i25_4_lut (.A(n12108), .B(n247), .C(n17925), .D(n2572), 
         .Z(n2347)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i25_4_lut.init = 16'hc0ca;
    CCU2C add_3831_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1890[17]), .C0(n54_adj_5591), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1890[17]), 
          .C1(n51_adj_5590), .D1(VCC_net), .CIN(n16683), .COUT(n16684), 
          .S0(n918), .S1(n917));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3831_17.INIT0 = 16'h6969;
    defparam add_3831_17.INIT1 = 16'h6969;
    defparam add_3831_17.INJECT1_0 = "NO";
    defparam add_3831_17.INJECT1_1 = "NO";
    CCU2C add_3831_15 (.A0(d_out_d_11__N_1890[17]), .B0(n60_adj_5593), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1890[17]), 
          .C1(n57_adj_5592), .D1(VCC_net), .CIN(n16682), .COUT(n16683), 
          .S0(n920), .S1(n919));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3831_15.INIT0 = 16'h9995;
    defparam add_3831_15.INIT1 = 16'h6969;
    defparam add_3831_15.INJECT1_0 = "NO";
    defparam add_3831_15.INJECT1_1 = "NO";
    CCU2C add_3831_13 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n66_adj_5595), .D0(VCC_net), .A1(d_out_d_11__N_1890[17]), 
          .B1(n17938), .C1(n63_adj_5594), .D1(VCC_net), .CIN(n16681), 
          .COUT(n16682), .S0(n922), .S1(n921));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3831_13.INIT0 = 16'h9696;
    defparam add_3831_13.INIT1 = 16'h6969;
    defparam add_3831_13.INJECT1_0 = "NO";
    defparam add_3831_13.INJECT1_1 = "NO";
    LUT4 mux_325_i26_4_lut (.A(n12110), .B(n244), .C(n17925), .D(n2572), 
         .Z(n2346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i26_4_lut.init = 16'hcfca;
    LUT4 i2288_3_lut_4_lut (.A(n18075), .B(n17937), .C(led_c_3), .D(n283_adj_5682), 
         .Z(n12086)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2288_3_lut_4_lut.init = 16'hf404;
    LUT4 i2278_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(led_c_3), .D(n301_adj_5688), 
         .Z(n12076)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2278_3_lut_4_lut.init = 16'hf404;
    LUT4 i26_4_lut (.A(n2572), .B(n253), .C(n17925), .D(n13_adj_4794), 
         .Z(n11_adj_4791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i26_4_lut.init = 16'hcacf;
    LUT4 mux_325_i24_4_lut (.A(n12106), .B(n250), .C(n17925), .D(n2572), 
         .Z(n2348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i24_4_lut.init = 16'hcfca;
    LUT4 mux_325_i21_4_lut (.A(n12102), .B(n259), .C(n17925), .D(n2572), 
         .Z(n2351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i21_4_lut.init = 16'hcfca;
    LUT4 i2480_4_lut (.A(n256), .B(n250_adj_5671), .C(led_c_3), .D(n17932), 
         .Z(n12294)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2480_4_lut.init = 16'hcac0;
    LUT4 mux_325_i19_4_lut (.A(n12098), .B(n265), .C(n17925), .D(n2572), 
         .Z(n2353)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i19_4_lut.init = 16'hcfca;
    LUT4 i2478_4_lut (.A(n262), .B(n256_adj_5673), .C(led_c_3), .D(n17932), 
         .Z(n12292)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2478_4_lut.init = 16'hcac0;
    LUT4 mux_325_i17_4_lut (.A(n12094), .B(n271), .C(n17925), .D(n2572), 
         .Z(n2355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i17_4_lut.init = 16'hcfca;
    LUT4 mux_325_i18_4_lut (.A(n2554), .B(n268), .C(n17925), .D(n2572), 
         .Z(n2354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i18_4_lut.init = 16'hcfca;
    LUT4 i2362_3_lut_4_lut (.A(n18075), .B(n17937), .C(n18076), .D(n154_adj_5639), 
         .Z(n12160)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2362_3_lut_4_lut.init = 16'hf707;
    LUT4 i3287_2_lut (.A(n262_adj_5675), .B(n18076), .Z(n2554)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i3287_2_lut.init = 16'h8888;
    CCU2C add_3831_11 (.A0(d_out_d_11__N_1878[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n72_adj_5597), .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(n69_adj_5596), .D1(VCC_net), 
          .CIN(n16680), .COUT(n16681), .S0(n924), .S1(n923));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3831_11.INIT0 = 16'h9696;
    defparam add_3831_11.INIT1 = 16'h9696;
    defparam add_3831_11.INJECT1_0 = "NO";
    defparam add_3831_11.INJECT1_1 = "NO";
    LUT4 mux_325_i15_4_lut (.A(n12092), .B(n277), .C(n17925), .D(n2572), 
         .Z(n2357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i15_4_lut.init = 16'hcfca;
    LUT4 i2310_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(led_c_3), .D(n241_adj_5668), 
         .Z(n12108)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2310_3_lut_4_lut.init = 16'hfb0b;
    CCU2C add_3831_9 (.A0(d_out_d_11__N_1882[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n78_adj_5599), .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(n75_adj_5598), .D1(VCC_net), 
          .CIN(n16679), .COUT(n16680), .S0(n926), .S1(n925));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3831_9.INIT0 = 16'h9696;
    defparam add_3831_9.INIT1 = 16'h9696;
    defparam add_3831_9.INJECT1_0 = "NO";
    defparam add_3831_9.INJECT1_1 = "NO";
    LUT4 i2300_3_lut_4_lut (.A(n18075), .B(n17937), .C(led_c_3), .D(n259_adj_5674), 
         .Z(n12098)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2300_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i3089_4_lut (.A(n27_adj_5727), .B(n274), .C(n17925), .D(n2422), 
         .Z(n2356)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i3089_4_lut.init = 16'hc5c0;
    CCU2C add_3831_7 (.A0(d_out_d_11__N_1886[17]), .B0(d_out_d_11__N_1890[17]), 
          .C0(n84_adj_5601), .D0(VCC_net), .A1(d_out_d_11__N_1884[17]), 
          .B1(d_out_d_11__N_1890[17]), .C1(n81_adj_5600), .D1(VCC_net), 
          .CIN(n16678), .COUT(n16679), .S0(n928), .S1(n927));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3831_7.INIT0 = 16'h9696;
    defparam add_3831_7.INIT1 = 16'h9696;
    defparam add_3831_7.INJECT1_0 = "NO";
    defparam add_3831_7.INJECT1_1 = "NO";
    LUT4 i3081_4_lut (.A(n27_adj_5727), .B(n283), .C(n17925), .D(n2425), 
         .Z(n2359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i3081_4_lut.init = 16'hcfca;
    CCU2C add_3831_5 (.A0(n90_adj_5603), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1888[17]), .B1(d_out_d_11__N_1890[17]), .C1(n87_adj_5602), 
          .D1(VCC_net), .CIN(n16677), .COUT(n16678), .S0(n930), .S1(n929));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3831_5.INIT0 = 16'haaa0;
    defparam add_3831_5.INIT1 = 16'h9696;
    defparam add_3831_5.INJECT1_0 = "NO";
    defparam add_3831_5.INJECT1_1 = "NO";
    LUT4 i3227_2_lut (.A(n277_adj_5680), .B(n18076), .Z(n2425)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i3227_2_lut.init = 16'h8888;
    CCU2C add_3831_3 (.A0(d_out_d_11__N_1890[17]), .B0(ISquare[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16676), .COUT(n16677), .S1(n931));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3831_3.INIT0 = 16'h666a;
    defparam add_3831_3.INIT1 = 16'h555f;
    defparam add_3831_3.INJECT1_0 = "NO";
    defparam add_3831_3.INJECT1_1 = "NO";
    LUT4 mux_325_i14_4_lut (.A(n2558), .B(n280), .C(n17925), .D(n2572), 
         .Z(n2358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i14_4_lut.init = 16'hcfca;
    CCU2C add_3831_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1890[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16676));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3831_1.INIT0 = 16'h0000;
    defparam add_3831_1.INIT1 = 16'haaaf;
    defparam add_3831_1.INJECT1_0 = "NO";
    defparam add_3831_1.INJECT1_1 = "NO";
    LUT4 i3286_2_lut (.A(n274_adj_5679), .B(led_c_3), .Z(n2558)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i3286_2_lut.init = 16'h8888;
    CCU2C add_3832_17 (.A0(d_out_d_11__N_1877), .B0(d_out_d_11__N_1878[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1877), .B1(d_out_d_11__N_1878[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16670), .S0(n41), .S1(d_out_d_11__N_1880[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3832_17.INIT0 = 16'h666a;
    defparam add_3832_17.INIT1 = 16'h666a;
    defparam add_3832_17.INJECT1_0 = "NO";
    defparam add_3832_17.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_15 (.A0(d1_adj_5740[48]), .B0(cout_adj_5344), 
          .C0(n147), .D0(d2_adj_5741[48]), .A1(d1_adj_5740[49]), .B1(cout_adj_5344), 
          .C1(n144), .D1(d2_adj_5741[49]), .CIN(n16493), .COUT(n16494), 
          .S0(d2_71__N_490_adj_5757[48]), .S1(d2_71__N_490_adj_5757[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_15.INJECT1_1 = "NO";
    CCU2C add_3832_15 (.A0(d_out_d_11__N_1878[17]), .B0(n40), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n37_adj_5614), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16669), .COUT(n16670), .S0(n47), 
          .S1(n44));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3832_15.INIT0 = 16'h9995;
    defparam add_3832_15.INIT1 = 16'h9995;
    defparam add_3832_15.INJECT1_0 = "NO";
    defparam add_3832_15.INJECT1_1 = "NO";
    CCU2C add_3832_13 (.A0(d_out_d_11__N_1878[17]), .B0(n46), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n43), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16668), .COUT(n16669), .S0(n53), .S1(n50));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3832_13.INIT0 = 16'h9995;
    defparam add_3832_13.INIT1 = 16'h9995;
    defparam add_3832_13.INJECT1_0 = "NO";
    defparam add_3832_13.INJECT1_1 = "NO";
    CCU2C add_3832_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1878[17]), .C0(n52), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1878[17]), 
          .C1(n49), .D1(VCC_net), .CIN(n16667), .COUT(n16668), .S0(n59), 
          .S1(n56));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3832_11.INIT0 = 16'h6969;
    defparam add_3832_11.INIT1 = 16'h6969;
    defparam add_3832_11.INJECT1_0 = "NO";
    defparam add_3832_11.INJECT1_1 = "NO";
    CCU2C add_3832_9 (.A0(d_out_d_11__N_1878[17]), .B0(n58), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1878[17]), 
          .C1(n55), .D1(VCC_net), .CIN(n16666), .COUT(n16667), .S0(n65_adj_5604), 
          .S1(n62));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3832_9.INIT0 = 16'h9995;
    defparam add_3832_9.INIT1 = 16'h6969;
    defparam add_3832_9.INJECT1_0 = "NO";
    defparam add_3832_9.INJECT1_1 = "NO";
    CCU2C add_3832_7 (.A0(d_out_d_11__N_1874[17]), .B0(d_out_d_11__N_1878[17]), 
          .C0(n64_adj_5615), .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(n17938), .C1(n61), .D1(VCC_net), .CIN(n16665), .COUT(n16666), 
          .S0(n71), .S1(n68));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3832_7.INIT0 = 16'h9696;
    defparam add_3832_7.INIT1 = 16'h6969;
    defparam add_3832_7.INJECT1_0 = "NO";
    defparam add_3832_7.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_13 (.A0(d1_adj_5740[46]), .B0(cout_adj_5344), 
          .C0(n153), .D0(d2_adj_5741[46]), .A1(d1_adj_5740[47]), .B1(cout_adj_5344), 
          .C1(n150), .D1(d2_adj_5741[47]), .CIN(n16492), .COUT(n16493), 
          .S0(d2_71__N_490_adj_5757[46]), .S1(d2_71__N_490_adj_5757[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_13.INJECT1_1 = "NO";
    CCU2C add_3832_5 (.A0(n70), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1876[17]), .B1(d_out_d_11__N_1878[17]), .C1(n67), 
          .D1(VCC_net), .CIN(n16664), .COUT(n16665), .S0(n77), .S1(n74));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3832_5.INIT0 = 16'haaa0;
    defparam add_3832_5.INIT1 = 16'h9696;
    defparam add_3832_5.INJECT1_0 = "NO";
    defparam add_3832_5.INJECT1_1 = "NO";
    CCU2C add_3832_3 (.A0(d_out_d_11__N_1878[17]), .B0(ISquare[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16663), .COUT(n16664), .S1(n80));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3832_3.INIT0 = 16'h666a;
    defparam add_3832_3.INIT1 = 16'h555f;
    defparam add_3832_3.INJECT1_0 = "NO";
    defparam add_3832_3.INJECT1_1 = "NO";
    CCU2C add_3832_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1878[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16663));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3832_1.INIT0 = 16'h0000;
    defparam add_3832_1.INIT1 = 16'haaaf;
    defparam add_3832_1.INJECT1_0 = "NO";
    defparam add_3832_1.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_11 (.A0(d1_adj_5740[44]), .B0(cout_adj_5344), 
          .C0(n159), .D0(d2_adj_5741[44]), .A1(d1_adj_5740[45]), .B1(cout_adj_5344), 
          .C1(n156), .D1(d2_adj_5741[45]), .CIN(n16491), .COUT(n16492), 
          .S0(d2_71__N_490_adj_5757[44]), .S1(d2_71__N_490_adj_5757[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_11.INJECT1_1 = "NO";
    CCU2C add_3833_19 (.A0(d_out_d_11__N_1888[17]), .B0(n48_adj_5276), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n45_adj_5275), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16657), .S0(n45_adj_5588), 
          .S1(d_out_d_11__N_1890[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3833_19.INIT0 = 16'h9995;
    defparam add_3833_19.INIT1 = 16'h9995;
    defparam add_3833_19.INJECT1_0 = "NO";
    defparam add_3833_19.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_9 (.A0(d1_adj_5740[42]), .B0(cout_adj_5344), 
          .C0(n165), .D0(d2_adj_5741[42]), .A1(d1_adj_5740[43]), .B1(cout_adj_5344), 
          .C1(n162), .D1(d2_adj_5741[43]), .CIN(n16490), .COUT(n16491), 
          .S0(d2_71__N_490_adj_5757[42]), .S1(d2_71__N_490_adj_5757[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_9.INJECT1_1 = "NO";
    CCU2C add_3833_17 (.A0(ISquare[31]), .B0(d_out_d_11__N_1888[17]), .C0(n54_adj_5278), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n51_adj_5277), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16656), .COUT(n16657), .S0(n51_adj_5590), 
          .S1(n48_adj_5589));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3833_17.INIT0 = 16'h6969;
    defparam add_3833_17.INIT1 = 16'h9995;
    defparam add_3833_17.INJECT1_0 = "NO";
    defparam add_3833_17.INJECT1_1 = "NO";
    CCU2C add_3833_15 (.A0(ISquare[31]), .B0(d_out_d_11__N_1888[17]), .C0(n60_adj_5280), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1888[17]), 
          .C1(n57_adj_5279), .D1(VCC_net), .CIN(n16655), .COUT(n16656), 
          .S0(n57_adj_5592), .S1(n54_adj_5591));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3833_15.INIT0 = 16'h6969;
    defparam add_3833_15.INIT1 = 16'h6969;
    defparam add_3833_15.INJECT1_0 = "NO";
    defparam add_3833_15.INJECT1_1 = "NO";
    CCU2C add_3833_13 (.A0(d_out_d_11__N_1888[17]), .B0(n17938), .C0(n66_adj_5282), 
          .D0(VCC_net), .A1(d_out_d_11__N_1888[17]), .B1(n63_adj_5281), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16654), .COUT(n16655), .S0(n63_adj_5594), 
          .S1(n60_adj_5593));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3833_13.INIT0 = 16'h6969;
    defparam add_3833_13.INIT1 = 16'h9995;
    defparam add_3833_13.INJECT1_0 = "NO";
    defparam add_3833_13.INJECT1_1 = "NO";
    CCU2C add_3833_11 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(n72), .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), .B1(d_out_d_11__N_1888[17]), 
          .C1(n69), .D1(VCC_net), .CIN(n16653), .COUT(n16654), .S0(n69_adj_5596), 
          .S1(n66_adj_5595));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3833_11.INIT0 = 16'h9696;
    defparam add_3833_11.INIT1 = 16'h9696;
    defparam add_3833_11.INJECT1_0 = "NO";
    defparam add_3833_11.INJECT1_1 = "NO";
    CCU2C add_3833_9 (.A0(d_out_d_11__N_1880[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(n78_adj_5283), .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(n75), .D1(VCC_net), .CIN(n16652), 
          .COUT(n16653), .S0(n75_adj_5598), .S1(n72_adj_5597));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3833_9.INIT0 = 16'h9696;
    defparam add_3833_9.INIT1 = 16'h9696;
    defparam add_3833_9.INJECT1_0 = "NO";
    defparam add_3833_9.INJECT1_1 = "NO";
    CCU2C add_3833_7 (.A0(d_out_d_11__N_1884[17]), .B0(d_out_d_11__N_1888[17]), 
          .C0(n84_adj_5285), .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), 
          .B1(d_out_d_11__N_1888[17]), .C1(n81_adj_5284), .D1(VCC_net), 
          .CIN(n16651), .COUT(n16652), .S0(n81_adj_5600), .S1(n78_adj_5599));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3833_7.INIT0 = 16'h9696;
    defparam add_3833_7.INIT1 = 16'h9696;
    defparam add_3833_7.INJECT1_0 = "NO";
    defparam add_3833_7.INJECT1_1 = "NO";
    CCU2C add_3833_5 (.A0(n90_adj_5287), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1886[17]), .B1(d_out_d_11__N_1888[17]), .C1(n87_adj_5286), 
          .D1(VCC_net), .CIN(n16650), .COUT(n16651), .S0(n87_adj_5602), 
          .S1(n84_adj_5601));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3833_5.INIT0 = 16'haaa0;
    defparam add_3833_5.INIT1 = 16'h9696;
    defparam add_3833_5.INJECT1_0 = "NO";
    defparam add_3833_5.INJECT1_1 = "NO";
    CCU2C add_3833_3 (.A0(d_out_d_11__N_1888[17]), .B0(ISquare[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16649), .COUT(n16650), .S1(n90_adj_5603));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3833_3.INIT0 = 16'h666a;
    defparam add_3833_3.INIT1 = 16'h555f;
    defparam add_3833_3.INJECT1_0 = "NO";
    defparam add_3833_3.INJECT1_1 = "NO";
    CCU2C add_3833_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1888[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16649));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3833_1.INIT0 = 16'h0000;
    defparam add_3833_1.INIT1 = 16'haaaf;
    defparam add_3833_1.INJECT1_0 = "NO";
    defparam add_3833_1.INJECT1_1 = "NO";
    CCU2C add_3828_65 (.A0(phase_inc_carrGen[62]), .B0(n17926), .C0(n12304), 
          .D0(n3660), .A1(phase_inc_carrGen[63]), .B1(n17926), .C1(n12306), 
          .D1(n3660), .CIN(n16643), .S0(n137), .S1(n134_adj_5111));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_65.INIT0 = 16'h74b8;
    defparam add_3828_65.INIT1 = 16'h74b8;
    defparam add_3828_65.INJECT1_0 = "NO";
    defparam add_3828_65.INJECT1_1 = "NO";
    CCU2C add_3828_63 (.A0(phase_inc_carrGen[60]), .B0(n17926), .C0(n2311), 
          .D0(n3660), .A1(phase_inc_carrGen[61]), .B1(n17926), .C1(n12302), 
          .D1(n3660), .CIN(n16642), .COUT(n16643), .S0(n143), .S1(n140));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_63.INIT0 = 16'h74b8;
    defparam add_3828_63.INIT1 = 16'h74b8;
    defparam add_3828_63.INJECT1_0 = "NO";
    defparam add_3828_63.INJECT1_1 = "NO";
    CCU2C add_3828_61 (.A0(phase_inc_carrGen[58]), .B0(n17926), .C0(n2313), 
          .D0(n3660), .A1(phase_inc_carrGen[59]), .B1(n17926), .C1(n2312), 
          .D1(n3660), .CIN(n16641), .COUT(n16642), .S0(n149), .S1(n146));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_61.INIT0 = 16'h74b8;
    defparam add_3828_61.INIT1 = 16'h74b8;
    defparam add_3828_61.INJECT1_0 = "NO";
    defparam add_3828_61.INJECT1_1 = "NO";
    CCU2C add_3828_59 (.A0(phase_inc_carrGen[56]), .B0(n17926), .C0(n2315), 
          .D0(n3660), .A1(phase_inc_carrGen[57]), .B1(n17926), .C1(n12300), 
          .D1(n3660), .CIN(n16640), .COUT(n16641), .S0(n155), .S1(n152));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_59.INIT0 = 16'h74b8;
    defparam add_3828_59.INIT1 = 16'h74b8;
    defparam add_3828_59.INJECT1_0 = "NO";
    defparam add_3828_59.INJECT1_1 = "NO";
    CCU2C add_3828_57 (.A0(phase_inc_carrGen[54]), .B0(n17926), .C0(n2317), 
          .D0(n3660), .A1(phase_inc_carrGen[55]), .B1(n17926), .C1(n21_adj_5729), 
          .D1(n3660), .CIN(n16639), .COUT(n16640), .S0(n161), .S1(n158));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_57.INIT0 = 16'h74b8;
    defparam add_3828_57.INIT1 = 16'h74b8;
    defparam add_3828_57.INJECT1_0 = "NO";
    defparam add_3828_57.INJECT1_1 = "NO";
    CCU2C add_3828_55 (.A0(phase_inc_carrGen[52]), .B0(n17926), .C0(n12298), 
          .D0(n3660), .A1(phase_inc_carrGen[53]), .B1(n17926), .C1(n2318), 
          .D1(n3660), .CIN(n16638), .COUT(n16639), .S0(n167), .S1(n164));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_55.INIT0 = 16'h74b8;
    defparam add_3828_55.INIT1 = 16'h74b8;
    defparam add_3828_55.INJECT1_0 = "NO";
    defparam add_3828_55.INJECT1_1 = "NO";
    CCU2C add_3828_53 (.A0(phase_inc_carrGen[50]), .B0(n17926), .C0(n2321), 
          .D0(n3657), .A1(phase_inc_carrGen[51]), .B1(n17926), .C1(n2320), 
          .D1(n3660), .CIN(n16637), .COUT(n16638), .S0(n173), .S1(n170));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_53.INIT0 = 16'h74b8;
    defparam add_3828_53.INIT1 = 16'h74b8;
    defparam add_3828_53.INJECT1_0 = "NO";
    defparam add_3828_53.INJECT1_1 = "NO";
    CCU2C add_3828_51 (.A0(phase_inc_carrGen[48]), .B0(n17926), .C0(n2323), 
          .D0(n3657), .A1(phase_inc_carrGen[49]), .B1(n17926), .C1(n2322), 
          .D1(n3657), .CIN(n16636), .COUT(n16637), .S0(n179), .S1(n176));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_51.INIT0 = 16'h74b8;
    defparam add_3828_51.INIT1 = 16'h74b8;
    defparam add_3828_51.INJECT1_0 = "NO";
    defparam add_3828_51.INJECT1_1 = "NO";
    CCU2C add_3828_49 (.A0(phase_inc_carrGen[46]), .B0(n17926), .C0(n2325), 
          .D0(n11804), .A1(phase_inc_carrGen[47]), .B1(n17926), .C1(n2324), 
          .D1(n11804), .CIN(n16635), .COUT(n16636), .S0(n185), .S1(n182));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_49.INIT0 = 16'h74b8;
    defparam add_3828_49.INIT1 = 16'h74b8;
    defparam add_3828_49.INJECT1_0 = "NO";
    defparam add_3828_49.INJECT1_1 = "NO";
    CCU2C add_3828_47 (.A0(phase_inc_carrGen[44]), .B0(n17926), .C0(n2327), 
          .D0(n17930), .A1(phase_inc_carrGen[45]), .B1(n17926), .C1(n2326), 
          .D1(n3660), .CIN(n16634), .COUT(n16635), .S0(n191), .S1(n188));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_47.INIT0 = 16'h74b8;
    defparam add_3828_47.INIT1 = 16'h74b8;
    defparam add_3828_47.INJECT1_0 = "NO";
    defparam add_3828_47.INJECT1_1 = "NO";
    CCU2C add_3828_45 (.A0(phase_inc_carrGen[42]), .B0(n17926), .C0(n2329), 
          .D0(n17929), .A1(phase_inc_carrGen[43]), .B1(n17926), .C1(n2328), 
          .D1(n3677), .CIN(n16633), .COUT(n16634), .S0(n197), .S1(n194));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_45.INIT0 = 16'h74b8;
    defparam add_3828_45.INIT1 = 16'h74b8;
    defparam add_3828_45.INJECT1_0 = "NO";
    defparam add_3828_45.INJECT1_1 = "NO";
    CCU2C add_3828_43 (.A0(phase_inc_carrGen[40]), .B0(n17926), .C0(n11_adj_5725), 
          .D0(n3657), .A1(phase_inc_carrGen[41]), .B1(n17926), .C1(n12296), 
          .D1(n3677), .CIN(n16632), .COUT(n16633), .S0(n203), .S1(n200));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_43.INIT0 = 16'h74b8;
    defparam add_3828_43.INIT1 = 16'h74b8;
    defparam add_3828_43.INJECT1_0 = "NO";
    defparam add_3828_43.INJECT1_1 = "NO";
    CCU2C add_3828_41 (.A0(phase_inc_carrGen[38]), .B0(n17926), .C0(n2333), 
          .D0(n3660), .A1(phase_inc_carrGen[39]), .B1(n17926), .C1(n2332), 
          .D1(n3660), .CIN(n16631), .COUT(n16632), .S0(n209), .S1(n206));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_41.INIT0 = 16'h74b8;
    defparam add_3828_41.INIT1 = 16'h74b8;
    defparam add_3828_41.INJECT1_0 = "NO";
    defparam add_3828_41.INJECT1_1 = "NO";
    CCU2C add_3828_39 (.A0(phase_inc_carrGen[36]), .B0(n17926), .C0(n2335), 
          .D0(n17930), .A1(phase_inc_carrGen[37]), .B1(n17926), .C1(n2334), 
          .D1(n3678), .CIN(n16630), .COUT(n16631), .S0(n215), .S1(n212));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_39.INIT0 = 16'h74b8;
    defparam add_3828_39.INIT1 = 16'h74b8;
    defparam add_3828_39.INJECT1_0 = "NO";
    defparam add_3828_39.INJECT1_1 = "NO";
    CCU2C add_3828_37 (.A0(phase_inc_carrGen[34]), .B0(n17926), .C0(n2337), 
          .D0(n17930), .A1(phase_inc_carrGen[35]), .B1(n17926), .C1(n2336), 
          .D1(n3660), .CIN(n16629), .COUT(n16630), .S0(n221), .S1(n218));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_37.INIT0 = 16'h74b8;
    defparam add_3828_37.INIT1 = 16'h74b8;
    defparam add_3828_37.INJECT1_0 = "NO";
    defparam add_3828_37.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_7 (.A0(d1_adj_5740[40]), .B0(cout_adj_5344), 
          .C0(n171), .D0(d2_adj_5741[40]), .A1(d1_adj_5740[41]), .B1(cout_adj_5344), 
          .C1(n168), .D1(d2_adj_5741[41]), .CIN(n16489), .COUT(n16490), 
          .S0(d2_71__N_490_adj_5757[40]), .S1(d2_71__N_490_adj_5757[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_7.INJECT1_1 = "NO";
    CCU2C add_3828_35 (.A0(phase_inc_carrGen[32]), .B0(n17926), .C0(n2339), 
          .D0(n3657), .A1(phase_inc_carrGen[33]), .B1(n17926), .C1(n2338), 
          .D1(n3678), .CIN(n16628), .COUT(n16629), .S0(n227), .S1(n224));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_35.INIT0 = 16'h74b8;
    defparam add_3828_35.INIT1 = 16'h74b8;
    defparam add_3828_35.INJECT1_0 = "NO";
    defparam add_3828_35.INJECT1_1 = "NO";
    CCU2C add_3828_33 (.A0(phase_inc_carrGen[30]), .B0(n17926), .C0(n2341), 
          .D0(n3657), .A1(phase_inc_carrGen[31]), .B1(n17926), .C1(n2340), 
          .D1(n3692), .CIN(n16627), .COUT(n16628), .S0(n233), .S1(n230));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_33.INIT0 = 16'h74b8;
    defparam add_3828_33.INIT1 = 16'h74b8;
    defparam add_3828_33.INJECT1_0 = "NO";
    defparam add_3828_33.INJECT1_1 = "NO";
    CCU2C add_3828_31 (.A0(phase_inc_carrGen[28]), .B0(n17926), .C0(n2343), 
          .D0(n3677), .A1(phase_inc_carrGen[29]), .B1(n17926), .C1(n2342), 
          .D1(n17929), .CIN(n16626), .COUT(n16627), .S0(n239), .S1(n236));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_31.INIT0 = 16'h74b8;
    defparam add_3828_31.INIT1 = 16'h74b8;
    defparam add_3828_31.INJECT1_0 = "NO";
    defparam add_3828_31.INJECT1_1 = "NO";
    CCU2C add_3828_29 (.A0(phase_inc_carrGen[26]), .B0(n17926), .C0(n2345), 
          .D0(n3660), .A1(phase_inc_carrGen[27]), .B1(n17926), .C1(n2344), 
          .D1(n3678), .CIN(n16625), .COUT(n16626), .S0(n245), .S1(n242));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_29.INIT0 = 16'h74b8;
    defparam add_3828_29.INIT1 = 16'h74b8;
    defparam add_3828_29.INJECT1_0 = "NO";
    defparam add_3828_29.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_5 (.A0(d1_adj_5740[38]), .B0(cout_adj_5344), 
          .C0(n177), .D0(d2_adj_5741[38]), .A1(d1_adj_5740[39]), .B1(cout_adj_5344), 
          .C1(n174), .D1(d2_adj_5741[39]), .CIN(n16488), .COUT(n16489), 
          .S0(d2_71__N_490_adj_5757[38]), .S1(d2_71__N_490_adj_5757[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_5.INJECT1_1 = "NO";
    CCU2C add_3828_27 (.A0(phase_inc_carrGen[24]), .B0(n17926), .C0(n2347), 
          .D0(n3660), .A1(phase_inc_carrGen[25]), .B1(n17926), .C1(n2346), 
          .D1(n3660), .CIN(n16624), .COUT(n16625), .S0(n251), .S1(n248));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_27.INIT0 = 16'h74b8;
    defparam add_3828_27.INIT1 = 16'h74b8;
    defparam add_3828_27.INJECT1_0 = "NO";
    defparam add_3828_27.INJECT1_1 = "NO";
    CCU2C add_3828_25 (.A0(phase_inc_carrGen[22]), .B0(n17926), .C0(n11_adj_4791), 
          .D0(n17930), .A1(phase_inc_carrGen[23]), .B1(n17926), .C1(n2348), 
          .D1(n17929), .CIN(n16623), .COUT(n16624), .S0(n257), .S1(n254));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_25.INIT0 = 16'h74b8;
    defparam add_3828_25.INIT1 = 16'h74b8;
    defparam add_3828_25.INJECT1_0 = "NO";
    defparam add_3828_25.INJECT1_1 = "NO";
    CCU2C add_3828_23 (.A0(phase_inc_carrGen[20]), .B0(n17926), .C0(n2351), 
          .D0(n3660), .A1(phase_inc_carrGen[21]), .B1(n17926), .C1(n12294), 
          .D1(n3657), .CIN(n16622), .COUT(n16623), .S0(n263), .S1(n260));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_23.INIT0 = 16'h74b8;
    defparam add_3828_23.INIT1 = 16'h74b8;
    defparam add_3828_23.INJECT1_0 = "NO";
    defparam add_3828_23.INJECT1_1 = "NO";
    CCU2C add_3828_21 (.A0(phase_inc_carrGen[18]), .B0(n17926), .C0(n2353), 
          .D0(n17929), .A1(phase_inc_carrGen[19]), .B1(n17926), .C1(n12292), 
          .D1(n3678), .CIN(n16621), .COUT(n16622), .S0(n269), .S1(n266));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_21.INIT0 = 16'h74b8;
    defparam add_3828_21.INIT1 = 16'h74b8;
    defparam add_3828_21.INJECT1_0 = "NO";
    defparam add_3828_21.INJECT1_1 = "NO";
    CCU2C add_3828_19 (.A0(phase_inc_carrGen[16]), .B0(n17926), .C0(n2355), 
          .D0(n3692), .A1(phase_inc_carrGen[17]), .B1(n17926), .C1(n2354), 
          .D1(n11804), .CIN(n16620), .COUT(n16621), .S0(n275), .S1(n272));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_19.INIT0 = 16'h74b8;
    defparam add_3828_19.INIT1 = 16'h74b8;
    defparam add_3828_19.INJECT1_0 = "NO";
    defparam add_3828_19.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_3 (.A0(d1_adj_5740[36]), .B0(cout_adj_5344), 
          .C0(n183), .D0(d2_adj_5741[36]), .A1(d1_adj_5740[37]), .B1(cout_adj_5344), 
          .C1(n180), .D1(d2_adj_5741[37]), .CIN(n16487), .COUT(n16488), 
          .S0(d2_71__N_490_adj_5757[36]), .S1(d2_71__N_490_adj_5757[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1501_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1501_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_3.INJECT1_1 = "NO";
    CCU2C add_3828_17 (.A0(phase_inc_carrGen[14]), .B0(n17926), .C0(n2357), 
          .D0(n17930), .A1(phase_inc_carrGen[15]), .B1(n17926), .C1(n2356), 
          .D1(n3678), .CIN(n16619), .COUT(n16620), .S0(n281), .S1(n278));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_17.INIT0 = 16'h74b8;
    defparam add_3828_17.INIT1 = 16'h74b8;
    defparam add_3828_17.INJECT1_0 = "NO";
    defparam add_3828_17.INJECT1_1 = "NO";
    CCU2C add_3828_15 (.A0(phase_inc_carrGen[12]), .B0(n17926), .C0(n2359), 
          .D0(n17930), .A1(phase_inc_carrGen[13]), .B1(n17926), .C1(n2358), 
          .D1(n3692), .CIN(n16618), .COUT(n16619), .S0(n287), .S1(n284));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_15.INIT0 = 16'h74b8;
    defparam add_3828_15.INIT1 = 16'h74b8;
    defparam add_3828_15.INJECT1_0 = "NO";
    defparam add_3828_15.INJECT1_1 = "NO";
    CCU2C add_3828_13 (.A0(phase_inc_carrGen[10]), .B0(n17926), .C0(n2361), 
          .D0(n3692), .A1(phase_inc_carrGen[11]), .B1(n17926), .C1(n12290), 
          .D1(n3660), .CIN(n16617), .COUT(n16618), .S0(n293), .S1(n290));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_13.INIT0 = 16'h74b8;
    defparam add_3828_13.INIT1 = 16'h74b8;
    defparam add_3828_13.INJECT1_0 = "NO";
    defparam add_3828_13.INJECT1_1 = "NO";
    CCU2C add_3828_11 (.A0(phase_inc_carrGen[8]), .B0(n17926), .C0(n2363), 
          .D0(n3677), .A1(phase_inc_carrGen[9]), .B1(n17926), .C1(n2362), 
          .D1(n17929), .CIN(n16616), .COUT(n16617), .S0(n299), .S1(n296));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_11.INIT0 = 16'h74b8;
    defparam add_3828_11.INIT1 = 16'h74b8;
    defparam add_3828_11.INJECT1_0 = "NO";
    defparam add_3828_11.INJECT1_1 = "NO";
    CCU2C add_3828_9 (.A0(phase_inc_carrGen[6]), .B0(n17926), .C0(n2365), 
          .D0(n3678), .A1(phase_inc_carrGen[7]), .B1(n17926), .C1(n2364), 
          .D1(n17929), .CIN(n16615), .COUT(n16616), .S0(n305), .S1(n302));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_9.INIT0 = 16'h74b8;
    defparam add_3828_9.INIT1 = 16'h74b8;
    defparam add_3828_9.INJECT1_0 = "NO";
    defparam add_3828_9.INJECT1_1 = "NO";
    CCU2C add_3828_7 (.A0(phase_inc_carrGen[4]), .B0(n17926), .C0(n2367), 
          .D0(n3678), .A1(phase_inc_carrGen[5]), .B1(n17926), .C1(n2366), 
          .D1(n3678), .CIN(n16614), .COUT(n16615), .S0(n311), .S1(n308));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_7.INIT0 = 16'h74b8;
    defparam add_3828_7.INIT1 = 16'h74b8;
    defparam add_3828_7.INJECT1_0 = "NO";
    defparam add_3828_7.INJECT1_1 = "NO";
    CCU2C add_3828_5 (.A0(phase_inc_carrGen[2]), .B0(n17926), .C0(n17955), 
          .D0(n11804), .A1(phase_inc_carrGen[3]), .B1(n17926), .C1(n17961), 
          .D1(n11804), .CIN(n16613), .COUT(n16614), .S0(n317), .S1(n314));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_5.INIT0 = 16'h74b8;
    defparam add_3828_5.INIT1 = 16'h74b8;
    defparam add_3828_5.INJECT1_0 = "NO";
    defparam add_3828_5.INJECT1_1 = "NO";
    CCU2C add_3828_3 (.A0(phase_inc_carrGen[0]), .B0(n17926), .C0(n16718), 
          .D0(n17929), .A1(phase_inc_carrGen[1]), .B1(n17926), .C1(n17954), 
          .D1(n3692), .CIN(n16612), .COUT(n16613), .S0(n323), .S1(n320));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_3.INIT0 = 16'h74b8;
    defparam add_3828_3.INIT1 = 16'h74b8;
    defparam add_3828_3.INJECT1_0 = "NO";
    defparam add_3828_3.INJECT1_1 = "NO";
    CCU2C _add_1_1501_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5344), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16487));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(63[15:24])
    defparam _add_1_1501_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1501_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1501_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1501_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_37 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n81_adj_2859), .D0(d1_adj_5740[70]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n78_adj_2860), .D1(d1_adj_5740[71]), 
          .CIN(n16482), .S0(d1_71__N_418_adj_5756[70]), .S1(d1_71__N_418_adj_5756[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_35 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n87_adj_2857), .D0(d1_adj_5740[68]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n84_adj_2858), .D1(d1_adj_5740[69]), 
          .CIN(n16481), .COUT(n16482), .S0(d1_71__N_418_adj_5756[68]), 
          .S1(d1_71__N_418_adj_5756[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_35.INJECT1_1 = "NO";
    LUT4 i5368_2_lut (.A(phase_inc_carrGen1[0]), .B(phase_accum_adj_5732[0]), 
         .Z(n321)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5368_2_lut.init = 16'h6666;
    CCU2C _add_1_1504_add_4_33 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n93_adj_2855), .D0(d1_adj_5740[66]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n90_adj_2856), .D1(d1_adj_5740[67]), 
          .CIN(n16480), .COUT(n16481), .S0(d1_71__N_418_adj_5756[66]), 
          .S1(d1_71__N_418_adj_5756[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_31 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n99_adj_2853), .D0(d1_adj_5740[64]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n96_adj_2854), .D1(d1_adj_5740[65]), 
          .CIN(n16479), .COUT(n16480), .S0(d1_71__N_418_adj_5756[64]), 
          .S1(d1_71__N_418_adj_5756[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_29 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n105_adj_2851), .D0(d1_adj_5740[62]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n102_adj_2852), .D1(d1_adj_5740[63]), 
          .CIN(n16478), .COUT(n16479), .S0(d1_71__N_418_adj_5756[62]), 
          .S1(d1_71__N_418_adj_5756[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_27 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n111_adj_2849), .D0(d1_adj_5740[60]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n108_adj_2850), .D1(d1_adj_5740[61]), 
          .CIN(n16477), .COUT(n16478), .S0(d1_71__N_418_adj_5756[60]), 
          .S1(d1_71__N_418_adj_5756[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_25 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n117_adj_2847), .D0(d1_adj_5740[58]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n114_adj_2848), .D1(d1_adj_5740[59]), 
          .CIN(n16476), .COUT(n16477), .S0(d1_71__N_418_adj_5756[58]), 
          .S1(d1_71__N_418_adj_5756[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_23 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n123_adj_2845), .D0(d1_adj_5740[56]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n120_adj_2846), .D1(d1_adj_5740[57]), 
          .CIN(n16475), .COUT(n16476), .S0(d1_71__N_418_adj_5756[56]), 
          .S1(d1_71__N_418_adj_5756[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_21 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n129_adj_2843), .D0(d1_adj_5740[54]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n126_adj_2844), .D1(d1_adj_5740[55]), 
          .CIN(n16474), .COUT(n16475), .S0(d1_71__N_418_adj_5756[54]), 
          .S1(d1_71__N_418_adj_5756[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_19 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n135_adj_2841), .D0(d1_adj_5740[52]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n132_adj_2842), .D1(d1_adj_5740[53]), 
          .CIN(n16473), .COUT(n16474), .S0(d1_71__N_418_adj_5756[52]), 
          .S1(d1_71__N_418_adj_5756[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_17 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n141_adj_2839), .D0(d1_adj_5740[50]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n138_adj_2840), .D1(d1_adj_5740[51]), 
          .CIN(n16472), .COUT(n16473), .S0(d1_71__N_418_adj_5756[50]), 
          .S1(d1_71__N_418_adj_5756[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_15 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n147_adj_2837), .D0(d1_adj_5740[48]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n144_adj_2838), .D1(d1_adj_5740[49]), 
          .CIN(n16471), .COUT(n16472), .S0(d1_71__N_418_adj_5756[48]), 
          .S1(d1_71__N_418_adj_5756[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_13 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n153_adj_2835), .D0(d1_adj_5740[46]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n150_adj_2836), .D1(d1_adj_5740[47]), 
          .CIN(n16470), .COUT(n16471), .S0(d1_71__N_418_adj_5756[46]), 
          .S1(d1_71__N_418_adj_5756[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_11 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n159_adj_2833), .D0(d1_adj_5740[44]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n156_adj_2834), .D1(d1_adj_5740[45]), 
          .CIN(n16469), .COUT(n16470), .S0(d1_71__N_418_adj_5756[44]), 
          .S1(d1_71__N_418_adj_5756[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_9 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n165_adj_2831), .D0(d1_adj_5740[42]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n162_adj_2832), .D1(d1_adj_5740[43]), 
          .CIN(n16468), .COUT(n16469), .S0(d1_71__N_418_adj_5756[42]), 
          .S1(d1_71__N_418_adj_5756[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_7 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n171_adj_2829), .D0(d1_adj_5740[40]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n168_adj_2830), .D1(d1_adj_5740[41]), 
          .CIN(n16467), .COUT(n16468), .S0(d1_71__N_418_adj_5756[40]), 
          .S1(d1_71__N_418_adj_5756[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_5 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n177_adj_2827), .D0(d1_adj_5740[38]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n174_adj_2828), .D1(d1_adj_5740[39]), 
          .CIN(n16466), .COUT(n16467), .S0(d1_71__N_418_adj_5756[38]), 
          .S1(d1_71__N_418_adj_5756[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_3 (.A0(MixerOutCos[11]), .B0(cout_adj_5327), 
          .C0(n183_adj_2825), .D0(d1_adj_5740[36]), .A1(MixerOutCos[11]), 
          .B1(cout_adj_5327), .C1(n180_adj_2826), .D1(d1_adj_5740[37]), 
          .CIN(n16465), .COUT(n16466), .S0(d1_71__N_418_adj_5756[36]), 
          .S1(d1_71__N_418_adj_5756[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1504_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1504_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1504_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5327), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16465));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1504_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1504_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1504_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1504_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_38 (.A0(d_d_tmp[71]), .B0(d_tmp[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16461), .S0(n78_adj_5480));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1552_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_36 (.A0(d_d_tmp[69]), .B0(d_tmp[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[70]), .B1(d_tmp[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16460), .COUT(n16461), .S0(n84_adj_5482), 
          .S1(n81_adj_5481));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_34 (.A0(d_d_tmp[67]), .B0(d_tmp[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[68]), .B1(d_tmp[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16459), .COUT(n16460), .S0(n90_adj_5484), 
          .S1(n87_adj_5483));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_32 (.A0(d_d_tmp[65]), .B0(d_tmp[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[66]), .B1(d_tmp[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16458), .COUT(n16459), .S0(n96_adj_5486), 
          .S1(n93_adj_5485));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_30 (.A0(d_d_tmp[63]), .B0(d_tmp[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[64]), .B1(d_tmp[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16457), .COUT(n16458), .S0(n102_adj_5488), 
          .S1(n99_adj_5487));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_28 (.A0(d_d_tmp[61]), .B0(d_tmp[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[62]), .B1(d_tmp[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16456), .COUT(n16457), .S0(n108_adj_5490), 
          .S1(n105_adj_5489));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_26 (.A0(d_d_tmp[59]), .B0(d_tmp[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[60]), .B1(d_tmp[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16455), .COUT(n16456), .S0(n114_adj_5492), 
          .S1(n111_adj_5491));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_24 (.A0(d_d_tmp[57]), .B0(d_tmp[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[58]), .B1(d_tmp[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16454), .COUT(n16455), .S0(n120_adj_5494), 
          .S1(n117_adj_5493));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_22 (.A0(d_d_tmp[55]), .B0(d_tmp[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[56]), .B1(d_tmp[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16453), .COUT(n16454), .S0(n126_adj_5496), 
          .S1(n123_adj_5495));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_20 (.A0(d_d_tmp[53]), .B0(d_tmp[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[54]), .B1(d_tmp[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16452), .COUT(n16453), .S0(n132_adj_5498), 
          .S1(n129_adj_5497));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_18 (.A0(d_d_tmp[51]), .B0(d_tmp[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[52]), .B1(d_tmp[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16451), .COUT(n16452), .S0(n138_adj_5500), 
          .S1(n135_adj_5499));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_16 (.A0(d_d_tmp[49]), .B0(d_tmp[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[50]), .B1(d_tmp[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16450), .COUT(n16451), .S0(n144_adj_5502), 
          .S1(n141_adj_5501));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_14 (.A0(d_d_tmp[47]), .B0(d_tmp[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[48]), .B1(d_tmp[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16449), .COUT(n16450), .S0(n150_adj_5504), 
          .S1(n147_adj_5503));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_12 (.A0(d_d_tmp[45]), .B0(d_tmp[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[46]), .B1(d_tmp[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16448), .COUT(n16449), .S0(n156_adj_5506), 
          .S1(n153_adj_5505));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_10 (.A0(d_d_tmp[43]), .B0(d_tmp[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[44]), .B1(d_tmp[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16447), .COUT(n16448), .S0(n162_adj_5508), 
          .S1(n159_adj_5507));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_8 (.A0(d_d_tmp[41]), .B0(d_tmp[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[42]), .B1(d_tmp[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16446), .COUT(n16447), .S0(n168_adj_5510), 
          .S1(n165_adj_5509));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_6 (.A0(d_d_tmp[39]), .B0(d_tmp[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[40]), .B1(d_tmp[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16445), .COUT(n16446), .S0(n174_adj_5512), 
          .S1(n171_adj_5511));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_4 (.A0(d_d_tmp[37]), .B0(d_tmp[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[38]), .B1(d_tmp[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16444), .COUT(n16445), .S0(n180_adj_5514), 
          .S1(n177_adj_5513));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1552_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1552_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d_tmp[36]), .B1(d_tmp[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16444), .S1(n183_adj_5515));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam _add_1_1552_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1552_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1552_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1552_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_37 (.A0(d7[70]), .B0(cout_adj_5325), .C0(n81_adj_5040), 
          .D0(n3_adj_4750), .A1(d7[71]), .B1(cout_adj_5325), .C1(n78_adj_5039), 
          .D1(n2_adj_4751), .CIN(n16442), .S0(d8_71__N_1603[70]), .S1(d8_71__N_1603[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_35 (.A0(d7[68]), .B0(cout_adj_5325), .C0(n87_adj_5042), 
          .D0(n5_adj_4748), .A1(d7[69]), .B1(cout_adj_5325), .C1(n84_adj_5041), 
          .D1(n4_adj_4749), .CIN(n16441), .COUT(n16442), .S0(d8_71__N_1603[68]), 
          .S1(d8_71__N_1603[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_33 (.A0(d7[66]), .B0(cout_adj_5325), .C0(n93_adj_5044), 
          .D0(n7_adj_4717), .A1(d7[67]), .B1(cout_adj_5325), .C1(n90_adj_5043), 
          .D1(n6_adj_4746), .CIN(n16440), .COUT(n16441), .S0(d8_71__N_1603[66]), 
          .S1(d8_71__N_1603[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_31 (.A0(d7[64]), .B0(cout_adj_5325), .C0(n99_adj_5046), 
          .D0(n9_adj_4684), .A1(d7[65]), .B1(cout_adj_5325), .C1(n96_adj_5045), 
          .D1(n8_adj_4714), .CIN(n16439), .COUT(n16440), .S0(d8_71__N_1603[64]), 
          .S1(d8_71__N_1603[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_29 (.A0(d7[62]), .B0(cout_adj_5325), .C0(n105_adj_5048), 
          .D0(n11_adj_4651), .A1(d7[63]), .B1(cout_adj_5325), .C1(n102_adj_5047), 
          .D1(n10_adj_4676), .CIN(n16438), .COUT(n16439), .S0(d8_71__N_1603[62]), 
          .S1(d8_71__N_1603[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_27 (.A0(d7[60]), .B0(cout_adj_5325), .C0(n111_adj_5050), 
          .D0(n13_adj_4636), .A1(d7[61]), .B1(cout_adj_5325), .C1(n108_adj_5049), 
          .D1(n12_adj_4638), .CIN(n16437), .COUT(n16438), .S0(d8_71__N_1603[60]), 
          .S1(d8_71__N_1603[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_25 (.A0(d7[58]), .B0(cout_adj_5325), .C0(n117_adj_5052), 
          .D0(n15_adj_4634), .A1(d7[59]), .B1(cout_adj_5325), .C1(n114_adj_5051), 
          .D1(n14_adj_4635), .CIN(n16436), .COUT(n16437), .S0(d8_71__N_1603[58]), 
          .S1(d8_71__N_1603[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_23 (.A0(d7[56]), .B0(cout_adj_5325), .C0(n123_adj_5054), 
          .D0(n17_adj_4632), .A1(d7[57]), .B1(cout_adj_5325), .C1(n120_adj_5053), 
          .D1(n16_adj_4633), .CIN(n16435), .COUT(n16436), .S0(d8_71__N_1603[56]), 
          .S1(d8_71__N_1603[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_21 (.A0(d7[54]), .B0(cout_adj_5325), .C0(n129_adj_5056), 
          .D0(n19_adj_4630), .A1(d7[55]), .B1(cout_adj_5325), .C1(n126_adj_5055), 
          .D1(n18_adj_4631), .CIN(n16434), .COUT(n16435), .S0(d8_71__N_1603[54]), 
          .S1(d8_71__N_1603[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_19 (.A0(d7[52]), .B0(cout_adj_5325), .C0(n135_adj_5058), 
          .D0(n21_adj_4628), .A1(d7[53]), .B1(cout_adj_5325), .C1(n132_adj_5057), 
          .D1(n20_adj_4629), .CIN(n16433), .COUT(n16434), .S0(d8_71__N_1603[52]), 
          .S1(d8_71__N_1603[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_17 (.A0(d7[50]), .B0(cout_adj_5325), .C0(n141_adj_5060), 
          .D0(n23_adj_4856), .A1(d7[51]), .B1(cout_adj_5325), .C1(n138_adj_5059), 
          .D1(n22_adj_4879), .CIN(n16432), .COUT(n16433), .S0(d8_71__N_1603[50]), 
          .S1(d8_71__N_1603[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_17.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_30 (.A0(phase_inc_carrGen1[28]), .B0(phase_accum_adj_5732[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[29]), .B1(phase_accum_adj_5732[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15936), .COUT(n15937), .S0(n237), 
          .S1(n234));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_30.INIT0 = 16'h666a;
    defparam phase_accum_add_4_30.INIT1 = 16'h666a;
    defparam phase_accum_add_4_30.INJECT1_0 = "NO";
    defparam phase_accum_add_4_30.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_28 (.A0(phase_inc_carrGen1[26]), .B0(phase_accum_adj_5732[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[27]), .B1(phase_accum_adj_5732[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15935), .COUT(n15936), .S0(n243), 
          .S1(n240));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_28.INIT0 = 16'h666a;
    defparam phase_accum_add_4_28.INIT1 = 16'h666a;
    defparam phase_accum_add_4_28.INJECT1_0 = "NO";
    defparam phase_accum_add_4_28.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_26 (.A0(phase_inc_carrGen1[24]), .B0(phase_accum_adj_5732[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[25]), .B1(phase_accum_adj_5732[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15934), .COUT(n15935), .S0(n249), 
          .S1(n246));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_26.INIT0 = 16'h666a;
    defparam phase_accum_add_4_26.INIT1 = 16'h666a;
    defparam phase_accum_add_4_26.INJECT1_0 = "NO";
    defparam phase_accum_add_4_26.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_24 (.A0(phase_inc_carrGen1[22]), .B0(phase_accum_adj_5732[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[23]), .B1(phase_accum_adj_5732[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15933), .COUT(n15934), .S0(n255), 
          .S1(n252));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_24.INIT0 = 16'h666a;
    defparam phase_accum_add_4_24.INIT1 = 16'h666a;
    defparam phase_accum_add_4_24.INJECT1_0 = "NO";
    defparam phase_accum_add_4_24.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_22 (.A0(phase_inc_carrGen1[20]), .B0(phase_accum_adj_5732[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[21]), .B1(phase_accum_adj_5732[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15932), .COUT(n15933), .S0(n261), 
          .S1(n258));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_22.INIT0 = 16'h666a;
    defparam phase_accum_add_4_22.INIT1 = 16'h666a;
    defparam phase_accum_add_4_22.INJECT1_0 = "NO";
    defparam phase_accum_add_4_22.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_20 (.A0(phase_inc_carrGen1[18]), .B0(phase_accum_adj_5732[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[19]), .B1(phase_accum_adj_5732[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15931), .COUT(n15932), .S0(n267), 
          .S1(n264));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_20.INIT0 = 16'h666a;
    defparam phase_accum_add_4_20.INIT1 = 16'h666a;
    defparam phase_accum_add_4_20.INJECT1_0 = "NO";
    defparam phase_accum_add_4_20.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_18 (.A0(phase_inc_carrGen1[16]), .B0(phase_accum_adj_5732[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[17]), .B1(phase_accum_adj_5732[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15930), .COUT(n15931), .S0(n273), 
          .S1(n270));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_18.INIT0 = 16'h666a;
    defparam phase_accum_add_4_18.INIT1 = 16'h666a;
    defparam phase_accum_add_4_18.INJECT1_0 = "NO";
    defparam phase_accum_add_4_18.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_16 (.A0(phase_inc_carrGen1[14]), .B0(phase_accum_adj_5732[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[15]), .B1(phase_accum_adj_5732[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15929), .COUT(n15930), .S0(n279), 
          .S1(n276));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_16.INIT0 = 16'h666a;
    defparam phase_accum_add_4_16.INIT1 = 16'h666a;
    defparam phase_accum_add_4_16.INJECT1_0 = "NO";
    defparam phase_accum_add_4_16.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_14 (.A0(phase_inc_carrGen1[12]), .B0(phase_accum_adj_5732[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[13]), .B1(phase_accum_adj_5732[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15928), .COUT(n15929), .S0(n285), 
          .S1(n282));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_14.INIT0 = 16'h666a;
    defparam phase_accum_add_4_14.INIT1 = 16'h666a;
    defparam phase_accum_add_4_14.INJECT1_0 = "NO";
    defparam phase_accum_add_4_14.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_12 (.A0(phase_inc_carrGen1[10]), .B0(phase_accum_adj_5732[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[11]), .B1(phase_accum_adj_5732[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15927), .COUT(n15928), .S0(n291), 
          .S1(n288));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_12.INIT0 = 16'h666a;
    defparam phase_accum_add_4_12.INIT1 = 16'h666a;
    defparam phase_accum_add_4_12.INJECT1_0 = "NO";
    defparam phase_accum_add_4_12.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_10 (.A0(phase_inc_carrGen1[8]), .B0(phase_accum_adj_5732[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[9]), .B1(phase_accum_adj_5732[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15926), .COUT(n15927), .S0(n297), 
          .S1(n294));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_10.INIT0 = 16'h666a;
    defparam phase_accum_add_4_10.INIT1 = 16'h666a;
    defparam phase_accum_add_4_10.INJECT1_0 = "NO";
    defparam phase_accum_add_4_10.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_8 (.A0(phase_inc_carrGen1[6]), .B0(phase_accum_adj_5732[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[7]), .B1(phase_accum_adj_5732[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15925), .COUT(n15926), .S0(n303), 
          .S1(n300));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_8.INIT0 = 16'h666a;
    defparam phase_accum_add_4_8.INIT1 = 16'h666a;
    defparam phase_accum_add_4_8.INJECT1_0 = "NO";
    defparam phase_accum_add_4_8.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_6 (.A0(phase_inc_carrGen1[4]), .B0(phase_accum_adj_5732[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[5]), .B1(phase_accum_adj_5732[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15924), .COUT(n15925), .S0(n309), 
          .S1(n306));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_6.INIT0 = 16'h666a;
    defparam phase_accum_add_4_6.INIT1 = 16'h666a;
    defparam phase_accum_add_4_6.INJECT1_0 = "NO";
    defparam phase_accum_add_4_6.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_4 (.A0(phase_inc_carrGen1[2]), .B0(phase_accum_adj_5732[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[3]), .B1(phase_accum_adj_5732[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15923), .COUT(n15924), .S0(n315), 
          .S1(n312));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_4.INIT0 = 16'h666a;
    defparam phase_accum_add_4_4.INIT1 = 16'h666a;
    defparam phase_accum_add_4_4.INJECT1_0 = "NO";
    defparam phase_accum_add_4_4.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_2 (.A0(phase_inc_carrGen1[0]), .B0(phase_accum_adj_5732[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_carrGen1[1]), .B1(phase_accum_adj_5732[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15923), .S1(n318));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(39[24:52])
    defparam phase_accum_add_4_2.INIT0 = 16'h0008;
    defparam phase_accum_add_4_2.INIT1 = 16'h666a;
    defparam phase_accum_add_4_2.INJECT1_0 = "NO";
    defparam phase_accum_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_38 (.A0(d_d6[71]), .B0(d6[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15921), .S0(n78_adj_5075));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1648_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_36 (.A0(d_d6[69]), .B0(d6[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[70]), .B1(d6[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15920), .COUT(n15921), .S0(n84_adj_5077), .S1(n81_adj_5076));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_34 (.A0(d_d6[67]), .B0(d6[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[68]), .B1(d6[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15919), .COUT(n15920), .S0(n90_adj_5079), .S1(n87_adj_5078));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_32 (.A0(d_d6[65]), .B0(d6[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[66]), .B1(d6[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15918), .COUT(n15919), .S0(n96_adj_5081), .S1(n93_adj_5080));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_30 (.A0(d_d6[63]), .B0(d6[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[64]), .B1(d6[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15917), .COUT(n15918), .S0(n102_adj_5083), .S1(n99_adj_5082));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_28 (.A0(d_d6[61]), .B0(d6[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[62]), .B1(d6[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15916), .COUT(n15917), .S0(n108_adj_5085), .S1(n105_adj_5084));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_26 (.A0(d_d6[59]), .B0(d6[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[60]), .B1(d6[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15915), .COUT(n15916), .S0(n114_adj_5087), .S1(n111_adj_5086));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_24 (.A0(d_d6[57]), .B0(d6[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[58]), .B1(d6[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15914), .COUT(n15915), .S0(n120_adj_5089), .S1(n117_adj_5088));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_22 (.A0(d_d6[55]), .B0(d6[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[56]), .B1(d6[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15913), .COUT(n15914), .S0(n126_adj_5091), .S1(n123_adj_5090));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_20 (.A0(d_d6[53]), .B0(d6[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[54]), .B1(d6[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15912), .COUT(n15913), .S0(n132_adj_5093), .S1(n129_adj_5092));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_18 (.A0(d_d6[51]), .B0(d6[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[52]), .B1(d6[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15911), .COUT(n15912), .S0(n138_adj_5095), .S1(n135_adj_5094));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_16 (.A0(d_d6[49]), .B0(d6[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[50]), .B1(d6[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15910), .COUT(n15911), .S0(n144_adj_5097), .S1(n141_adj_5096));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_14 (.A0(d_d6[47]), .B0(d6[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[48]), .B1(d6[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15909), .COUT(n15910), .S0(n150_adj_5099), .S1(n147_adj_5098));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_12 (.A0(d_d6[45]), .B0(d6[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[46]), .B1(d6[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15908), .COUT(n15909), .S0(n156_adj_5101), .S1(n153_adj_5100));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_10 (.A0(d_d6[43]), .B0(d6[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[44]), .B1(d6[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15907), .COUT(n15908), .S0(n162_adj_5103), .S1(n159_adj_5102));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_8 (.A0(d_d6[41]), .B0(d6[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[42]), .B1(d6[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15906), .COUT(n15907), .S0(n168_adj_5105), .S1(n165_adj_5104));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_6 (.A0(d_d6[39]), .B0(d6[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[40]), .B1(d6[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15905), .COUT(n15906), .S0(n174_adj_5107), .S1(n171_adj_5106));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_4 (.A0(d_d6[37]), .B0(d6[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[38]), .B1(d6[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15904), .COUT(n15905), .S0(n180_adj_5109), .S1(n177_adj_5108));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1648_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1648_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6[36]), .B1(d6[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15904), .S1(n183_adj_5110));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1648_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1648_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1648_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1648_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_17 (.A0(count_adj_5755[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15903), .S0(n36_adj_5400));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1442_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1442_add_4_17.INIT1 = 16'h0000;
    defparam _add_1_1442_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_15 (.A0(count_adj_5755[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5755[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15902), .COUT(n15903), .S0(n42_adj_5402), 
          .S1(n39_adj_5401));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1442_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1442_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1442_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_13 (.A0(count_adj_5755[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5755[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15901), .COUT(n15902), .S0(n48_adj_5404), 
          .S1(n45_adj_5403));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1442_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1442_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1442_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_11 (.A0(count_adj_5755[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5755[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15900), .COUT(n15901), .S0(n54_adj_5406), 
          .S1(n51_adj_5405));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1442_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1442_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1442_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_9 (.A0(count_adj_5755[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5755[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15899), .COUT(n15900), .S0(n60_adj_5408), 
          .S1(n57_adj_5407));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1442_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1442_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1442_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_7 (.A0(count_adj_5755[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5755[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15898), .COUT(n15899), .S0(n66_adj_5410), 
          .S1(n63_adj_5409));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1442_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1442_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1442_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_5 (.A0(count_adj_5755[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5755[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15897), .COUT(n15898), .S0(n72_adj_5412), 
          .S1(n69_adj_5411));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1442_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1442_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1442_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_3 (.A0(count_adj_5755[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_5755[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15896), .COUT(n15897), .S0(n78_adj_5414), 
          .S1(n75_adj_5413));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1442_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1442_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1442_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1442_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_adj_5755[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15896), .S1(n81_adj_5415));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(79[26:39])
    defparam _add_1_1442_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1442_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1442_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1442_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_38 (.A0(d3[71]), .B0(d2[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15895), .S0(n78_adj_5552));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1561_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1561_add_4_36 (.A0(d3[69]), .B0(d2[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(d3[70]), .B1(d2[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15894), .COUT(n15895), .S0(n84_adj_5554), .S1(n81_adj_5553));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1561_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1561_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1561_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1561_add_4_36.INJECT1_1 = "NO";
    LUT4 mux_325_i7_4_lut (.A(n2565), .B(n301), .C(n17925), .D(n2572), 
         .Z(n2365)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i7_4_lut.init = 16'hc0ca;
    LUT4 i1_2_lut_rep_160 (.A(led_c_4), .B(n17069), .Z(n17932)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_160.init = 16'h8888;
    LUT4 mux_325_i11_4_lut (.A(n12086), .B(n289), .C(n17925), .D(n2572), 
         .Z(n2361)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i11_4_lut.init = 16'hc0ca;
    LUT4 i2490_4_lut (.A(n133_adj_5416), .B(n127), .C(led_c_3), .D(n17932), 
         .Z(n12304)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2490_4_lut.init = 16'hcac0;
    LUT4 i2476_4_lut (.A(n286), .B(n280_adj_5681), .C(led_c_3), .D(n17932), 
         .Z(n12290)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2476_4_lut.init = 16'hcac0;
    LUT4 i13_4_lut_then_4_lut (.A(led_c_3), .B(n17937), .C(n17069), .D(led_c_4), 
         .Z(n17953)) /* synthesis lut_function=(!(A+!(B (C (D))+!B ((D)+!C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i13_4_lut_then_4_lut.init = 16'h5101;
    LUT4 i13_4_lut_else_4_lut (.A(led_c_3), .B(n17937), .C(n17069), .Z(n17952)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i13_4_lut_else_4_lut.init = 16'h0101;
    LUT4 i3155_2_lut (.A(led_c_4), .B(n2824), .Z(n3660)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i3155_2_lut.init = 16'h4444;
    FD1S3AX o_Rx_Byte_i4_rep_181 (.D(o_Rx_Byte1[3]), .CK(clk_80mhz), .Q(n18076));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam o_Rx_Byte_i4_rep_181.GSR = "ENABLED";
    LUT4 i2492_4_lut (.A(n130), .B(n124), .C(led_c_3), .D(n17932), .Z(n12306)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2492_4_lut.init = 16'hcac0;
    LUT4 mux_325_i9_4_lut (.A(n12082), .B(n295), .C(n17925), .D(n2572), 
         .Z(n2363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i9_4_lut.init = 16'hcfca;
    LUT4 i6354_4_lut (.A(n18121), .B(led_c_3), .C(n17926), .D(n17932), 
         .Z(clk_80mhz_enable_1470)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))) */ ;
    defparam i6354_4_lut.init = 16'ha0a2;
    LUT4 i6362_4_lut (.A(led_c_2), .B(n17939), .C(led_c_3), .D(led_c_6), 
         .Z(clk_80mhz_enable_1407)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i6362_4_lut.init = 16'h0004;
    LUT4 i6298_4_lut (.A(r_Rx_Byte[6]), .B(r_Rx_Data), .C(n17397), .D(n17943), 
         .Z(n17664)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i6298_4_lut.init = 16'hcaaa;
    LUT4 i5379_2_lut (.A(d1_adj_5740[0]), .B(MixerOutCos[0]), .Z(d1_71__N_418_adj_5756[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5379_2_lut.init = 16'h6666;
    LUT4 i5357_2_lut (.A(MultResult2[0]), .B(MultResult1[0]), .Z(n126_adj_5442)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5357_2_lut.init = 16'h6666;
    LUT4 i2334_3_lut_4_lut (.A(n18075), .B(n17937), .C(led_c_3), .D(n205_adj_5656), 
         .Z(n12132)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2334_3_lut_4_lut.init = 16'hf404;
    LUT4 i1_3_lut_rep_165_4_lut_4_lut (.A(led_c_0), .B(n17951), .C(n17948), 
         .D(led_c_6), .Z(n17937)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_3_lut_rep_165_4_lut_4_lut.init = 16'h4000;
    CCU2C add_3828_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n17205), .B1(n12983), .C1(led_c_4), .D1(n2824), .COUT(n16612));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam add_3828_1.INIT0 = 16'h0000;
    defparam add_3828_1.INIT1 = 16'hf7ff;
    defparam add_3828_1.INJECT1_0 = "NO";
    defparam add_3828_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut (.A(led_c_0), .B(n18076), .C(led_c_1), .D(led_c_2), 
         .Z(n17097)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_4_lut.init = 16'hfffd;
    LUT4 i1_4_lut (.A(n18075), .B(n17940), .C(led_c_0), .D(led_c_1), 
         .Z(n17069)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut.init = 16'h0040;
    LUT4 i2304_3_lut_4_lut (.A(n18075), .B(n17937), .C(led_c_3), .D(n253_adj_5672), 
         .Z(n12102)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2304_3_lut_4_lut.init = 16'hf707;
    LUT4 i5347_2_lut (.A(d2[0]), .B(d1[0]), .Z(d2_71__N_490[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5347_2_lut.init = 16'h6666;
    LUT4 i3293_2_lut_2_lut (.A(led_c_3), .B(n226_adj_5663), .Z(n2542)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i3293_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2294_3_lut_4_lut (.A(n18075), .B(n17937), .C(n18076), .D(n271_adj_5678), 
         .Z(n12092)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2294_3_lut_4_lut.init = 16'hf808;
    LUT4 i3299_2_lut_2_lut (.A(n18076), .B(n145_adj_5636), .Z(n2515)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i3299_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2284_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(led_c_3), .D(n289_adj_5684), 
         .Z(n12082)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2284_3_lut_4_lut.init = 16'hf808;
    LUT4 i3226_2_lut_2_lut (.A(led_c_3), .B(n292_adj_5685), .Z(n2430)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i3226_2_lut_2_lut.init = 16'hdddd;
    LUT4 i359_2_lut_3_lut_3_lut (.A(led_c_3), .B(n17069), .C(led_c_4), 
         .Z(n2572)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i359_2_lut_3_lut_3_lut.init = 16'h0404;
    LUT4 i3228_2_lut_2_lut (.A(led_c_3), .B(n268_adj_5677), .Z(n2422)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i3228_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2332_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(led_c_3), .D(n208_adj_5657), 
         .Z(n12130)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2332_3_lut_4_lut.init = 16'hf404;
    LUT4 i2324_3_lut_4_lut (.A(n18075), .B(n17937), .C(n18076), .D(n220_adj_5661), 
         .Z(n12122)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2324_3_lut_4_lut.init = 16'hf404;
    LUT4 i348_2_lut_rep_153_3_lut_3_lut (.A(led_c_3), .B(n17069), .C(led_c_4), 
         .Z(n17925)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i348_2_lut_rep_153_3_lut_3_lut.init = 16'h4040;
    CCU2C add_3826_11 (.A0(ISquare[31]), .B0(n17942), .C0(n17938), .D0(VCC_net), 
          .A1(ISquare[31]), .B1(n17942), .C1(n17938), .D1(VCC_net), 
          .CIN(n16607), .S0(n29_adj_5606), .S1(d_out_d_11__N_1874[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3826_11.INIT0 = 16'he1e1;
    defparam add_3826_11.INIT1 = 16'he1e1;
    defparam add_3826_11.INJECT1_0 = "NO";
    defparam add_3826_11.INJECT1_1 = "NO";
    LUT4 i2_2_lut_3_lut_3_lut (.A(led_c_3), .B(n17937), .C(led_c_2), .Z(n16718)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i2_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 i5342_2_lut (.A(d3[0]), .B(d2[0]), .Z(d3_71__N_562[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5342_2_lut.init = 16'h6666;
    LUT4 i2318_3_lut_4_lut (.A(n18075), .B(n17937), .C(n18076), .D(n229_adj_5664), 
         .Z(n12116)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2318_3_lut_4_lut.init = 16'hf404;
    LUT4 i5348_2_lut (.A(d4[0]), .B(d3[0]), .Z(d4_71__N_634[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5348_2_lut.init = 16'h6666;
    LUT4 i27_3_lut_3_lut (.A(n18076), .B(n17937), .C(n247_adj_5670), .Z(n13_adj_4794)) /* synthesis lut_function=(!(A (C)+!A !(B))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i27_3_lut_3_lut.init = 16'h4e4e;
    LUT4 i2286_3_lut_4_lut (.A(n18075), .B(n17937), .C(n18076), .D(n286_adj_5683), 
         .Z(n12084)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2286_3_lut_4_lut.init = 16'hf707;
    LUT4 i5381_2_lut (.A(d5[0]), .B(d4[0]), .Z(d5_71__N_706[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5381_2_lut.init = 16'h6666;
    CCU2C add_3826_9 (.A0(n17938), .B0(ISquare[31]), .C0(ISquare[23]), 
          .D0(ISquare[22]), .A1(n23_adj_2823), .B1(n15173), .C1(n213_adj_4637), 
          .D1(ISquare[31]), .CIN(n16606), .COUT(n16607), .S0(n35_adj_5608), 
          .S1(n32_adj_5607));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3826_9.INIT0 = 16'h6665;
    defparam add_3826_9.INIT1 = 16'h556a;
    defparam add_3826_9.INJECT1_0 = "NO";
    defparam add_3826_9.INJECT1_1 = "NO";
    LUT4 i2312_3_lut_4_lut (.A(n18075), .B(n17937), .C(n18076), .D(n238_adj_5667), 
         .Z(n12110)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2312_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_325_i61_4_lut (.A(n12172), .B(n139), .C(n17925), .D(n2572), 
         .Z(n2311)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i61_4_lut.init = 16'hc0ca;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(led_c_3), .B(n17937), .C(n17069), 
         .D(led_c_4), .Z(n27_adj_5727)) /* synthesis lut_function=(!(A+!(B+!((D)+!C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h4454;
    CCU2C add_3826_7 (.A0(n32_adj_2822), .B0(ISquare[31]), .C0(ISquare[23]), 
          .D0(ISquare[22]), .A1(n17942), .B1(ISquare[31]), .C1(ISquare[23]), 
          .D1(ISquare[22]), .CIN(n16605), .COUT(n16606), .S0(n41_adj_5609), 
          .S1(n38));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3826_7.INIT0 = 16'h999a;
    defparam add_3826_7.INIT1 = 16'haaa9;
    defparam add_3826_7.INJECT1_0 = "NO";
    defparam add_3826_7.INJECT1_1 = "NO";
    CCU2C add_3826_5 (.A0(ISquare[22]), .B0(ISquare[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[23]), .B1(ISquare[22]), .C1(ISquare[31]), 
          .D1(n15173), .CIN(n16604), .COUT(n16605), .S0(n47_adj_5611), 
          .S1(n44_adj_5610));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3826_5.INIT0 = 16'h9999;
    defparam add_3826_5.INIT1 = 16'heee1;
    defparam add_3826_5.INJECT1_0 = "NO";
    defparam add_3826_5.INJECT1_1 = "NO";
    CCU2C add_3826_3 (.A0(ISquare[31]), .B0(n17942), .C0(ISquare[20]), 
          .D0(VCC_net), .A1(ISquare[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16603), .COUT(n16604), .S1(n50_adj_5612));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3826_3.INIT0 = 16'he1e1;
    defparam add_3826_3.INIT1 = 16'h555f;
    defparam add_3826_3.INJECT1_0 = "NO";
    defparam add_3826_3.INJECT1_1 = "NO";
    CCU2C add_3826_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(ISquare[22]), .B1(ISquare[23]), .C1(n213_adj_4637), .D1(ISquare[31]), 
          .COUT(n16603));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3826_1.INIT0 = 16'h0000;
    defparam add_3826_1.INIT1 = 16'h001f;
    defparam add_3826_1.INJECT1_0 = "NO";
    defparam add_3826_1.INJECT1_1 = "NO";
    LUT4 mux_325_i8_4_lut (.A(n27_adj_5727), .B(n298), .C(n17925), .D(n2430), 
         .Z(n2364)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i8_4_lut.init = 16'hc5c0;
    LUT4 i2488_4_lut (.A(n136_adj_5417), .B(n130_adj_5631), .C(led_c_3), 
         .D(n17932), .Z(n12302)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2488_4_lut.init = 16'hcac0;
    LUT4 mux_325_i5_4_lut (.A(n12076), .B(n307), .C(n17925), .D(n2572), 
         .Z(n2367)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i5_4_lut.init = 16'hcfca;
    LUT4 i2350_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(n18076), .D(n175_adj_5646), 
         .Z(n12148)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2350_3_lut_4_lut.init = 16'hf707;
    LUT4 i2344_3_lut_4_lut (.A(n18075), .B(n17937), .C(led_c_3), .D(n187_adj_5650), 
         .Z(n12142)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2344_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_325_i6_4_lut (.A(n12078), .B(n304), .C(n17925), .D(n2572), 
         .Z(n2366)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i6_4_lut.init = 16'hc0ca;
    LUT4 i27_3_lut_3_lut_adj_61 (.A(led_c_3), .B(n17937), .C(n193_adj_5652), 
         .Z(n13_adj_5726)) /* synthesis lut_function=(!(A (C)+!A !(B))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i27_3_lut_3_lut_adj_61.init = 16'h4e4e;
    LUT4 i3231_2_lut_2_lut (.A(led_c_3), .B(n181_adj_5648), .Z(n2393)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i3231_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2308_3_lut_4_lut (.A(n18075), .B(n17937), .C(led_c_3), .D(n244_adj_5669), 
         .Z(n12106)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2308_3_lut_4_lut.init = 16'hf404;
    LUT4 i3283_2_lut_2_lut (.A(n18076), .B(n295_adj_5686), .Z(n2565)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i3283_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut_3_lut (.A(led_c_3), .B(led_c_0), .C(led_c_4), .Z(n17401)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i1_3_lut_3_lut.init = 16'h5454;
    LUT4 i2336_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(n18076), .D(n202_adj_5655), 
         .Z(n12134)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2336_3_lut_4_lut.init = 16'hf707;
    LUT4 i6297_4_lut (.A(r_Rx_Byte[4]), .B(r_Rx_Data), .C(n17946), .D(n17945), 
         .Z(n17663)) /* synthesis lut_function=(A (B+(C+(D)))+!A !((C+(D))+!B)) */ ;
    defparam i6297_4_lut.init = 16'haaac;
    LUT4 i2330_3_lut_4_lut (.A(n18075), .B(n17937), .C(n18076), .D(n211_adj_5658), 
         .Z(n12128)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2330_3_lut_4_lut.init = 16'hf808;
    CCU2C _add_1_1439_add_4_28 (.A0(d5_adj_5744[26]), .B0(d4_adj_5743[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[27]), .B1(d4_adj_5743[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16112), .COUT(n16113), .S0(d5_71__N_706_adj_5760[26]), 
          .S1(d5_71__N_706_adj_5760[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_15 (.A0(d7[48]), .B0(cout_adj_5325), .C0(n147_adj_5062), 
          .D0(n25), .A1(d7[49]), .B1(cout_adj_5325), .C1(n144_adj_5061), 
          .D1(n24), .CIN(n16431), .COUT(n16432), .S0(d8_71__N_1603[48]), 
          .S1(d8_71__N_1603[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_2 (.A0(d5[0]), .B0(d4[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[1]), .B1(d4[1]), .C1(GND_net), .D1(VCC_net), .COUT(n16360), 
          .S1(d5_71__N_706[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1421_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_2.INJECT1_1 = "NO";
    CCU2C add_3834_13 (.A0(d_out_d_11__N_1873), .B0(d_out_d_11__N_1874[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1873), .B1(d_out_d_11__N_1874[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16597), .S0(n33_adj_5186), 
          .S1(d_out_d_11__N_1876[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3834_13.INIT0 = 16'h666a;
    defparam add_3834_13.INIT1 = 16'h666a;
    defparam add_3834_13.INJECT1_0 = "NO";
    defparam add_3834_13.INJECT1_1 = "NO";
    CCU2C add_3834_11 (.A0(d_out_d_11__N_1874[17]), .B0(n32_adj_5607), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), .B1(n29_adj_5606), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16596), .COUT(n16597), .S0(n39), 
          .S1(n36_adj_5187));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3834_11.INIT0 = 16'h9995;
    defparam add_3834_11.INIT1 = 16'h9995;
    defparam add_3834_11.INJECT1_0 = "NO";
    defparam add_3834_11.INJECT1_1 = "NO";
    CCU2C add_3834_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1874[17]), .C0(n38), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1874[17]), 
          .C1(n35_adj_5608), .D1(VCC_net), .CIN(n16595), .COUT(n16596), 
          .S0(n45), .S1(n42));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3834_9.INIT0 = 16'h6969;
    defparam add_3834_9.INIT1 = 16'h6969;
    defparam add_3834_9.INJECT1_0 = "NO";
    defparam add_3834_9.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_13 (.A0(d7[46]), .B0(cout_adj_5325), .C0(n153_adj_5064), 
          .D0(n27), .A1(d7[47]), .B1(cout_adj_5325), .C1(n150_adj_5063), 
          .D1(n26), .CIN(n16430), .COUT(n16431), .S0(d8_71__N_1603[46]), 
          .S1(d8_71__N_1603[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_30 (.A0(d1[28]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[29]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16336), .COUT(n16337), .S0(d1_71__N_418[28]), 
          .S1(d1_71__N_418[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_30.INJECT1_1 = "NO";
    CCU2C add_3834_7 (.A0(d_out_d_11__N_1874[17]), .B0(n44_adj_5610), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1874[17]), 
          .C1(n41_adj_5609), .D1(VCC_net), .CIN(n16594), .COUT(n16595), 
          .S0(n51), .S1(n48));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3834_7.INIT0 = 16'h9995;
    defparam add_3834_7.INIT1 = 16'h6969;
    defparam add_3834_7.INJECT1_0 = "NO";
    defparam add_3834_7.INJECT1_1 = "NO";
    CCU2C add_3834_5 (.A0(n50_adj_5612), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(n17938), .C1(n47_adj_5611), 
          .D1(VCC_net), .CIN(n16593), .COUT(n16594), .S0(n57), .S1(n54));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3834_5.INIT0 = 16'haaa0;
    defparam add_3834_5.INIT1 = 16'h6969;
    defparam add_3834_5.INJECT1_0 = "NO";
    defparam add_3834_5.INJECT1_1 = "NO";
    CCU2C add_3834_3 (.A0(d_out_d_11__N_1874[17]), .B0(ISquare[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16592), .COUT(n16593), .S1(n60));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3834_3.INIT0 = 16'h666a;
    defparam add_3834_3.INIT1 = 16'h555f;
    defparam add_3834_3.INJECT1_0 = "NO";
    defparam add_3834_3.INJECT1_1 = "NO";
    CCU2C add_3834_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16592));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3834_1.INIT0 = 16'h0000;
    defparam add_3834_1.INIT1 = 16'haaaf;
    defparam add_3834_1.INJECT1_0 = "NO";
    defparam add_3834_1.INJECT1_1 = "NO";
    CCU2C add_3827_17 (.A0(ISquare[31]), .B0(n917), .C0(GND_net), .D0(VCC_net), 
          .A1(n916), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16586), 
          .S1(d_out_d_11__N_2401[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3827_17.INIT0 = 16'h666a;
    defparam add_3827_17.INIT1 = 16'haaa0;
    defparam add_3827_17.INJECT1_0 = "NO";
    defparam add_3827_17.INJECT1_1 = "NO";
    CCU2C add_3827_15 (.A0(ISquare[31]), .B0(n919), .C0(GND_net), .D0(VCC_net), 
          .A1(ISquare[31]), .B1(n918), .C1(GND_net), .D1(VCC_net), .CIN(n16585), 
          .COUT(n16586));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3827_15.INIT0 = 16'h666a;
    defparam add_3827_15.INIT1 = 16'h666a;
    defparam add_3827_15.INJECT1_0 = "NO";
    defparam add_3827_15.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_11 (.A0(d7[44]), .B0(cout_adj_5325), .C0(n159_adj_5066), 
          .D0(n29), .A1(d7[45]), .B1(cout_adj_5325), .C1(n156_adj_5065), 
          .D1(n28), .CIN(n16429), .COUT(n16430), .S0(d8_71__N_1603[44]), 
          .S1(d8_71__N_1603[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_11.INJECT1_1 = "NO";
    CCU2C add_3827_13 (.A0(n921), .B0(n15173), .C0(n213_adj_4637), .D0(ISquare[31]), 
          .A1(n920), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n16584), 
          .COUT(n16585));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3827_13.INIT0 = 16'h556a;
    defparam add_3827_13.INIT1 = 16'haaa0;
    defparam add_3827_13.INJECT1_0 = "NO";
    defparam add_3827_13.INJECT1_1 = "NO";
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    CCU2C add_3827_11 (.A0(d_out_d_11__N_1876[17]), .B0(n923), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), .B1(n922), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16583), .COUT(n16584));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3827_11.INIT0 = 16'h9995;
    defparam add_3827_11.INIT1 = 16'h9995;
    defparam add_3827_11.INJECT1_0 = "NO";
    defparam add_3827_11.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_28 (.A0(d1[26]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[27]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16335), .COUT(n16336), .S0(d1_71__N_418[26]), 
          .S1(d1_71__N_418[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_28.INJECT1_1 = "NO";
    CCU2C add_3827_9 (.A0(d_out_d_11__N_1880[17]), .B0(n925), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1878[17]), .B1(n924), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16582), .COUT(n16583));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3827_9.INIT0 = 16'h9995;
    defparam add_3827_9.INIT1 = 16'h9995;
    defparam add_3827_9.INJECT1_0 = "NO";
    defparam add_3827_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_161_3_lut_4_lut_4_lut (.A(led_c_1), .B(led_c_4), .C(n17948), 
         .D(led_c_6), .Z(n17933)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;
    defparam i1_2_lut_rep_161_3_lut_4_lut_4_lut.init = 16'hdfff;
    LUT4 i2316_3_lut_4_lut (.A(n18075), .B(n17937), .C(led_c_3), .D(n232_adj_5665), 
         .Z(n12114)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2316_3_lut_4_lut.init = 16'hf707;
    LUT4 i2314_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(n18076), .D(n235_adj_5666), 
         .Z(n12112)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2314_3_lut_4_lut.init = 16'hf808;
    FD1S3AX o_Rx_Byte_i3_rep_180 (.D(o_Rx_Byte1[2]), .CK(clk_80mhz), .Q(n18075));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam o_Rx_Byte_i3_rep_180.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut_4_lut_4_lut (.A(led_c_1), .B(led_c_0), .C(led_c_4), 
         .D(led_c_3), .Z(n17317)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_4_lut_4_lut_4_lut.init = 16'h0010;
    LUT4 mux_325_i59_4_lut (.A(n12168), .B(n145), .C(n17925), .D(n2572), 
         .Z(n2313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i59_4_lut.init = 16'hcfca;
    LUT4 i2280_3_lut_4_lut (.A(n18075), .B(n17937), .C(n18076), .D(n298_adj_5687), 
         .Z(n12078)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2280_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_3_lut_rep_176 (.A(led_c_5), .B(led_c_7), .C(o_Rx_DV), .Z(n17948)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam i1_3_lut_rep_176.init = 16'h2020;
    LUT4 mux_325_i60_4_lut (.A(n12170), .B(n142), .C(n17925), .D(n2572), 
         .Z(n2312)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i60_4_lut.init = 16'hc0ca;
    LUT4 mux_325_i57_4_lut (.A(n2515), .B(n151), .C(n17925), .D(n2572), 
         .Z(n2315)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i57_4_lut.init = 16'hc0ca;
    LUT4 i2486_4_lut (.A(n148), .B(n142_adj_5635), .C(led_c_3), .D(n17932), 
         .Z(n12300)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2486_4_lut.init = 16'hcac0;
    LUT4 mux_325_i55_4_lut (.A(n12162), .B(n157), .C(n17925), .D(n2572), 
         .Z(n2317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i55_4_lut.init = 16'hcfca;
    LUT4 i25_4_lut (.A(n40_adj_5728), .B(n154), .C(n17925), .D(n27_adj_5727), 
         .Z(n21_adj_5729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i25_4_lut.init = 16'hcfca;
    LUT4 i60_2_lut (.A(led_c_3), .B(n148_adj_5637), .Z(n40_adj_5728)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(44[22:25])
    defparam i60_2_lut.init = 16'h8888;
    LUT4 i2484_4_lut (.A(n163), .B(n157_adj_5640), .C(led_c_3), .D(n17932), 
         .Z(n12298)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2484_4_lut.init = 16'hcac0;
    LUT4 i5416_2_lut_rep_167_4_lut (.A(led_c_5), .B(led_c_7), .C(o_Rx_DV), 
         .D(led_c_4), .Z(n17939)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam i5416_2_lut_rep_167_4_lut.init = 16'h2000;
    LUT4 i5380_2_lut (.A(d1[0]), .B(MixerOutSin[0]), .Z(d1_71__N_418[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5380_2_lut.init = 16'h6666;
    LUT4 i5414_2_lut_rep_168_4_lut (.A(led_c_5), .B(led_c_7), .C(o_Rx_DV), 
         .D(led_c_6), .Z(n17940)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam i5414_2_lut_rep_168_4_lut.init = 16'h2000;
    CCU2C _add_1_add_4_4 (.A0(d_d8[1]), .B0(d8[1]), .C0(GND_net), .D0(VCC_net), 
          .A1(d_d8[2]), .B1(d8[2]), .C1(GND_net), .D1(VCC_net), .CIN(n15198), 
          .COUT(n15199), .S0(d9_71__N_1675[1]), .S1(d9_71__N_1675[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_add_4_4.INJECT1_1 = "NO";
    LUT4 mux_325_i54_4_lut (.A(n12160), .B(n160), .C(n17925), .D(n2572), 
         .Z(n2318)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i54_4_lut.init = 16'hc0ca;
    LUT4 mux_325_i51_4_lut (.A(n2521), .B(n169), .C(n17925), .D(n2572), 
         .Z(n2321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i51_4_lut.init = 16'hcfca;
    LUT4 i5378_2_lut (.A(d2_adj_5741[0]), .B(d1_adj_5740[0]), .Z(d2_71__N_490_adj_5757[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5378_2_lut.init = 16'h6666;
    PLL PLL_inst (.clk_25mhz_c(clk_25mhz_c), .clk_80mhz(clk_80mhz), .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(97[8] 100[5])
    CCU2C _add_1_1439_add_4_26 (.A0(d5_adj_5744[24]), .B0(d4_adj_5743[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(d5_adj_5744[25]), .B1(d4_adj_5743[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16111), .COUT(n16112), .S0(d5_71__N_706_adj_5760[24]), 
          .S1(d5_71__N_706_adj_5760[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1439_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1439_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1439_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1439_add_4_26.INJECT1_1 = "NO";
    CCU2C add_3827_7 (.A0(d_out_d_11__N_1884[17]), .B0(n927), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1882[17]), .B1(n926), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16581), .COUT(n16582));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3827_7.INIT0 = 16'h9995;
    defparam add_3827_7.INIT1 = 16'h9995;
    defparam add_3827_7.INJECT1_0 = "NO";
    defparam add_3827_7.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_9 (.A0(d7[42]), .B0(cout_adj_5325), .C0(n165_adj_5068), 
          .D0(n31), .A1(d7[43]), .B1(cout_adj_5325), .C1(n162_adj_5067), 
          .D1(n30), .CIN(n16428), .COUT(n16429), .S0(d8_71__N_1603[42]), 
          .S1(d8_71__N_1603[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_7 (.A0(d7[40]), .B0(cout_adj_5325), .C0(n171_adj_5070), 
          .D0(n33_adj_4755), .A1(d7[41]), .B1(cout_adj_5325), .C1(n168_adj_5069), 
          .D1(n32_adj_4855), .CIN(n16427), .COUT(n16428), .S0(d8_71__N_1603[40]), 
          .S1(d8_71__N_1603[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_5 (.A0(d7[38]), .B0(cout_adj_5325), .C0(n177_adj_5072), 
          .D0(n35_adj_4753), .A1(d7[39]), .B1(cout_adj_5325), .C1(n174_adj_5071), 
          .D1(n34_adj_4754), .CIN(n16426), .COUT(n16427), .S0(d8_71__N_1603[38]), 
          .S1(d8_71__N_1603[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_26 (.A0(d1[24]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[25]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16334), .COUT(n16335), .S0(d1_71__N_418[24]), 
          .S1(d1_71__N_418[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_26.INJECT1_1 = "NO";
    CCU2C add_3827_5 (.A0(d_out_d_11__N_1888[17]), .B0(n929), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1886[17]), .B1(n928), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16580), .COUT(n16581));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3827_5.INIT0 = 16'h9995;
    defparam add_3827_5.INIT1 = 16'h9995;
    defparam add_3827_5.INJECT1_0 = "NO";
    defparam add_3827_5.INJECT1_1 = "NO";
    LUT4 i3297_2_lut (.A(n163_adj_5642), .B(n18076), .Z(n2521)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i3297_2_lut.init = 16'h8888;
    CCU2C _add_1_1519_add_4_9 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n165_adj_5318), .D0(d1[42]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n162_adj_5317), .D1(d1[43]), .CIN(n16183), .COUT(n16184), 
          .S0(d1_71__N_418[42]), .S1(d1_71__N_418[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_3 (.A0(d7[36]), .B0(cout_adj_5325), .C0(n183_adj_5074), 
          .D0(n37_adj_4747), .A1(d7[37]), .B1(cout_adj_5325), .C1(n180_adj_5073), 
          .D1(n36_adj_4752), .CIN(n16425), .COUT(n16426), .S0(d8_71__N_1603[36]), 
          .S1(d8_71__N_1603[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1465_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1465_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1465_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5325), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16425));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1465_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1465_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1465_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1465_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_24 (.A0(d1[22]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[23]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16333), .COUT(n16334), .S0(d1_71__N_418[22]), 
          .S1(d1_71__N_418[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_37 (.A0(d2_adj_5741[70]), .B0(cout_adj_5345), 
          .C0(n81_adj_5115), .D0(d3_adj_5742[70]), .A1(d2_adj_5741[71]), 
          .B1(cout_adj_5345), .C1(n78_adj_5114), .D1(d3_adj_5742[71]), 
          .CIN(n16420), .S0(d3_71__N_562_adj_5758[70]), .S1(d3_71__N_562_adj_5758[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_37.INJECT1_1 = "NO";
    FD1P3AX phase_inc_carrGen_i0_i0 (.D(n323), .SP(clk_80mhz_enable_1470), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i0.GSR = "ENABLED";
    CCU2C _add_1_1519_add_4_37 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n81_adj_5290), .D0(d1[70]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n78_adj_5289), .D1(d1[71]), .CIN(n16197), .S0(d1_71__N_418[70]), 
          .S1(d1_71__N_418[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_35 (.A0(d2_adj_5741[68]), .B0(cout_adj_5345), 
          .C0(n87_adj_5117), .D0(d3_adj_5742[68]), .A1(d2_adj_5741[69]), 
          .B1(cout_adj_5345), .C1(n84_adj_5116), .D1(d3_adj_5742[69]), 
          .CIN(n16419), .COUT(n16420), .S0(d3_71__N_562_adj_5758[68]), 
          .S1(d3_71__N_562_adj_5758[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_33 (.A0(d2_adj_5741[66]), .B0(cout_adj_5345), 
          .C0(n93_adj_5119), .D0(d3_adj_5742[66]), .A1(d2_adj_5741[67]), 
          .B1(cout_adj_5345), .C1(n90_adj_5118), .D1(d3_adj_5742[67]), 
          .CIN(n16418), .COUT(n16419), .S0(d3_71__N_562_adj_5758[66]), 
          .S1(d3_71__N_562_adj_5758[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_31 (.A0(d2_adj_5741[64]), .B0(cout_adj_5345), 
          .C0(n99_adj_5121), .D0(d3_adj_5742[64]), .A1(d2_adj_5741[65]), 
          .B1(cout_adj_5345), .C1(n96_adj_5120), .D1(d3_adj_5742[65]), 
          .CIN(n16417), .COUT(n16418), .S0(d3_71__N_562_adj_5758[64]), 
          .S1(d3_71__N_562_adj_5758[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_31.INJECT1_1 = "NO";
    LUT4 mux_750_i22_3_lut (.A(led_c_2), .B(led_c_4), .C(n2824), .Z(n3657)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_750_i22_3_lut.init = 16'h3a3a;
    CCU2C _add_1_1406_add_4_22 (.A0(d1[20]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[21]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16332), .COUT(n16333), .S0(d1_71__N_418[20]), 
          .S1(d1_71__N_418[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_22.INJECT1_1 = "NO";
    CCU2C add_3827_3 (.A0(d_out_d_11__N_1892[17]), .B0(n931), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1890[17]), .B1(n930), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16579), .COUT(n16580));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3827_3.INIT0 = 16'h9995;
    defparam add_3827_3.INIT1 = 16'h9995;
    defparam add_3827_3.INJECT1_0 = "NO";
    defparam add_3827_3.INJECT1_1 = "NO";
    LUT4 mux_325_i52_4_lut (.A(n12156), .B(n166), .C(n17925), .D(n2572), 
         .Z(n2320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i52_4_lut.init = 16'hcfca;
    CCU2C _add_1_1633_add_4_38 (.A0(d_d6_adj_5746[71]), .B0(d6_adj_5745[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16358), .S0(n78_adj_4916));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1633_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_29 (.A0(d2_adj_5741[62]), .B0(cout_adj_5345), 
          .C0(n105_adj_5123), .D0(d3_adj_5742[62]), .A1(d2_adj_5741[63]), 
          .B1(cout_adj_5345), .C1(n102_adj_5122), .D1(d3_adj_5742[63]), 
          .CIN(n16416), .COUT(n16417), .S0(d3_71__N_562_adj_5758[62]), 
          .S1(d3_71__N_562_adj_5758[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_20 (.A0(d1[18]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[19]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16331), .COUT(n16332), .S0(d1_71__N_418[18]), 
          .S1(d1_71__N_418[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_27 (.A0(d2_adj_5741[60]), .B0(cout_adj_5345), 
          .C0(n111_adj_5125), .D0(d3_adj_5742[60]), .A1(d2_adj_5741[61]), 
          .B1(cout_adj_5345), .C1(n108_adj_5124), .D1(d3_adj_5742[61]), 
          .CIN(n16415), .COUT(n16416), .S0(d3_71__N_562_adj_5758[60]), 
          .S1(d3_71__N_562_adj_5758[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_36 (.A0(d_d6_adj_5746[69]), .B0(d6_adj_5745[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[70]), .B1(d6_adj_5745[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16357), .COUT(n16358), .S0(n84_adj_4918), 
          .S1(n81_adj_4917));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_25 (.A0(d2_adj_5741[58]), .B0(cout_adj_5345), 
          .C0(n117_adj_5127), .D0(d3_adj_5742[58]), .A1(d2_adj_5741[59]), 
          .B1(cout_adj_5345), .C1(n114_adj_5126), .D1(d3_adj_5742[59]), 
          .CIN(n16414), .COUT(n16415), .S0(d3_71__N_562_adj_5758[58]), 
          .S1(d3_71__N_562_adj_5758[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_34 (.A0(d_d6_adj_5746[67]), .B0(d6_adj_5745[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[68]), .B1(d6_adj_5745[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16356), .COUT(n16357), .S0(n90_adj_4920), 
          .S1(n87_adj_4919));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_23 (.A0(d2_adj_5741[56]), .B0(cout_adj_5345), 
          .C0(n123_adj_5129), .D0(d3_adj_5742[56]), .A1(d2_adj_5741[57]), 
          .B1(cout_adj_5345), .C1(n120_adj_5128), .D1(d3_adj_5742[57]), 
          .CIN(n16413), .COUT(n16414), .S0(d3_71__N_562_adj_5758[56]), 
          .S1(d3_71__N_562_adj_5758[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_21 (.A0(d2_adj_5741[54]), .B0(cout_adj_5345), 
          .C0(n129_adj_5131), .D0(d3_adj_5742[54]), .A1(d2_adj_5741[55]), 
          .B1(cout_adj_5345), .C1(n126_adj_5130), .D1(d3_adj_5742[55]), 
          .CIN(n16412), .COUT(n16413), .S0(d3_71__N_562_adj_5758[54]), 
          .S1(d3_71__N_562_adj_5758[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_19 (.A0(d2_adj_5741[52]), .B0(cout_adj_5345), 
          .C0(n135_adj_5133), .D0(d3_adj_5742[52]), .A1(d2_adj_5741[53]), 
          .B1(cout_adj_5345), .C1(n132_adj_5132), .D1(d3_adj_5742[53]), 
          .CIN(n16411), .COUT(n16412), .S0(d3_71__N_562_adj_5758[52]), 
          .S1(d3_71__N_562_adj_5758[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_19.INJECT1_1 = "NO";
    VLO i1 (.Z(GND_net));
    CCU2C _add_1_1498_add_4_17 (.A0(d2_adj_5741[50]), .B0(cout_adj_5345), 
          .C0(n141_adj_5135), .D0(d3_adj_5742[50]), .A1(d2_adj_5741[51]), 
          .B1(cout_adj_5345), .C1(n138_adj_5134), .D1(d3_adj_5742[51]), 
          .CIN(n16410), .COUT(n16411), .S0(d3_71__N_562_adj_5758[50]), 
          .S1(d3_71__N_562_adj_5758[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_35 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n87_adj_5292), .D0(d1[68]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n84_adj_5291), .D1(d1[69]), .CIN(n16196), .COUT(n16197), 
          .S0(d1_71__N_418[68]), .S1(d1_71__N_418[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_15 (.A0(d2_adj_5741[48]), .B0(cout_adj_5345), 
          .C0(n147_adj_5137), .D0(d3_adj_5742[48]), .A1(d2_adj_5741[49]), 
          .B1(cout_adj_5345), .C1(n144_adj_5136), .D1(d3_adj_5742[49]), 
          .CIN(n16409), .COUT(n16410), .S0(d3_71__N_562_adj_5758[48]), 
          .S1(d3_71__N_562_adj_5758[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_13 (.A0(d2_adj_5741[46]), .B0(cout_adj_5345), 
          .C0(n153_adj_5139), .D0(d3_adj_5742[46]), .A1(d2_adj_5741[47]), 
          .B1(cout_adj_5345), .C1(n150_adj_5138), .D1(d3_adj_5742[47]), 
          .CIN(n16408), .COUT(n16409), .S0(d3_71__N_562_adj_5758[46]), 
          .S1(d3_71__N_562_adj_5758[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1519_add_4_33 (.A0(MixerOutSin[11]), .B0(cout_adj_5534), 
          .C0(n93_adj_5294), .D0(d1[66]), .A1(MixerOutSin[11]), .B1(cout_adj_5534), 
          .C1(n90_adj_5293), .D1(d1[67]), .CIN(n16195), .COUT(n16196), 
          .S0(d1_71__N_418[66]), .S1(d1_71__N_418[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1519_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1519_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1519_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1519_add_4_33.INJECT1_1 = "NO";
    CCU2C add_3827_1 (.A0(ISquare[0]), .B0(GND_net), .C0(GND_net), .D0(ISquare[0]), 
          .A1(d_out_d_11__N_1892[17]), .B1(ISquare[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16579));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(68[15:27])
    defparam add_3827_1.INIT0 = 16'h000A;
    defparam add_3827_1.INIT1 = 16'h666a;
    defparam add_3827_1.INJECT1_0 = "NO";
    defparam add_3827_1.INJECT1_1 = "NO";
    LUT4 i5377_2_lut (.A(d3_adj_5742[0]), .B(d2_adj_5741[0]), .Z(d3_71__N_562_adj_5758[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5377_2_lut.init = 16'h6666;
    CCU2C _add_1_1498_add_4_11 (.A0(d2_adj_5741[44]), .B0(cout_adj_5345), 
          .C0(n159_adj_5141), .D0(d3_adj_5742[44]), .A1(d2_adj_5741[45]), 
          .B1(cout_adj_5345), .C1(n156_adj_5140), .D1(d3_adj_5742[45]), 
          .CIN(n16407), .COUT(n16408), .S0(d3_71__N_562_adj_5758[44]), 
          .S1(d3_71__N_562_adj_5758[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_9 (.A0(d2_adj_5741[42]), .B0(cout_adj_5345), 
          .C0(n165_adj_5143), .D0(d3_adj_5742[42]), .A1(d2_adj_5741[43]), 
          .B1(cout_adj_5345), .C1(n162_adj_5142), .D1(d3_adj_5742[43]), 
          .CIN(n16406), .COUT(n16407), .S0(d3_71__N_562_adj_5758[42]), 
          .S1(d3_71__N_562_adj_5758[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_18 (.A0(d1[16]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[17]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16330), .COUT(n16331), .S0(d1_71__N_418[16]), 
          .S1(d1_71__N_418[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_18.INJECT1_1 = "NO";
    CCU2C add_3825_15 (.A0(d_out_d_11__N_1875), .B0(d_out_d_11__N_1876[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1875), .B1(d_out_d_11__N_1876[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16577), .S0(n37_adj_5614), 
          .S1(d_out_d_11__N_1878[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3825_15.INIT0 = 16'h666a;
    defparam add_3825_15.INIT1 = 16'h666a;
    defparam add_3825_15.INJECT1_0 = "NO";
    defparam add_3825_15.INJECT1_1 = "NO";
    CCU2C add_3825_13 (.A0(d_out_d_11__N_1876[17]), .B0(n36_adj_5187), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n33_adj_5186), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16576), .COUT(n16577), .S0(n43), 
          .S1(n40));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3825_13.INIT0 = 16'h9995;
    defparam add_3825_13.INIT1 = 16'h9995;
    defparam add_3825_13.INJECT1_0 = "NO";
    defparam add_3825_13.INJECT1_1 = "NO";
    LUT4 mux_325_i49_4_lut (.A(n12152), .B(n175), .C(n17925), .D(n2572), 
         .Z(n2323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i49_4_lut.init = 16'hcfca;
    \CIC(WIDTH=72,DECIMATION_RATIO=4096)  CIC_cos_inst (.d_tmp({d_tmp_adj_5738}), 
            .clk_80mhz(clk_80mhz), .d5({d5_adj_5744}), .d_d_tmp({d_d_tmp_adj_5739}), 
            .d2({d2_adj_5741}), .d2_71__N_490({d2_71__N_490_adj_5757}), 
            .d3({d3_adj_5742}), .d3_71__N_562({d3_71__N_562_adj_5758}), 
            .d4({d4_adj_5743}), .d4_71__N_634({d4_71__N_634_adj_5759}), 
            .d5_71__N_706({d5_71__N_706_adj_5760}), .d6({d6_adj_5745}), 
            .d6_71__N_1459({d6_71__N_1459_adj_5772}), .d_d6({d_d6_adj_5746}), 
            .d7({d7_adj_5747}), .d7_71__N_1531({d7_71__N_1531_adj_5773}), 
            .d_d7({d_d7_adj_5748}), .d8({d8_adj_5749}), .d8_71__N_1603({d8_71__N_1603_adj_5774}), 
            .d_d8({d_d8_adj_5750}), .d9({d9_adj_5751}), .d9_71__N_1675({d9_71__N_1675_adj_5775}), 
            .d_d9({d_d9_adj_5752}), .n19(n19_adj_4696), .CIC1_outCos({CIC1_outCos}), 
            .d1({d1_adj_5740}), .d1_71__N_418({d1_71__N_418_adj_5756}), 
            .n22(n22), .n8(n8), .n37(n37_adj_4715), .n11(n11), .n10(n10), 
            .n13(n13), .count({count_adj_5755}), .n31(n31_adj_2808), .\CICGain[0] (CICGain[0]), 
            .n66(n66_adj_4798), .n18(n18_adj_4697), .n30(n30_adj_2809), 
            .n21(n21_adj_4694), .n3(n3_adj_4712), .n2(n2_adj_4713), .n5(n5_adj_4710), 
            .n4(n4_adj_4711), .n7(n7_adj_4708), .n6(n6_adj_4709), .n9(n9_adj_4706), 
            .n8_adj_127(n8_adj_4707), .n15(n15_adj_4700), .n14(n14_adj_4701), 
            .\CICGain[1] (CICGain[1]), .\d10[68] (d10_adj_5753[68]), .\d10[69] (d10_adj_5753[69]), 
            .\d10[67] (d10_adj_5753[67]), .n11_adj_128(n11_adj_4704), .n10_adj_129(n10_adj_4705), 
            .n13_adj_130(n13_adj_4702), .n12(n12_adj_4703), .n63(n63), 
            .n131(n131), .\d_out_11__N_1819[2] (d_out_11__N_1819[2]), .n64(n64), 
            .n132(n132_adj_4792), .\d_out_11__N_1819[3] (d_out_11__N_1819[3]), 
            .n65(n65), .n133(n133), .\d_out_11__N_1819[4] (d_out_11__N_1819[4]), 
            .n66_adj_131(n66), .n134(n134), .\d_out_11__N_1819[5] (d_out_11__N_1819[5]), 
            .\d10[66] (d10[66]), .n135(n135_adj_4793), .\d_out_11__N_1819[6] (d_out_11__N_1819[6]), 
            .n12_adj_132(n12), .\d10[67]_adj_133 (d10[67]), .n136(n136), 
            .\d_out_11__N_1819[7] (d_out_11__N_1819[7]), .n63_adj_134(n63_adj_4795), 
            .n131_adj_135(n131_adj_4799), .n15_adj_136(n15), .n64_adj_137(n64_adj_4796), 
            .n132_adj_138(n132_adj_4800), .n65_adj_139(n65_adj_4797), .n133_adj_140(n133_adj_4801), 
            .n134_adj_141(n134_adj_4802), .n135_adj_142(n135_adj_4803), 
            .n136_adj_143(n136_adj_4804), .n36(n36_adj_4716), .n25(n25_adj_4690), 
            .n24(n24_adj_4691), .n25_adj_144(n25_adj_2814), .n33(n33), 
            .n24_adj_145(n24_adj_2815), .n27(n27_adj_4688), .n27_adj_146(n27_adj_2812), 
            .n26(n26_adj_2813), .n32(n32), .n14_adj_147(n14), .n35(n35), 
            .\d10[60] (d10_adj_5753[60]), .n26_adj_148(n26_adj_4689), .n34(n34), 
            .n17(n17), .\d10[59] (d10_adj_5753[59]), .\d10[61] (d10_adj_5753[61]), 
            .\d10[62] (d10_adj_5753[62]), .\d10[63] (d10_adj_5753[63]), 
            .\d10[64] (d10_adj_5753[64]), .\d10[70] (d10_adj_5753[70]), 
            .\d10[71] (d10_adj_5753[71]), .\d_out_11__N_1819[10] (d_out_11__N_1819_adj_5778[10]), 
            .\d_out_11__N_1819[11] (d_out_11__N_1819_adj_5778[11]), .n20(n20_adj_4695), 
            .n29(n29_adj_4686), .n16(n16), .n37_adj_149(n37), .n29_adj_150(n29_adj_2810), 
            .n17610(n17610), .\d10[65] (d10[65]), .\d10[68]_adj_151 (d10[68]), 
            .n87_adj_252({n36_adj_5400, n39_adj_5401, n42_adj_5402, n45_adj_5403, 
            n48_adj_5404, n51_adj_5405, n54_adj_5406, n57_adj_5407, 
            n60_adj_5408, n63_adj_5409, n66_adj_5410, n69_adj_5411, 
            n72_adj_5412, n75_adj_5413, n78_adj_5414, n81_adj_5415}), 
            .n28(n28_adj_4687), .n31_adj_155(n31_adj_4683), .n17630(n17630), 
            .n19_adj_156(n19), .n28_adj_157(n28_adj_2811), .n18_adj_158(n18), 
            .n21_adj_159(n21), .n20_adj_160(n20), .n36_adj_161(n36), .n30_adj_162(n30_adj_4685), 
            .n37_adj_163(n37_adj_4677), .n36_adj_164(n36_adj_4678), .n3_adj_165(n3_adj_4674), 
            .n2_adj_166(n2_adj_4675), .n5_adj_167(n5_adj_4672), .n4_adj_168(n4_adj_4673), 
            .n7_adj_169(n7_adj_4670), .n6_adj_170(n6_adj_4671), .n9_adj_171(n9_adj_4668), 
            .n8_adj_172(n8_adj_4669), .n11_adj_173(n11_adj_4666), .n10_adj_174(n10_adj_4667), 
            .n35_adj_175(n35_adj_4679), .n13_adj_176(n13_adj_4664), .n12_adj_177(n12_adj_4665), 
            .n15_adj_178(n15_adj_4662), .n14_adj_179(n14_adj_4663), .n17_adj_180(n17_adj_4660), 
            .n34_adj_181(n34_adj_4680), .n16_adj_182(n16_adj_4661), .n19_adj_183(n19_adj_4658), 
            .n18_adj_184(n18_adj_4659), .n21_adj_185(n21_adj_4656), .n20_adj_186(n20_adj_4657), 
            .n23(n23_adj_4654), .n22_adj_187(n22_adj_4655), .n23_adj_188(n23), 
            .n25_adj_189(n25_adj_4652), .n24_adj_190(n24_adj_4653), .n27_adj_191(n27_adj_4649), 
            .n26_adj_192(n26_adj_4650), .n29_adj_193(n29_adj_4647), .n28_adj_194(n28_adj_4648), 
            .n3_adj_195(n3), .n2_adj_196(n2), .n5_adj_197(n5), .n31_adj_198(n31_adj_4645), 
            .n4_adj_199(n4), .n7_adj_200(n7), .n6_adj_201(n6), .n9_adj_202(n9_adj_4741), 
            .n8_adj_203(n8_adj_4745), .n30_adj_204(n30_adj_4646), .n33_adj_205(n33_adj_4643), 
            .n32_adj_206(n32_adj_4644), .n35_adj_207(n35_adj_4641), .n34_adj_208(n34_adj_4642), 
            .n37_adj_209(n37_adj_4639), .n36_adj_210(n36_adj_4640), .n17_adj_211(n17_adj_4698), 
            .n16_adj_212(n16_adj_4699), .n11_adj_213(n11_adj_4743), .n10_adj_214(n10_adj_4742), 
            .n13_adj_215(n13_adj_4740), .n12_adj_216(n12_adj_4744), .n15_adj_217(n15_adj_4738), 
            .n14_adj_218(n14_adj_4739), .n17_adj_219(n17_adj_4736), .n16_adj_220(n16_adj_4737), 
            .n19_adj_221(n19_adj_4734), .n18_adj_222(n18_adj_4735), .n21_adj_223(n21_adj_4732), 
            .n23_adj_224(n23_adj_4692), .n22_adj_225(n22_adj_4693), .n20_adj_226(n20_adj_4733), 
            .n23_adj_227(n23_adj_4730), .n22_adj_228(n22_adj_4731), .n25_adj_229(n25_adj_4728), 
            .n24_adj_230(n24_adj_4729), .n27_adj_231(n27_adj_4726), .n26_adj_232(n26_adj_4727), 
            .n29_adj_233(n29_adj_4724), .\d_out_11__N_1819[8] (d_out_11__N_1819[8]), 
            .n28_adj_234(n28_adj_4725), .n31_adj_235(n31_adj_4722), .n30_adj_236(n30_adj_4723), 
            .n118(n118_adj_5630), .n120(n120_adj_5038), .cout(cout_adj_5516), 
            .n115(n115_adj_5629), .n117(n117_adj_5037), .n112(n112_adj_5628), 
            .n114(n114_adj_5036), .n109(n109_adj_5627), .n111(n111_adj_5035), 
            .n33_adj_237(n33_adj_4720), .n32_adj_238(n32_adj_4721), .n106(n106_adj_5626), 
            .n108(n108_adj_5034), .n103(n103_adj_5625), .n105(n105_adj_5033), 
            .n100(n100_adj_5624), .n102(n102_adj_5032), .n97(n97_adj_5623), 
            .n99(n99_adj_5031), .n94(n94_adj_5622), .n96(n96_adj_5030), 
            .n91(n91_adj_5621), .n93(n93_adj_5029), .n88(n88_adj_5620), 
            .n90(n90_adj_5028), .n35_adj_239(n35_adj_4718), .n85(n85_adj_5619), 
            .n87(n87_adj_5027), .n82(n82_adj_5618), .n84(n84_adj_5026), 
            .n79(n79_adj_5617), .n81_adj_240(n81_adj_5025), .n76(n76_adj_5616), 
            .n78_adj_241(n78_adj_5024), .n34_adj_242(n34_adj_4719), .n33_adj_243(n33_adj_4681), 
            .n32_adj_244(n32_adj_4682), .n3_adj_245(n3_adj_2820), .n2_adj_246(n2_adj_2821), 
            .n5_adj_247(n5_adj_2818), .n4_adj_248(n4_adj_2819), .n7_adj_249(n7_adj_2816), 
            .n6_adj_250(n6_adj_2817), .n9_adj_251(n9)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(148[4] 154[5])
    CCU2C _add_1_1636_add_4_10 (.A0(d_d7_adj_5748[43]), .B0(d7_adj_5747[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[44]), .B1(d7_adj_5747[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16121), .COUT(n16122), .S0(n162_adj_4980), 
          .S1(n159_adj_4979));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_10.INJECT1_1 = "NO";
    LUT4 mux_325_i50_4_lut (.A(n27_adj_5727), .B(n172), .C(n17925), .D(n2388), 
         .Z(n2322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i50_4_lut.init = 16'hcfca;
    CCU2C _add_1_1636_add_4_6 (.A0(d_d7_adj_5748[39]), .B0(d7_adj_5747[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[40]), .B1(d7_adj_5747[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16119), .COUT(n16120), .S0(n174_adj_4984), 
          .S1(n171_adj_4983));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1636_add_4_8 (.A0(d_d7_adj_5748[41]), .B0(d7_adj_5747[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d7_adj_5748[42]), .B1(d7_adj_5747[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16120), .COUT(n16121), .S0(n168_adj_4982), 
          .S1(n165_adj_4981));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam _add_1_1636_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1636_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1636_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1636_add_4_8.INJECT1_1 = "NO";
    LUT4 i3232_2_lut (.A(n166_adj_5643), .B(led_c_3), .Z(n2388)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i3232_2_lut.init = 16'h8888;
    CCU2C _add_1_1633_add_4_32 (.A0(d_d6_adj_5746[65]), .B0(d6_adj_5745[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[66]), .B1(d6_adj_5745[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16355), .COUT(n16356), .S0(n96_adj_4922), 
          .S1(n93_adj_4921));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_32.INJECT1_1 = "NO";
    CCU2C add_3825_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1876[17]), .C0(n42), 
          .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n39), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16575), .COUT(n16576), .S0(n49), .S1(n46));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3825_11.INIT0 = 16'h6969;
    defparam add_3825_11.INIT1 = 16'h9995;
    defparam add_3825_11.INJECT1_0 = "NO";
    defparam add_3825_11.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_30 (.A0(d_d6_adj_5746[63]), .B0(d6_adj_5745[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[64]), .B1(d6_adj_5745[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16354), .COUT(n16355), .S0(n102_adj_4924), 
          .S1(n99_adj_4923));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_30.INJECT1_1 = "NO";
    CCU2C add_3825_9 (.A0(ISquare[31]), .B0(d_out_d_11__N_1876[17]), .C0(n48), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1876[17]), 
          .C1(n45), .D1(VCC_net), .CIN(n16574), .COUT(n16575), .S0(n55), 
          .S1(n52));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3825_9.INIT0 = 16'h6969;
    defparam add_3825_9.INIT1 = 16'h6969;
    defparam add_3825_9.INJECT1_0 = "NO";
    defparam add_3825_9.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_28 (.A0(d_d6_adj_5746[61]), .B0(d6_adj_5745[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[62]), .B1(d6_adj_5745[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16353), .COUT(n16354), .S0(n108_adj_4926), 
          .S1(n105_adj_4925));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_28.INJECT1_1 = "NO";
    CCU2C add_3825_7 (.A0(d_out_d_11__N_1876[17]), .B0(n17938), .C0(n54), 
          .D0(VCC_net), .A1(d_out_d_11__N_1876[17]), .B1(n51), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16573), .COUT(n16574), .S0(n61), .S1(n58));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3825_7.INIT0 = 16'h6969;
    defparam add_3825_7.INIT1 = 16'h9995;
    defparam add_3825_7.INJECT1_0 = "NO";
    defparam add_3825_7.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_26 (.A0(d_d6_adj_5746[59]), .B0(d6_adj_5745[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[60]), .B1(d6_adj_5745[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16352), .COUT(n16353), .S0(n114_adj_4928), 
          .S1(n111_adj_4927));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_26.INJECT1_1 = "NO";
    CCU2C add_3825_5 (.A0(n60), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1874[17]), .B1(d_out_d_11__N_1876[17]), .C1(n57), 
          .D1(VCC_net), .CIN(n16572), .COUT(n16573), .S0(n67), .S1(n64_adj_5615));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3825_5.INIT0 = 16'haaa0;
    defparam add_3825_5.INIT1 = 16'h9696;
    defparam add_3825_5.INJECT1_0 = "NO";
    defparam add_3825_5.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_24 (.A0(d_d6_adj_5746[57]), .B0(d6_adj_5745[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[58]), .B1(d6_adj_5745[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16351), .COUT(n16352), .S0(n120_adj_4930), 
          .S1(n117_adj_4929));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_24.INJECT1_1 = "NO";
    CCU2C add_3825_3 (.A0(d_out_d_11__N_1876[17]), .B0(ISquare[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16571), .COUT(n16572), .S1(n70));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3825_3.INIT0 = 16'h666a;
    defparam add_3825_3.INIT1 = 16'h555f;
    defparam add_3825_3.INJECT1_0 = "NO";
    defparam add_3825_3.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_22 (.A0(d_d6_adj_5746[55]), .B0(d6_adj_5745[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[56]), .B1(d6_adj_5745[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16350), .COUT(n16351), .S0(n126_adj_4932), 
          .S1(n123_adj_4931));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_22.INJECT1_1 = "NO";
    CCU2C add_3825_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1876[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16571));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3825_1.INIT0 = 16'h0000;
    defparam add_3825_1.INIT1 = 16'haaaf;
    defparam add_3825_1.INJECT1_0 = "NO";
    defparam add_3825_1.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_20 (.A0(d_d6_adj_5746[53]), .B0(d6_adj_5745[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[54]), .B1(d6_adj_5745[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16349), .COUT(n16350), .S0(n132_adj_4934), 
          .S1(n129_adj_4933));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_18 (.A0(d_d6_adj_5746[51]), .B0(d6_adj_5745[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[52]), .B1(d6_adj_5745[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16348), .COUT(n16349), .S0(n138_adj_4936), 
          .S1(n135_adj_4935));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_16 (.A0(d_d6_adj_5746[49]), .B0(d6_adj_5745[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[50]), .B1(d6_adj_5745[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16347), .COUT(n16348), .S0(n144_adj_4938), 
          .S1(n141_adj_4937));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_16.INJECT1_1 = "NO";
    CCU2C add_3835_19 (.A0(d_out_d_11__N_1879), .B0(d_out_d_11__N_1880[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_out_d_11__N_1879), .B1(d_out_d_11__N_1880[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16565), .S0(n45_adj_5346), 
          .S1(d_out_d_11__N_1882[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3835_19.INIT0 = 16'h666a;
    defparam add_3835_19.INIT1 = 16'h666a;
    defparam add_3835_19.INJECT1_0 = "NO";
    defparam add_3835_19.INJECT1_1 = "NO";
    CCU2C add_3835_17 (.A0(d_out_d_11__N_1880[17]), .B0(n44), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n41), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16564), .COUT(n16565), .S0(n51_adj_5348), 
          .S1(n48_adj_5347));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3835_17.INIT0 = 16'h9995;
    defparam add_3835_17.INIT1 = 16'h9995;
    defparam add_3835_17.INJECT1_0 = "NO";
    defparam add_3835_17.INJECT1_1 = "NO";
    GSR GSR_INST (.GSR(VCC_net));
    FD1P3AX phase_inc_carrGen_i0_i1 (.D(n320), .SP(clk_80mhz_enable_1471), 
            .CK(clk_80mhz), .Q(phase_inc_carrGen[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam phase_inc_carrGen_i0_i1.GSR = "ENABLED";
    LUT4 mux_325_i47_4_lut (.A(n12148), .B(n181), .C(n17925), .D(n2572), 
         .Z(n2325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i47_4_lut.init = 16'hcfca;
    LUT4 mux_325_i48_4_lut (.A(n12150), .B(n178), .C(n17925), .D(n2572), 
         .Z(n2324)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i48_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1498_add_4_7 (.A0(d2_adj_5741[40]), .B0(cout_adj_5345), 
          .C0(n171_adj_5145), .D0(d3_adj_5742[40]), .A1(d2_adj_5741[41]), 
          .B1(cout_adj_5345), .C1(n168_adj_5144), .D1(d3_adj_5742[41]), 
          .CIN(n16405), .COUT(n16406), .S0(d3_71__N_562_adj_5758[40]), 
          .S1(d3_71__N_562_adj_5758[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1498_add_4_5 (.A0(d2_adj_5741[38]), .B0(cout_adj_5345), 
          .C0(n177_adj_5147), .D0(d3_adj_5742[38]), .A1(d2_adj_5741[39]), 
          .B1(cout_adj_5345), .C1(n174_adj_5146), .D1(d3_adj_5742[39]), 
          .CIN(n16404), .COUT(n16405), .S0(d3_71__N_562_adj_5758[38]), 
          .S1(d3_71__N_562_adj_5758[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_5.INJECT1_1 = "NO";
    LUT4 i3085_4_lut (.A(n27_adj_5727), .B(n187), .C(n17925), .D(n2393), 
         .Z(n2327)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i3085_4_lut.init = 16'hc5c0;
    CCU2C _add_1_1498_add_4_3 (.A0(d2_adj_5741[36]), .B0(cout_adj_5345), 
          .C0(n183_adj_5149), .D0(d3_adj_5742[36]), .A1(d2_adj_5741[37]), 
          .B1(cout_adj_5345), .C1(n180_adj_5148), .D1(d3_adj_5742[37]), 
          .CIN(n16403), .COUT(n16404), .S0(d3_71__N_562_adj_5758[36]), 
          .S1(d3_71__N_562_adj_5758[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1498_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1498_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_3.INJECT1_1 = "NO";
    LUT4 mux_325_i46_4_lut (.A(n12146), .B(n184), .C(n17925), .D(n2572), 
         .Z(n2326)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i46_4_lut.init = 16'hc0ca;
    LUT4 mux_325_i43_4_lut (.A(n12142), .B(n193), .C(n17925), .D(n2572), 
         .Z(n2329)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i43_4_lut.init = 16'hc0ca;
    LUT4 i2296_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(led_c_3), .D(n265_adj_5676), 
         .Z(n12094)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2296_3_lut_4_lut.init = 16'hf404;
    LUT4 i5372_2_lut (.A(d4_adj_5743[0]), .B(d3_adj_5742[0]), .Z(d4_71__N_634_adj_5759[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5372_2_lut.init = 16'h6666;
    LUT4 i5369_2_lut (.A(d5_adj_5744[0]), .B(d4_adj_5743[0]), .Z(d5_71__N_706_adj_5760[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5369_2_lut.init = 16'h6666;
    LUT4 mux_325_i44_4_lut (.A(n12144), .B(n190), .C(n17925), .D(n2572), 
         .Z(n2328)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i44_4_lut.init = 16'hc0ca;
    LUT4 i26_4_lut_adj_62 (.A(n2572), .B(n199), .C(n17925), .D(n13_adj_5726), 
         .Z(n11_adj_5725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i26_4_lut_adj_62.init = 16'hcacf;
    LUT4 i2482_4_lut (.A(n196), .B(n190_adj_5651), .C(led_c_3), .D(n17932), 
         .Z(n12296)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2482_4_lut.init = 16'hcac0;
    CCU2C _add_1_1498_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5345), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16403));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(64[15:24])
    defparam _add_1_1498_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1498_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1498_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1498_add_4_1.INJECT1_1 = "NO";
    LUT4 mux_325_i39_4_lut (.A(n12136), .B(n205), .C(n17925), .D(n2572), 
         .Z(n2333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i39_4_lut.init = 16'hcfca;
    LUT4 mux_325_i40_4_lut (.A(n12138), .B(n202), .C(n17925), .D(n2572), 
         .Z(n2332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i40_4_lut.init = 16'hcfca;
    LUT4 mux_325_i37_4_lut (.A(n12132), .B(n211), .C(n17925), .D(n2572), 
         .Z(n2335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i37_4_lut.init = 16'hcfca;
    LUT4 i1_2_lut_rep_179 (.A(led_c_1), .B(led_c_4), .Z(n17951)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(186[11] 212[6])
    defparam i1_2_lut_rep_179.init = 16'h2222;
    LUT4 mux_325_i38_4_lut (.A(n12134), .B(n208), .C(n17925), .D(n2572), 
         .Z(n2334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i38_4_lut.init = 16'hcfca;
    LUT4 i3145_2_lut (.A(led_c_4), .B(n2824), .Z(n3678)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i3145_2_lut.init = 16'hbbbb;
    LUT4 mux_325_i35_4_lut (.A(n12128), .B(n217), .C(n17925), .D(n2572), 
         .Z(n2337)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i35_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1471_add_4_37 (.A0(d8_adj_5749[70]), .B0(cout_adj_5517), 
          .C0(n81_adj_4989), .D0(n3_adj_4674), .A1(d8_adj_5749[71]), .B1(cout_adj_5517), 
          .C1(n78_adj_4988), .D1(n2_adj_4675), .CIN(n16398), .S0(d9_71__N_1675_adj_5775[70]), 
          .S1(d9_71__N_1675_adj_5775[71]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_35 (.A0(d8_adj_5749[68]), .B0(cout_adj_5517), 
          .C0(n87_adj_4991), .D0(n5_adj_4672), .A1(d8_adj_5749[69]), .B1(cout_adj_5517), 
          .C1(n84_adj_4990), .D1(n4_adj_4673), .CIN(n16397), .COUT(n16398), 
          .S0(d9_71__N_1675_adj_5775[68]), .S1(d9_71__N_1675_adj_5775[69]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_33 (.A0(d8_adj_5749[66]), .B0(cout_adj_5517), 
          .C0(n93_adj_4993), .D0(n7_adj_4670), .A1(d8_adj_5749[67]), .B1(cout_adj_5517), 
          .C1(n90_adj_4992), .D1(n6_adj_4671), .CIN(n16396), .COUT(n16397), 
          .S0(d9_71__N_1675_adj_5775[66]), .S1(d9_71__N_1675_adj_5775[67]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_33.INJECT1_1 = "NO";
    nco_sig nco_sig_inst (.\phase_accum[63] (phase_accum[63]), .sinGen_c(sinGen_c)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(114[4] 120[5])
    CCU2C _add_1_1627_add_4_34 (.A0(d_d9[31]), .B0(d9[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d9[32]), .B1(d9[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16292), .COUT(n16293));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam _add_1_1627_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1627_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1627_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1627_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_31 (.A0(d8_adj_5749[64]), .B0(cout_adj_5517), 
          .C0(n99_adj_4995), .D0(n9_adj_4668), .A1(d8_adj_5749[65]), .B1(cout_adj_5517), 
          .C1(n96_adj_4994), .D1(n8_adj_4669), .CIN(n16395), .COUT(n16396), 
          .S0(d9_71__N_1675_adj_5775[64]), .S1(d9_71__N_1675_adj_5775[65]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_31.INJECT1_1 = "NO";
    LUT4 i2374_3_lut_4_lut (.A(n18075), .B(n17937), .C(n18076), .D(n133_adj_5632), 
         .Z(n12172)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2374_3_lut_4_lut.init = 16'hfb0b;
    CCU2C _add_1_1471_add_4_29 (.A0(d8_adj_5749[62]), .B0(cout_adj_5517), 
          .C0(n105_adj_4997), .D0(n11_adj_4666), .A1(d8_adj_5749[63]), 
          .B1(cout_adj_5517), .C1(n102_adj_4996), .D1(n10_adj_4667), .CIN(n16394), 
          .COUT(n16395), .S0(d9_71__N_1675_adj_5775[62]), .S1(d9_71__N_1675_adj_5775[63]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_29.INJECT1_1 = "NO";
    PFUMX i6419 (.BLUT(n17959), .ALUT(n17960), .C0(n17069), .Z(n17961));
    CCU2C _add_1_1471_add_4_27 (.A0(d8_adj_5749[60]), .B0(cout_adj_5517), 
          .C0(n111_adj_4999), .D0(n13_adj_4664), .A1(d8_adj_5749[61]), 
          .B1(cout_adj_5517), .C1(n108_adj_4998), .D1(n12_adj_4665), .CIN(n16393), 
          .COUT(n16394), .S0(d9_71__N_1675_adj_5775[60]), .S1(d9_71__N_1675_adj_5775[61]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_25 (.A0(d8_adj_5749[58]), .B0(cout_adj_5517), 
          .C0(n117_adj_5001), .D0(n15_adj_4662), .A1(d8_adj_5749[59]), 
          .B1(cout_adj_5517), .C1(n114_adj_5000), .D1(n14_adj_4663), .CIN(n16392), 
          .COUT(n16393), .S0(d9_71__N_1675_adj_5775[58]), .S1(d9_71__N_1675_adj_5775[59]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_23 (.A0(d8_adj_5749[56]), .B0(cout_adj_5517), 
          .C0(n123_adj_5003), .D0(n17_adj_4660), .A1(d8_adj_5749[57]), 
          .B1(cout_adj_5517), .C1(n120_adj_5002), .D1(n16_adj_4661), .CIN(n16391), 
          .COUT(n16392), .S0(d9_71__N_1675_adj_5775[56]), .S1(d9_71__N_1675_adj_5775[57]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_21 (.A0(d8_adj_5749[54]), .B0(cout_adj_5517), 
          .C0(n129_adj_5005), .D0(n19_adj_4658), .A1(d8_adj_5749[55]), 
          .B1(cout_adj_5517), .C1(n126_adj_5004), .D1(n18_adj_4659), .CIN(n16390), 
          .COUT(n16391), .S0(d9_71__N_1675_adj_5775[54]), .S1(d9_71__N_1675_adj_5775[55]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_19 (.A0(d8_adj_5749[52]), .B0(cout_adj_5517), 
          .C0(n135_adj_5007), .D0(n21_adj_4656), .A1(d8_adj_5749[53]), 
          .B1(cout_adj_5517), .C1(n132_adj_5006), .D1(n20_adj_4657), .CIN(n16389), 
          .COUT(n16390), .S0(d9_71__N_1675_adj_5775[52]), .S1(d9_71__N_1675_adj_5775[53]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_19.INJECT1_1 = "NO";
    LUT4 mux_325_i36_4_lut (.A(n12130), .B(n214), .C(n17925), .D(n2572), 
         .Z(n2336)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam mux_325_i36_4_lut.init = 16'hc0ca;
    LUT4 i2370_3_lut_4_lut (.A(led_c_2), .B(n17937), .C(led_c_3), .D(n139_adj_5634), 
         .Z(n12168)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(191[7] 211[11])
    defparam i2370_3_lut_4_lut.init = 16'hfb0b;
    CCU2C _add_1_1633_add_4_14 (.A0(d_d6_adj_5746[47]), .B0(d6_adj_5745[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[48]), .B1(d6_adj_5745[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16346), .COUT(n16347), .S0(n150_adj_4940), 
          .S1(n147_adj_4939));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_17 (.A0(d8_adj_5749[50]), .B0(cout_adj_5517), 
          .C0(n141_adj_5009), .D0(n23_adj_4654), .A1(d8_adj_5749[51]), 
          .B1(cout_adj_5517), .C1(n138_adj_5008), .D1(n22_adj_4655), .CIN(n16388), 
          .COUT(n16389), .S0(d9_71__N_1675_adj_5775[50]), .S1(d9_71__N_1675_adj_5775[51]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_12 (.A0(d_d6_adj_5746[45]), .B0(d6_adj_5745[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[46]), .B1(d6_adj_5745[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16345), .COUT(n16346), .S0(n156_adj_4942), 
          .S1(n153_adj_4941));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_15 (.A0(d8_adj_5749[48]), .B0(cout_adj_5517), 
          .C0(n147_adj_5011), .D0(n25_adj_4652), .A1(d8_adj_5749[49]), 
          .B1(cout_adj_5517), .C1(n144_adj_5010), .D1(n24_adj_4653), .CIN(n16387), 
          .COUT(n16388), .S0(d9_71__N_1675_adj_5775[48]), .S1(d9_71__N_1675_adj_5775[49]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_10 (.A0(d_d6_adj_5746[43]), .B0(d6_adj_5745[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[44]), .B1(d6_adj_5745[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16344), .COUT(n16345), .S0(n162_adj_4944), 
          .S1(n159_adj_4943));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_13 (.A0(d8_adj_5749[46]), .B0(cout_adj_5517), 
          .C0(n153_adj_5013), .D0(n27_adj_4649), .A1(d8_adj_5749[47]), 
          .B1(cout_adj_5517), .C1(n150_adj_5012), .D1(n26_adj_4650), .CIN(n16386), 
          .COUT(n16387), .S0(d9_71__N_1675_adj_5775[46]), .S1(d9_71__N_1675_adj_5775[47]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_8 (.A0(d_d6_adj_5746[41]), .B0(d6_adj_5745[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[42]), .B1(d6_adj_5745[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16343), .COUT(n16344), .S0(n168_adj_4946), 
          .S1(n165_adj_4945));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_11 (.A0(d8_adj_5749[44]), .B0(cout_adj_5517), 
          .C0(n159_adj_5015), .D0(n29_adj_4647), .A1(d8_adj_5749[45]), 
          .B1(cout_adj_5517), .C1(n156_adj_5014), .D1(n28_adj_4648), .CIN(n16385), 
          .COUT(n16386), .S0(d9_71__N_1675_adj_5775[44]), .S1(d9_71__N_1675_adj_5775[45]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_6 (.A0(d_d6_adj_5746[39]), .B0(d6_adj_5745[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[40]), .B1(d6_adj_5745[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16342), .COUT(n16343), .S0(n174_adj_4948), 
          .S1(n171_adj_4947));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_9 (.A0(d8_adj_5749[42]), .B0(cout_adj_5517), 
          .C0(n165_adj_5017), .D0(n31_adj_4645), .A1(d8_adj_5749[43]), 
          .B1(cout_adj_5517), .C1(n162_adj_5016), .D1(n30_adj_4646), .CIN(n16384), 
          .COUT(n16385), .S0(d9_71__N_1675_adj_5775[42]), .S1(d9_71__N_1675_adj_5775[43]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_4 (.A0(d_d6_adj_5746[37]), .B0(d6_adj_5745[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(d_d6_adj_5746[38]), .B1(d6_adj_5745[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16341), .COUT(n16342), .S0(n180_adj_4950), 
          .S1(n177_adj_4949));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1633_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_7 (.A0(d8_adj_5749[40]), .B0(cout_adj_5517), 
          .C0(n171_adj_5019), .D0(n33_adj_4643), .A1(d8_adj_5749[41]), 
          .B1(cout_adj_5517), .C1(n168_adj_5018), .D1(n32_adj_4644), .CIN(n16383), 
          .COUT(n16384), .S0(d9_71__N_1675_adj_5775[40]), .S1(d9_71__N_1675_adj_5775[41]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1633_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_d6_adj_5746[36]), .B1(d6_adj_5745[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n16341), .S1(n183_adj_4951));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam _add_1_1633_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1633_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1633_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1633_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_5 (.A0(d8_adj_5749[38]), .B0(cout_adj_5517), 
          .C0(n177_adj_5021), .D0(n35_adj_4641), .A1(d8_adj_5749[39]), 
          .B1(cout_adj_5517), .C1(n174_adj_5020), .D1(n34_adj_4642), .CIN(n16382), 
          .COUT(n16383), .S0(d9_71__N_1675_adj_5775[38]), .S1(d9_71__N_1675_adj_5775[39]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut (.A(led_c_3), .B(led_c_0), .C(led_c_4), 
         .D(led_c_1), .Z(n17090)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(199[11] 210[18])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0800;
    CCU2C _add_1_1471_add_4_3 (.A0(d8_adj_5749[36]), .B0(cout_adj_5517), 
          .C0(n183_adj_5023), .D0(n37_adj_4639), .A1(d8_adj_5749[37]), 
          .B1(cout_adj_5517), .C1(n180_adj_5022), .D1(n36_adj_4640), .CIN(n16381), 
          .COUT(n16382), .S0(d9_71__N_1675_adj_5775[36]), .S1(d9_71__N_1675_adj_5775[37]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1471_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1471_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_3.INJECT1_1 = "NO";
    CCU2C add_3835_15 (.A0(d_out_d_11__N_1880[17]), .B0(n50), .C0(GND_net), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n47), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16563), .COUT(n16564), .S0(n57_adj_5350), 
          .S1(n54_adj_5349));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3835_15.INIT0 = 16'h9995;
    defparam add_3835_15.INIT1 = 16'h9995;
    defparam add_3835_15.INJECT1_0 = "NO";
    defparam add_3835_15.INJECT1_1 = "NO";
    CCU2C _add_1_1471_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5517), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16381));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam _add_1_1471_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1471_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1471_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1471_add_4_1.INJECT1_1 = "NO";
    CCU2C add_3835_13 (.A0(ISquare[31]), .B0(d_out_d_11__N_1880[17]), .C0(n56), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n53), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16562), .COUT(n16563), .S0(n63_adj_5352), 
          .S1(n60_adj_5351));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3835_13.INIT0 = 16'h6969;
    defparam add_3835_13.INIT1 = 16'h9995;
    defparam add_3835_13.INJECT1_0 = "NO";
    defparam add_3835_13.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16377), .S0(cout_adj_5326));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1421_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1421_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_36 (.A0(d5[34]), .B0(d4[34]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[35]), .B1(d4[35]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16376), .COUT(n16377), .S0(d5_71__N_706[34]), .S1(d5_71__N_706[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_36.INJECT1_1 = "NO";
    CCU2C add_3835_11 (.A0(ISquare[31]), .B0(d_out_d_11__N_1880[17]), .C0(n62), 
          .D0(VCC_net), .A1(ISquare[31]), .B1(d_out_d_11__N_1880[17]), 
          .C1(n59), .D1(VCC_net), .CIN(n16561), .COUT(n16562), .S0(n69_adj_5354), 
          .S1(n66_adj_5353));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3835_11.INIT0 = 16'h6969;
    defparam add_3835_11.INIT1 = 16'h6969;
    defparam add_3835_11.INJECT1_0 = "NO";
    defparam add_3835_11.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_34 (.A0(d5[32]), .B0(d4[32]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[33]), .B1(d4[33]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16375), .COUT(n16376), .S0(d5_71__N_706[32]), .S1(d5_71__N_706[33]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_32 (.A0(d5[30]), .B0(d4[30]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[31]), .B1(d4[31]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16374), .COUT(n16375), .S0(d5_71__N_706[30]), .S1(d5_71__N_706[31]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_32.INJECT1_1 = "NO";
    CCU2C add_3835_9 (.A0(d_out_d_11__N_1880[17]), .B0(n17938), .C0(n68), 
          .D0(VCC_net), .A1(d_out_d_11__N_1880[17]), .B1(n65_adj_5604), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16560), .COUT(n16561), .S0(n75_adj_5356), 
          .S1(n72_adj_5355));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3835_9.INIT0 = 16'h6969;
    defparam add_3835_9.INIT1 = 16'h9995;
    defparam add_3835_9.INJECT1_0 = "NO";
    defparam add_3835_9.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_30 (.A0(d5[28]), .B0(d4[28]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[29]), .B1(d4[29]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16373), .COUT(n16374), .S0(d5_71__N_706[28]), .S1(d5_71__N_706[29]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_28 (.A0(d5[26]), .B0(d4[26]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[27]), .B1(d4[27]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16372), .COUT(n16373), .S0(d5_71__N_706[26]), .S1(d5_71__N_706[27]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_28.INJECT1_1 = "NO";
    AMDemodulator AMDemodulator_inst (.\DataInReg_11__N_1856[0] (DataInReg_11__N_1856[0]), 
            .CIC1_out_clkSin(CIC1_out_clkSin), .CIC1_outCos({CIC1_outCos}), 
            .MultResult2({MultResult2}), .\d_out_d_11__N_1880[17] (d_out_d_11__N_1880[17]), 
            .d_out_d_11__N_1879(d_out_d_11__N_1879), .\d_out_d_11__N_1878[17] (d_out_d_11__N_1878[17]), 
            .d_out_d_11__N_1877(d_out_d_11__N_1877), .\d_out_d_11__N_1876[17] (d_out_d_11__N_1876[17]), 
            .d_out_d_11__N_1875(d_out_d_11__N_1875), .MultDataB({MultDataB}), 
            .MultResult1({MultResult1}), .VCC_net(VCC_net), .GND_net(GND_net), 
            .\DataInReg_11__N_1856[1] (DataInReg_11__N_1856[1]), .\DataInReg_11__N_1856[2] (DataInReg_11__N_1856[2]), 
            .\DataInReg_11__N_1856[3] (DataInReg_11__N_1856[3]), .\DataInReg_11__N_1856[4] (DataInReg_11__N_1856[4]), 
            .\DataInReg_11__N_1856[5] (DataInReg_11__N_1856[5]), .\DataInReg_11__N_1856[6] (DataInReg_11__N_1856[6]), 
            .\DataInReg_11__N_1856[7] (DataInReg_11__N_1856[7]), .\DataInReg_11__N_1856[8] (DataInReg_11__N_1856[8]), 
            .\DemodOut[9] (DemodOut[9]), .\d_out_d_11__N_2383[17] (d_out_d_11__N_2383[17]), 
            .\d_out_d_11__N_2401[17] (d_out_d_11__N_2401[17]), .\d_out_d_11__N_1892[17] (d_out_d_11__N_1892[17]), 
            .\ISquare[31] (ISquare[31]), .n213(n213_adj_4637), .\d_out_d_11__N_1874[17] (d_out_d_11__N_1874[17]), 
            .d_out_d_11__N_1873(d_out_d_11__N_1873), .\d_out_d_11__N_1888[17] (d_out_d_11__N_1888[17]), 
            .\d_out_d_11__N_1890[17] (d_out_d_11__N_1890[17]), .\d_out_d_11__N_1886[17] (d_out_d_11__N_1886[17]), 
            .\d_out_d_11__N_1884[17] (d_out_d_11__N_1884[17]), .\d_out_d_11__N_1882[17] (d_out_d_11__N_1882[17])) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(171[18] 176[5])
    CCU2C _add_1_1421_add_4_26 (.A0(d5[24]), .B0(d4[24]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[25]), .B1(d4[25]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16371), .COUT(n16372), .S0(d5_71__N_706[24]), .S1(d5_71__N_706[25]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_26.INJECT1_1 = "NO";
    CCU2C add_3835_7 (.A0(d_out_d_11__N_1876[17]), .B0(d_out_d_11__N_1880[17]), 
          .C0(n74), .D0(VCC_net), .A1(d_out_d_11__N_1874[17]), .B1(d_out_d_11__N_1880[17]), 
          .C1(n71), .D1(VCC_net), .CIN(n16559), .COUT(n16560), .S0(n81_adj_5358), 
          .S1(n78_adj_5357));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3835_7.INIT0 = 16'h9696;
    defparam add_3835_7.INIT1 = 16'h9696;
    defparam add_3835_7.INJECT1_0 = "NO";
    defparam add_3835_7.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16340), .S0(cout_adj_5534));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1406_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1406_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_24 (.A0(d5[22]), .B0(d4[22]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[23]), .B1(d4[23]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16370), .COUT(n16371), .S0(d5_71__N_706[22]), .S1(d5_71__N_706[23]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_24.INJECT1_1 = "NO";
    PFUMX i6415 (.BLUT(n17952), .ALUT(n17953), .C0(n316), .Z(n17954));
    CCU2C _add_1_1421_add_4_22 (.A0(d5[20]), .B0(d4[20]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[21]), .B1(d4[21]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16369), .COUT(n16370), .S0(d5_71__N_706[20]), .S1(d5_71__N_706[21]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_22.INJECT1_1 = "NO";
    CCU2C add_3835_5 (.A0(n80), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1878[17]), .B1(d_out_d_11__N_1880[17]), .C1(n77), 
          .D1(VCC_net), .CIN(n16558), .COUT(n16559), .S0(n87_adj_5360), 
          .S1(n84_adj_5359));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3835_5.INIT0 = 16'haaa0;
    defparam add_3835_5.INIT1 = 16'h9696;
    defparam add_3835_5.INJECT1_0 = "NO";
    defparam add_3835_5.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_20 (.A0(d5[18]), .B0(d4[18]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[19]), .B1(d4[19]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16368), .COUT(n16369), .S0(d5_71__N_706[18]), .S1(d5_71__N_706[19]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_18 (.A0(d5[16]), .B0(d4[16]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[17]), .B1(d4[17]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16367), .COUT(n16368), .S0(d5_71__N_706[16]), .S1(d5_71__N_706[17]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_16 (.A0(d5[14]), .B0(d4[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[15]), .B1(d4[15]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16366), .COUT(n16367), .S0(d5_71__N_706[14]), .S1(d5_71__N_706[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_16.INJECT1_1 = "NO";
    CCU2C add_3835_3 (.A0(d_out_d_11__N_1880[17]), .B0(ISquare[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(ISquare[13]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16557), .COUT(n16558), .S1(n90_adj_5361));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3835_3.INIT0 = 16'h666a;
    defparam add_3835_3.INIT1 = 16'h555f;
    defparam add_3835_3.INJECT1_0 = "NO";
    defparam add_3835_3.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_14 (.A0(d5[12]), .B0(d4[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[13]), .B1(d4[13]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16365), .COUT(n16366), .S0(d5_71__N_706[12]), .S1(d5_71__N_706[13]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_12 (.A0(d5[10]), .B0(d4[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[11]), .B1(d4[11]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16364), .COUT(n16365), .S0(d5_71__N_706[10]), .S1(d5_71__N_706[11]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_12.INJECT1_1 = "NO";
    CCU2C add_3835_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(d_out_d_11__N_1880[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16557));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam add_3835_1.INIT0 = 16'h0000;
    defparam add_3835_1.INIT1 = 16'haaaf;
    defparam add_3835_1.INJECT1_0 = "NO";
    defparam add_3835_1.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_10 (.A0(d5[8]), .B0(d4[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(d5[9]), .B1(d4[9]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n16363), .COUT(n16364), .S0(d5_71__N_706[8]), .S1(d5_71__N_706[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_8 (.A0(d5[6]), .B0(d4[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[7]), .B1(d4[7]), .C1(GND_net), .D1(VCC_net), .CIN(n16362), 
          .COUT(n16363), .S0(d5_71__N_706[6]), .S1(d5_71__N_706[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_6 (.A0(d5[4]), .B0(d4[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[5]), .B1(d4[5]), .C1(GND_net), .D1(VCC_net), .CIN(n16361), 
          .COUT(n16362), .S0(d5_71__N_706[4]), .S1(d5_71__N_706[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1406_add_4_36 (.A0(d1[34]), .B0(MixerOutSin[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(d1[35]), .B1(MixerOutSin[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16339), .COUT(n16340), .S0(d1_71__N_418[34]), 
          .S1(d1_71__N_418[35]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(62[15:24])
    defparam _add_1_1406_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1406_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1406_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1406_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1421_add_4_4 (.A0(d5[2]), .B0(d4[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(d5[3]), .B1(d4[3]), .C1(GND_net), .D1(VCC_net), .CIN(n16360), 
          .COUT(n16361), .S0(d5_71__N_706[2]), .S1(d5_71__N_706[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(66[15:24])
    defparam _add_1_1421_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1421_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1421_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1421_add_4_4.INJECT1_1 = "NO";
    \CIC(WIDTH=72,DECIMATION_RATIO=4096)_U0  CIC_Sin_inst (.d_tmp({d_tmp}), 
            .clk_80mhz(clk_80mhz), .d5({d5}), .d_d_tmp({d_d_tmp}), .d2({d2}), 
            .d2_71__N_490({d2_71__N_490}), .d_d8({d_d8}), .n11(n11_adj_4869), 
            .d3({d3}), .d3_71__N_562({d3_71__N_562}), .d4({d4}), .d4_71__N_634({d4_71__N_634}), 
            .d5_71__N_706({d5_71__N_706}), .d6({d6}), .d6_71__N_1459({d6_71__N_1459}), 
            .d_d6({d_d6}), .CIC1_out_clkSin(CIC1_out_clkSin), .d7({d7}), 
            .d7_71__N_1531({d7_71__N_1531}), .d_d7({d_d7}), .d8({d8}), 
            .d8_71__N_1603({d8_71__N_1603}), .d9({d9}), .d9_71__N_1675({d9_71__N_1675}), 
            .d_d9({d_d9}), .n26(n26_adj_4830), .MultDataB({MultDataB}), 
            .d1({d1}), .d1_71__N_418({d1_71__N_418}), .count({count}), 
            .n29(n29_adj_4827), .n10(n10_adj_4870), .n13(n13_adj_4867), 
            .n12(n12_adj_4868), .n15(n15_adj_4865), .\CICGain[1] (CICGain[1]), 
            .n18(n18_adj_4776), .n21(n21_adj_4773), .n20(n20_adj_4774), 
            .n23(n23_adj_4771), .n22(n22_adj_4772), .n25(n25_adj_4769), 
            .n24(n24_adj_4770), .n27(n27_adj_4767), .n26_adj_1(n26_adj_4768), 
            .n29_adj_2(n29_adj_4765), .n28(n28_adj_4766), .n31(n31_adj_4763), 
            .n30(n30_adj_4764), .n33(n33_adj_4761), .n118(n118), .n120(n120_adj_5274), 
            .cout(cout_adj_4756), .n115(n115), .n117(n117_adj_5273), .n112(n112), 
            .n114(n114_adj_5272), .n32(n32_adj_4762), .n35(n35_adj_4759), 
            .n109(n109), .n111(n111_adj_5271), .n34(n34_adj_4760), .n106(n106), 
            .n108(n108_adj_5270), .n37(n37_adj_4757), .n103(n103), .n105(n105_adj_5269), 
            .n36(n36_adj_4758), .n3(n3_adj_4817), .n2(n2_adj_4818), .n100(n100), 
            .n102(n102_adj_5268), .n97(n97), .n99(n99_adj_5267), .n5(n5_adj_4815), 
            .n4(n4_adj_4816), .n94(n94), .n96(n96_adj_5266), .n91(n91), 
            .n93(n93_adj_5265), .n88(n88), .n90(n90_adj_5264), .n7(n7_adj_4813), 
            .n85(n85), .n87(n87_adj_5263), .n82(n82), .n84(n84_adj_5262), 
            .n79(n79), .n81(n81_adj_5261), .n76(n76), .n78(n78_adj_5260), 
            .n14(n14_adj_4866), .n6(n6_adj_4814), .n8(n8_adj_4714), .\d10[68] (d10[68]), 
            .\d10[66] (d10[66]), .\d10[67] (d10[67]), .n28_adj_3(n28_adj_4828), 
            .n31_adj_4(n31_adj_4825), .n11_adj_5(n11_adj_4651), .n9(n9_adj_4811), 
            .\d10[65] (d10[65]), .\d_out_11__N_1819[2] (d_out_11__N_1819[2]), 
            .\d_out_11__N_1819[3] (d_out_11__N_1819[3]), .\d_out_11__N_1819[4] (d_out_11__N_1819[4]), 
            .\d_out_11__N_1819[5] (d_out_11__N_1819[5]), .\d_out_11__N_1819[6] (d_out_11__N_1819[6]), 
            .\d_out_11__N_1819[7] (d_out_11__N_1819[7]), .\d_out_11__N_1819[8] (d_out_11__N_1819[8]), 
            .n87_adj_126({n36_adj_5328, n39_adj_5329, n42_adj_5330, n45_adj_5331, 
            n48_adj_5332, n51_adj_5333, n54_adj_5334, n57_adj_5335, 
            n60_adj_5336, n63_adj_5337, n66_adj_5338, n69_adj_5339, 
            n72_adj_5340, n75_adj_5341, n78_adj_5342, n81_adj_5343}), 
            .\CICGain[0] (CICGain[0]), .n30_adj_9(n30_adj_4826), .n63_adj_10(n63), 
            .n65(n65), .n135(n135_adj_4793), .n64(n64), .n134(n134), 
            .n133(n133), .n8_adj_11(n8_adj_4812), .n132(n132_adj_4792), 
            .n66_adj_12(n66), .n136(n136), .n11_adj_13(n11_adj_4809), 
            .n10_adj_14(n10_adj_4810), .n66_adj_15(n66_adj_4798), .\d10[64] (d10_adj_5753[64]), 
            .n136_adj_16(n136_adj_4804), .n65_adj_17(n65_adj_4797), .\d10[63] (d10_adj_5753[63]), 
            .n135_adj_18(n135_adj_4803), .n63_adj_19(n63_adj_4795), .\d10[61] (d10_adj_5753[61]), 
            .n133_adj_20(n133_adj_4801), .n13_adj_21(n13_adj_4807), .\d10[68]_adj_22 (d10_adj_5753[68]), 
            .\d10[69] (d10_adj_5753[69]), .\d10[71] (d10_adj_5753[71]), 
            .\d10[70] (d10_adj_5753[70]), .n64_adj_23(n64_adj_4796), .\d10[62] (d10_adj_5753[62]), 
            .n134_adj_24(n134_adj_4802), .n17(n17_adj_4863), .n16(n16_adj_4864), 
            .n19(n19_adj_4861), .n18_adj_25(n18_adj_4862), .n21_adj_26(n21_adj_4859), 
            .n20_adj_27(n20_adj_4860), .n23_adj_28(n23_adj_4857), .n22_adj_29(n22_adj_4858), 
            .n17610(n17610), .\d10[60] (d10_adj_5753[60]), .n132_adj_30(n132_adj_4800), 
            .n17630(n17630), .\d10[59] (d10_adj_5753[59]), .n131(n131_adj_4799), 
            .n12_adj_31(n12_adj_4808), .n3_adj_32(n3_adj_4626), .n2_adj_33(n2_adj_4627), 
            .n10_adj_34(n10_adj_4676), .n13_adj_35(n13_adj_4636), .n12_adj_36(n12_adj_4638), 
            .n15_adj_37(n15_adj_4634), .n14_adj_38(n14_adj_4635), .n17_adj_39(n17_adj_4632), 
            .n16_adj_40(n16_adj_4633), .n19_adj_41(n19_adj_4630), .n131_adj_42(n131), 
            .\d10[67]_adj_43 (d10_adj_5753[67]), .n18_adj_44(n18_adj_4631), 
            .n21_adj_45(n21_adj_4628), .n20_adj_46(n20_adj_4629), .n23_adj_47(n23_adj_4856), 
            .n22_adj_48(n22_adj_4879), .n25_adj_49(n25_adj_4831), .n24_adj_50(n24_adj_4832), 
            .n25_adj_51(n25), .n24_adj_52(n24), .n27_adj_53(n27), .n26_adj_54(n26), 
            .n29_adj_55(n29), .n28_adj_56(n28), .n31_adj_57(n31), .n30_adj_58(n30), 
            .n33_adj_59(n33_adj_4755), .n32_adj_60(n32_adj_4855), .n27_adj_61(n27_adj_4829), 
            .n35_adj_62(n35_adj_4753), .n34_adj_63(n34_adj_4754), .n37_adj_64(n37_adj_4747), 
            .n36_adj_65(n36_adj_4752), .n15_adj_66(n15_adj_4805), .n14_adj_67(n14_adj_4806), 
            .n17_adj_68(n17_adj_4833), .n16_adj_69(n16_adj_4834), .n5_adj_70(n5_adj_4789), 
            .n4_adj_71(n4_adj_4790), .n33_adj_72(n33_adj_4823), .n7_adj_73(n7_adj_4787), 
            .n32_adj_74(n32_adj_4824), .n35_adj_75(n35_adj_4821), .n34_adj_76(n34_adj_4822), 
            .n6_adj_77(n6_adj_4788), .n9_adj_78(n9_adj_4785), .n8_adj_79(n8_adj_4786), 
            .n11_adj_80(n11_adj_4783), .n37_adj_81(n37_adj_4819), .n10_adj_82(n10_adj_4784), 
            .n36_adj_83(n36_adj_4820), .n13_adj_84(n13_adj_4781), .n3_adj_85(n3_adj_4750), 
            .n2_adj_86(n2_adj_4751), .n5_adj_87(n5_adj_4748), .n12_adj_88(n12_adj_4782), 
            .n4_adj_89(n4_adj_4749), .n7_adj_90(n7_adj_4717), .n15_adj_91(n15_adj_4779), 
            .n14_adj_92(n14_adj_4780), .n6_adj_93(n6_adj_4746), .n17_adj_94(n17_adj_4777), 
            .n19_adj_95(n19_adj_4852), .n18_adj_96(n18_adj_4835), .n9_adj_97(n9_adj_4684), 
            .n16_adj_98(n16_adj_4778), .\d_out_11__N_1819[10] (d_out_11__N_1819_adj_5778[10]), 
            .n19_adj_99(n19_adj_4775), .n21_adj_100(n21_adj_4850), .n20_adj_101(n20_adj_4851), 
            .\d_out_11__N_1819[11] (d_out_11__N_1819_adj_5778[11]), .n23_adj_102(n23_adj_4848), 
            .n22_adj_103(n22_adj_4849), .n25_adj_104(n25_adj_4846), .n24_adj_105(n24_adj_4847), 
            .n27_adj_106(n27_adj_4844), .n26_adj_107(n26_adj_4845), .n29_adj_108(n29_adj_4842), 
            .n28_adj_109(n28_adj_4843), .n31_adj_110(n31_adj_4840), .n30_adj_111(n30_adj_4841), 
            .n33_adj_112(n33_adj_4838), .n32_adj_113(n32_adj_4839), .n35_adj_114(n35_adj_4836), 
            .n34_adj_115(n34_adj_4837), .n37_adj_116(n37_adj_4854), .n36_adj_117(n36_adj_4853), 
            .n3_adj_118(n3_adj_4877), .n2_adj_119(n2_adj_4878), .n5_adj_120(n5_adj_4875), 
            .n4_adj_121(n4_adj_4876), .n7_adj_122(n7_adj_4873), .n6_adj_123(n6_adj_4874), 
            .n9_adj_124(n9_adj_4871), .n8_adj_125(n8_adj_4872)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(136[4] 142[5])
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=87) 
//

module \uart_rx(CLKS_PER_BIT=87)  (clk_80mhz, i_Rx_Serial_c, r_Rx_Data, 
            o_Rx_Byte1, \r_Rx_Byte[4] , n17663, GND_net, VCC_net, 
            o_Rx_DV1, n17943, \r_Rx_Byte[6] , n17945, n17397, n17946, 
            n17664) /* synthesis syn_module_defined=1 */ ;
    input clk_80mhz;
    input i_Rx_Serial_c;
    output r_Rx_Data;
    output [7:0]o_Rx_Byte1;
    output \r_Rx_Byte[4] ;
    input n17663;
    input GND_net;
    input VCC_net;
    output o_Rx_DV1;
    output n17943;
    output \r_Rx_Byte[6] ;
    output n17945;
    output n17397;
    output n17946;
    input n17664;
    
    wire [7:0]UartClk /* synthesis SET_AS_NETWORK=\uart_rx_inst/UartClk[2], is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(37[14:21])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(61[23:32])
    wire [2:0]r_SM_Main;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(43[17:26])
    
    wire n17826, r_Rx_DV_last, r_Rx_DV, r_Rx_Data_R, UartClk_2_enable_15;
    wire [7:0]r_Rx_Byte;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(41[17:26])
    
    wire UartClk_2_enable_2, n17091, UartClk_2_enable_30;
    wire [2:0]r_Bit_Index;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(40[17:28])
    
    wire UartClk_2_enable_32, n17086, n18, n17935, n12696, UartClk_2_enable_4, 
        n17936, n17828, n16532;
    wire [2:0]n30;
    wire [2:0]n17;
    
    wire n17827, UartClk_2_enable_5, n12693, r_Rx_DV_last_N_2531, UartClk_2_enable_6, 
        n16531;
    wire [15:0]r_Clock_Count;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(39[18:31])
    wire [15:0]n69;
    
    wire n17107, UartClk_2_enable_7, n16530, n16529, n16528, n16527, 
        n16526, n16525, n16524, n17829, n17825, n193, n17085, 
        n17421, n17423, n17425, n17411, n16773, UartClk_2_enable_35, 
        n17060, UartClk_2_enable_36, n208, n17300, UartClk_2_enable_33, 
        n17928, n17824, n17373, n17365, n17183, n17361, n17135, 
        n17950, n17949, UartClk_2_enable_34, n17947, n17441;
    
    FD1S3IX r_SM_Main_i0 (.D(n17826), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i0.GSR = "ENABLED";
    FD1S3AX r_Rx_DV_last_60 (.D(r_Rx_DV), .CK(clk_80mhz), .Q(r_Rx_DV_last)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(47[11] 52[8])
    defparam r_Rx_DV_last_60.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_R_61 (.D(i_Rx_Serial_c), .CK(UartClk[2]), .Q(r_Rx_Data_R)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(57[11] 62[8])
    defparam r_Rx_Data_R_61.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_62 (.D(r_Rx_Data_R), .CK(UartClk[2]), .Q(r_Rx_Data)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(57[11] 62[8])
    defparam r_Rx_Data_62.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i0 (.D(r_Rx_Byte[0]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i0.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i4 (.D(n17663), .SP(UartClk_2_enable_2), .CK(UartClk[2]), 
            .Q(\r_Rx_Byte[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i4.GSR = "ENABLED";
    LUT4 i6360_4_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(n17091), 
         .D(r_Rx_Data), .Z(UartClk_2_enable_30)) /* synthesis lut_function=(!(A (B)+!A (B+(C (D))))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(69[7] 161[14])
    defparam i6360_4_lut.init = 16'h2333;
    FD1P3AX r_Bit_Index_i0 (.D(n17086), .SP(UartClk_2_enable_32), .CK(UartClk[2]), 
            .Q(r_Bit_Index[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i0.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(r_SM_Main[2]), .B(n18), .C(n17935), .D(r_SM_Main[1]), 
         .Z(n12696)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i1_4_lut.init = 16'h5044;
    FD1P3AX r_Rx_Byte_i3 (.D(r_Rx_Data), .SP(UartClk_2_enable_4), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i3.GSR = "ENABLED";
    LUT4 r_SM_Main_2__N_2466_2__bdd_3_lut (.A(r_Rx_Data), .B(r_SM_Main[0]), 
         .C(n17936), .Z(n17828)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam r_SM_Main_2__N_2466_2__bdd_3_lut.init = 16'h0404;
    CCU2C UartClk_1006_1032_add_4_3 (.A0(n30[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(UartClk[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16532), .S0(n17[1]), .S1(n17[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_1006_1032_add_4_3.INIT0 = 16'haaa0;
    defparam UartClk_1006_1032_add_4_3.INIT1 = 16'haaa0;
    defparam UartClk_1006_1032_add_4_3.INJECT1_0 = "NO";
    defparam UartClk_1006_1032_add_4_3.INJECT1_1 = "NO";
    LUT4 r_SM_Main_2__N_2466_2__bdd_2_lut (.A(n17935), .B(r_SM_Main[0]), 
         .Z(n17827)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam r_SM_Main_2__N_2466_2__bdd_2_lut.init = 16'h7777;
    LUT4 i6349_4_lut (.A(r_SM_Main[0]), .B(r_SM_Main[1]), .C(r_SM_Main[2]), 
         .D(n17935), .Z(UartClk_2_enable_32)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B (C)))) */ ;
    defparam i6349_4_lut.init = 16'h0501;
    FD1P3AX r_Rx_Byte_i2 (.D(r_Rx_Data), .SP(UartClk_2_enable_5), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i2.GSR = "ENABLED";
    FD1S3IX o_Rx_DV_59 (.D(r_Rx_DV_last_N_2531), .CK(clk_80mhz), .CD(n12693), 
            .Q(o_Rx_DV1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(47[11] 52[8])
    defparam o_Rx_DV_59.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i1 (.D(r_Rx_Data), .SP(UartClk_2_enable_6), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i1.GSR = "ENABLED";
    FD1S3AX UartClk_1006_1032__i0 (.D(n17[0]), .CK(clk_80mhz), .Q(n30[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_1006_1032__i0.GSR = "ENABLED";
    CCU2C UartClk_1006_1032_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n16532), .S1(n17[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_1006_1032_add_4_1.INIT0 = 16'h0000;
    defparam UartClk_1006_1032_add_4_1.INIT1 = 16'h555f;
    defparam UartClk_1006_1032_add_4_1.INJECT1_0 = "NO";
    defparam UartClk_1006_1032_add_4_1.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1008_add_4_17 (.A0(r_Clock_Count[15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n16531), .S0(n69[15]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008_add_4_17.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_17.INIT1 = 16'h0000;
    defparam r_Clock_Count_1008_add_4_17.INJECT1_0 = "NO";
    defparam r_Clock_Count_1008_add_4_17.INJECT1_1 = "NO";
    FD1S3IX r_SM_Main_i2 (.D(n17935), .CK(UartClk[2]), .CD(n17107), .Q(r_SM_Main[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i2.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i0 (.D(r_Rx_Data), .SP(UartClk_2_enable_7), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_171 (.A(r_SM_Main[1]), .B(r_SM_Main[0]), .Z(n17943)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i1_2_lut_rep_171.init = 16'h2222;
    LUT4 i1_2_lut_rep_155_3_lut (.A(r_SM_Main[1]), .B(r_SM_Main[0]), .C(n17935), 
         .Z(UartClk_2_enable_2)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i1_2_lut_rep_155_3_lut.init = 16'h2020;
    CCU2C r_Clock_Count_1008_add_4_15 (.A0(r_Clock_Count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16530), .COUT(n16531), .S0(n69[13]), 
          .S1(n69[14]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008_add_4_15.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_15.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_15.INJECT1_0 = "NO";
    defparam r_Clock_Count_1008_add_4_15.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1008_add_4_13 (.A0(r_Clock_Count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16529), .COUT(n16530), .S0(n69[11]), 
          .S1(n69[12]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008_add_4_13.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_13.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_13.INJECT1_0 = "NO";
    defparam r_Clock_Count_1008_add_4_13.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1008_add_4_11 (.A0(r_Clock_Count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16528), .COUT(n16529), .S0(n69[9]), 
          .S1(n69[10]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008_add_4_11.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_11.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_11.INJECT1_0 = "NO";
    defparam r_Clock_Count_1008_add_4_11.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1008_add_4_9 (.A0(r_Clock_Count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16527), .COUT(n16528), .S0(n69[7]), 
          .S1(n69[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008_add_4_9.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_9.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_9.INJECT1_0 = "NO";
    defparam r_Clock_Count_1008_add_4_9.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1008_add_4_7 (.A0(r_Clock_Count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16526), .COUT(n16527), .S0(n69[5]), 
          .S1(n69[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008_add_4_7.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_7.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_7.INJECT1_0 = "NO";
    defparam r_Clock_Count_1008_add_4_7.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1008_add_4_5 (.A0(r_Clock_Count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16525), .COUT(n16526), .S0(n69[3]), 
          .S1(n69[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008_add_4_5.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_5.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_5.INJECT1_0 = "NO";
    defparam r_Clock_Count_1008_add_4_5.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1008_add_4_3 (.A0(r_Clock_Count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n16524), .COUT(n16525), .S0(n69[1]), 
          .S1(n69[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008_add_4_3.INIT0 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_3.INIT1 = 16'haaa0;
    defparam r_Clock_Count_1008_add_4_3.INJECT1_0 = "NO";
    defparam r_Clock_Count_1008_add_4_3.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_1008_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(r_Clock_Count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16524), .S1(n69[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008_add_4_1.INIT0 = 16'h0000;
    defparam r_Clock_Count_1008_add_4_1.INIT1 = 16'h555f;
    defparam r_Clock_Count_1008_add_4_1.INJECT1_0 = "NO";
    defparam r_Clock_Count_1008_add_4_1.INJECT1_1 = "NO";
    FD1S3IX r_SM_Main_i1 (.D(n17829), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i1.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i1 (.D(r_Rx_Byte[1]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i0 (.D(n69[0]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i0.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i2 (.D(r_Rx_Byte[2]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i3 (.D(r_Rx_Byte[3]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i4 (.D(\r_Rx_Byte[4] ), .SP(UartClk_2_enable_15), 
            .CK(UartClk[2]), .Q(o_Rx_Byte1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i5 (.D(r_Rx_Byte[5]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i6 (.D(\r_Rx_Byte[6] ), .SP(UartClk_2_enable_15), 
            .CK(UartClk[2]), .Q(o_Rx_Byte1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i7 (.D(r_Rx_Byte[7]), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(o_Rx_Byte1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(r_SM_Main[1]), .B(r_SM_Main[0]), .C(r_Bit_Index[0]), 
         .D(n17935), .Z(n17086)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 r_SM_Main_2__N_2466_2__bdd_3_lut_6377 (.A(n17936), .B(r_Rx_Data), 
         .C(r_SM_Main[0]), .Z(n17825)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+(C))) */ ;
    defparam r_SM_Main_2__N_2466_2__bdd_3_lut_6377.init = 16'ha3a3;
    LUT4 i6339_2_lut_3_lut (.A(n193), .B(r_Bit_Index[1]), .C(r_Bit_Index[0]), 
         .Z(UartClk_2_enable_4)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i6339_2_lut_3_lut.init = 16'h4040;
    LUT4 i6337_2_lut_3_lut (.A(n193), .B(r_Bit_Index[1]), .C(r_Bit_Index[0]), 
         .Z(UartClk_2_enable_5)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i6337_2_lut_3_lut.init = 16'h0404;
    LUT4 i1_3_lut_4_lut (.A(n17935), .B(n17943), .C(r_Bit_Index[1]), .D(r_Bit_Index[0]), 
         .Z(n17085)) /* synthesis lut_function=(!(((C (D)+!C !(D))+!B)+!A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i1_3_lut_4_lut.init = 16'h0880;
    LUT4 i1_4_lut_adj_47 (.A(n17421), .B(n17423), .C(n17425), .D(n17411), 
         .Z(n16773)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_47.init = 16'hfffe;
    LUT4 i1_2_lut (.A(r_Clock_Count[15]), .B(r_Clock_Count[2]), .Z(n17421)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_48 (.A(r_Clock_Count[12]), .B(r_Clock_Count[11]), 
         .C(r_Clock_Count[7]), .D(r_Clock_Count[14]), .Z(n17423)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_48.init = 16'hfffe;
    LUT4 i1_4_lut_adj_49 (.A(r_Clock_Count[9]), .B(r_Clock_Count[10]), .C(r_Clock_Count[8]), 
         .D(r_Clock_Count[4]), .Z(n17425)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_49.init = 16'hfffe;
    LUT4 i208_2_lut_rep_173 (.A(r_Bit_Index[0]), .B(r_SM_Main[2]), .Z(n17945)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i208_2_lut_rep_173.init = 16'heeee;
    LUT4 i1_2_lut_adj_50 (.A(r_Clock_Count[13]), .B(r_Clock_Count[6]), .Z(n17411)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_50.init = 16'heeee;
    LUT4 i1_2_lut_adj_51 (.A(r_Bit_Index[2]), .B(n17935), .Z(UartClk_2_enable_35)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i1_2_lut_adj_51.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(r_Bit_Index[0]), .B(r_SM_Main[2]), .C(r_Bit_Index[1]), 
         .Z(n17397)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_rep_174 (.A(r_Bit_Index[1]), .B(r_Bit_Index[2]), .Z(n17946)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_174.init = 16'hbbbb;
    LUT4 i6342_2_lut_3_lut (.A(r_Bit_Index[1]), .B(r_Bit_Index[2]), .C(n17060), 
         .Z(UartClk_2_enable_36)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i6342_2_lut_3_lut.init = 16'h0404;
    LUT4 i1_4_lut_adj_52 (.A(n208), .B(n17935), .C(n17943), .D(r_Bit_Index[2]), 
         .Z(n17300)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C (D))))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i1_4_lut_adj_52.init = 16'h4080;
    LUT4 i6344_3_lut (.A(r_Bit_Index[1]), .B(n17060), .C(r_Bit_Index[2]), 
         .Z(UartClk_2_enable_33)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(114[17:39])
    defparam i6344_3_lut.init = 16'h2020;
    LUT4 i1_4_lut_adj_53 (.A(r_Bit_Index[0]), .B(n17928), .C(r_SM_Main[1]), 
         .D(r_SM_Main[0]), .Z(n17060)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i1_4_lut_adj_53.init = 16'hffdf;
    LUT4 i1_2_lut_adj_54 (.A(r_Bit_Index[1]), .B(r_Bit_Index[0]), .Z(n208)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(40[17:28])
    defparam i1_2_lut_adj_54.init = 16'h8888;
    LUT4 i6323_2_lut_3_lut (.A(r_Bit_Index[1]), .B(n193), .C(r_Bit_Index[0]), 
         .Z(UartClk_2_enable_7)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i6323_2_lut_3_lut.init = 16'h0101;
    LUT4 r_SM_Main_2__N_2466_2__bdd_4_lut (.A(n17935), .B(n208), .C(r_SM_Main[0]), 
         .D(r_Bit_Index[2]), .Z(n17824)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(C))) */ ;
    defparam r_SM_Main_2__N_2466_2__bdd_4_lut.init = 16'h5850;
    LUT4 i1_4_lut_rep_163 (.A(n17373), .B(n17365), .C(r_Clock_Count[6]), 
         .D(n17183), .Z(n17935)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_rep_163.init = 16'hfeee;
    LUT4 i1_2_lut_rep_156 (.A(r_SM_Main[2]), .B(n17935), .Z(n17928)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i1_2_lut_rep_156.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_55 (.A(r_Clock_Count[12]), .B(r_Clock_Count[7]), .C(r_Clock_Count[14]), 
         .D(r_Clock_Count[9]), .Z(n17373)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_55.init = 16'hfffe;
    LUT4 i1_4_lut_adj_56 (.A(r_Clock_Count[15]), .B(n17361), .C(r_Clock_Count[11]), 
         .D(r_Clock_Count[10]), .Z(n17365)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_56.init = 16'hfffe;
    LUT4 i5891_4_lut (.A(r_Clock_Count[5]), .B(r_Clock_Count[4]), .C(r_Clock_Count[3]), 
         .D(n17135), .Z(n17183)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i5891_4_lut.init = 16'heeea;
    LUT4 i2873_1_lut (.A(r_Rx_DV), .Z(n12693)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i2873_1_lut.init = 16'h5555;
    LUT4 r_Rx_DV_last_I_0_1_lut (.A(r_Rx_DV_last), .Z(r_Rx_DV_last_N_2531)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(50[30:43])
    defparam r_Rx_DV_last_I_0_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_adj_57 (.A(r_Clock_Count[13]), .B(r_Clock_Count[8]), .Z(n17361)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_57.init = 16'heeee;
    LUT4 i5844_2_lut (.A(r_Clock_Count[1]), .B(r_Clock_Count[2]), .Z(n17135)) /* synthesis lut_function=(A (B)) */ ;
    defparam i5844_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_4_lut (.A(n17950), .B(n17949), .C(n16773), .D(r_SM_Main[0]), 
         .Z(n17091)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0800;
    LUT4 i6334_2_lut_3_lut (.A(r_Bit_Index[1]), .B(n193), .C(r_Bit_Index[0]), 
         .Z(UartClk_2_enable_6)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i6334_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_3_lut_rep_151_4_lut (.A(r_SM_Main[2]), .B(n17935), .C(r_SM_Main[1]), 
         .D(r_SM_Main[0]), .Z(UartClk_2_enable_15)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i1_3_lut_rep_151_4_lut.init = 16'h4000;
    LUT4 i1_3_lut_3_lut_4_lut (.A(r_SM_Main[2]), .B(n17935), .C(r_SM_Main[1]), 
         .D(r_SM_Main[0]), .Z(UartClk_2_enable_34)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam i1_3_lut_3_lut_4_lut.init = 16'h400f;
    LUT4 i1_4_lut_4_lut (.A(n17935), .B(r_Bit_Index[2]), .C(r_SM_Main[0]), 
         .D(n17947), .Z(n193)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_4_lut.init = 16'hfffd;
    FD1P3IX r_Clock_Count_1008__i15 (.D(n69[15]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[15])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i15.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i14 (.D(n69[14]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[14])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i14.GSR = "ENABLED";
    PFUMX i6378 (.BLUT(n17828), .ALUT(n17827), .C0(r_SM_Main[1]), .Z(n17829));
    LUT4 i1_2_lut_rep_175 (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .Z(n17947)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_175.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_adj_58 (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(r_SM_Main[0]), 
         .Z(n17107)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_58.init = 16'hbfbf;
    PFUMX i6375 (.BLUT(n17825), .ALUT(n17824), .C0(r_SM_Main[1]), .Z(n17826));
    FD1S3AX UartClk_1006_1032__i1 (.D(n17[1]), .CK(clk_80mhz), .Q(n30[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_1006_1032__i1.GSR = "ENABLED";
    FD1S3AX UartClk_1006_1032__i2 (.D(n17[2]), .CK(clk_80mhz), .Q(UartClk[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(49[15:29])
    defparam UartClk_1006_1032__i2.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i13 (.D(n69[13]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[13])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i13.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_177 (.A(r_Clock_Count[1]), .B(r_Clock_Count[0]), .Z(n17949)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_177.init = 16'h8888;
    LUT4 i1_3_lut_rep_164_4_lut (.A(r_Clock_Count[1]), .B(r_Clock_Count[0]), 
         .C(n16773), .D(n17950), .Z(n17936)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i1_3_lut_rep_164_4_lut.init = 16'hf7ff;
    FD1P3IX r_Clock_Count_1008__i12 (.D(n69[12]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[12])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i12.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i11 (.D(n69[11]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[11])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i11.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i10 (.D(n69[10]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[10])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i10.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i9 (.D(n69[9]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i9.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i8 (.D(n69[8]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i8.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i7 (.D(n69[7]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i7.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i6 (.D(n69[6]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i6.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i5 (.D(n69[5]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i5.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i4 (.D(n69[4]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i4.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i3 (.D(n69[3]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i3.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i2 (.D(n69[2]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i2.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_1008__i1 (.D(n69[1]), .SP(UartClk_2_enable_30), 
            .CD(n12696), .CK(UartClk[2]), .Q(r_Clock_Count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_1008__i1.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i2 (.D(n17300), .SP(UartClk_2_enable_32), .CK(UartClk[2]), 
            .Q(r_Bit_Index[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i2.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i1 (.D(n17085), .SP(UartClk_2_enable_32), .CK(UartClk[2]), 
            .Q(r_Bit_Index[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i1.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i7 (.D(r_Rx_Data), .SP(UartClk_2_enable_33), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i7.GSR = "ENABLED";
    FD1P3AX r_Rx_DV_64 (.D(UartClk_2_enable_15), .SP(UartClk_2_enable_34), 
            .CK(UartClk[2]), .Q(r_Rx_DV)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_DV_64.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_178 (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), .Z(n17950)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_178.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_59 (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), 
         .C(r_Clock_Count[0]), .D(r_Clock_Count[1]), .Z(n17441)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_59.init = 16'h8000;
    LUT4 i1_4_lut_4_lut_adj_60 (.A(r_Rx_Data), .B(n17441), .C(n16773), 
         .D(r_SM_Main[0]), .Z(n18)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B (D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(87[21:38])
    defparam i1_4_lut_4_lut_adj_60.init = 16'h04ff;
    FD1P3AX r_Rx_Byte_i6 (.D(n17664), .SP(UartClk_2_enable_35), .CK(UartClk[2]), 
            .Q(\r_Rx_Byte[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i5 (.D(r_Rx_Data), .SP(UartClk_2_enable_36), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=33, LSE_RCOL=5, LSE_LLINE=179, LSE_RLINE=184 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i5.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module Mixer
//

module Mixer (MixerOutCos, clk_80mhz, MixerOutSin, DiffOut_c, RFIn_c, 
            \LOCosine[10] , MixerOutCos_11__N_250, \LOCosine[7] , \LOCosine[6] , 
            \LOCosine[11] , \LOCosine[5] , \LOCosine[4] , \LOCosine[3] , 
            \LOSine[1] , MixerOutSin_11__N_236, \LOCosine[2] , \LOCosine[12] , 
            \LOCosine[1] , \LOSine[12] , \LOCosine[9] , \LOCosine[8] , 
            \LOSine[11] , \LOSine[10] , \LOSine[9] , \LOSine[8] , \LOSine[7] , 
            \LOSine[6] , \LOSine[5] , \LOSine[4] , \LOSine[3] , \LOSine[2] ) /* synthesis syn_module_defined=1 */ ;
    output [11:0]MixerOutCos;
    input clk_80mhz;
    output [11:0]MixerOutSin;
    output DiffOut_c;
    input RFIn_c;
    input \LOCosine[10] ;
    input [11:0]MixerOutCos_11__N_250;
    input \LOCosine[7] ;
    input \LOCosine[6] ;
    input \LOCosine[11] ;
    input \LOCosine[5] ;
    input \LOCosine[4] ;
    input \LOCosine[3] ;
    input \LOSine[1] ;
    input [11:0]MixerOutSin_11__N_236;
    input \LOCosine[2] ;
    input \LOCosine[12] ;
    input \LOCosine[1] ;
    input \LOSine[12] ;
    input \LOCosine[9] ;
    input \LOCosine[8] ;
    input \LOSine[11] ;
    input \LOSine[10] ;
    input \LOSine[9] ;
    input \LOSine[8] ;
    input \LOSine[7] ;
    input \LOSine[6] ;
    input \LOSine[5] ;
    input \LOSine[4] ;
    input \LOSine[3] ;
    input \LOSine[2] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(61[23:32])
    wire [11:0]MixerOutCos_11__N_224;
    wire [11:0]MixerOutSin_11__N_212;
    
    wire RFInR;
    
    FD1S3AX MixerOutCos_i10 (.D(MixerOutCos_11__N_224[10]), .CK(clk_80mhz), 
            .Q(MixerOutCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i10.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i9 (.D(MixerOutCos_11__N_224[9]), .CK(clk_80mhz), 
            .Q(MixerOutCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i9.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i8 (.D(MixerOutCos_11__N_224[8]), .CK(clk_80mhz), 
            .Q(MixerOutCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i8.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i7 (.D(MixerOutCos_11__N_224[7]), .CK(clk_80mhz), 
            .Q(MixerOutCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i7.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i6 (.D(MixerOutCos_11__N_224[6]), .CK(clk_80mhz), 
            .Q(MixerOutCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i6.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i5 (.D(MixerOutCos_11__N_224[5]), .CK(clk_80mhz), 
            .Q(MixerOutCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i5.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i4 (.D(MixerOutCos_11__N_224[4]), .CK(clk_80mhz), 
            .Q(MixerOutCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i4.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i3 (.D(MixerOutCos_11__N_224[3]), .CK(clk_80mhz), 
            .Q(MixerOutCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i3.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i2 (.D(MixerOutCos_11__N_224[2]), .CK(clk_80mhz), 
            .Q(MixerOutCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i2.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i0 (.D(MixerOutSin_11__N_212[0]), .CK(clk_80mhz), 
            .Q(MixerOutSin[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i0.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i1 (.D(MixerOutCos_11__N_224[1]), .CK(clk_80mhz), 
            .Q(MixerOutCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i1.GSR = "ENABLED";
    FD1S3AY RFInR_14 (.D(DiffOut_c), .CK(clk_80mhz), .Q(RFInR)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(34[10] 37[6])
    defparam RFInR_14.GSR = "ENABLED";
    FD1S3AX MixerOutCos_i0 (.D(MixerOutCos_11__N_224[0]), .CK(clk_80mhz), 
            .Q(MixerOutCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i0.GSR = "ENABLED";
    FD1S3AY RFInR1_13 (.D(RFIn_c), .CK(clk_80mhz), .Q(DiffOut_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(34[10] 37[6])
    defparam RFInR1_13.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i11 (.D(MixerOutSin_11__N_212[11]), .CK(clk_80mhz), 
            .Q(MixerOutSin[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i11.GSR = "ENABLED";
    LUT4 MixerOutCos_11__I_0_i10_3_lut (.A(\LOCosine[10] ), .B(MixerOutCos_11__N_250[9]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i10_3_lut.init = 16'hcaca;
    FD1S3AX MixerOutSin_i10 (.D(MixerOutSin_11__N_212[10]), .CK(clk_80mhz), 
            .Q(MixerOutSin[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i10.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i9 (.D(MixerOutSin_11__N_212[9]), .CK(clk_80mhz), 
            .Q(MixerOutSin[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i9.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i8 (.D(MixerOutSin_11__N_212[8]), .CK(clk_80mhz), 
            .Q(MixerOutSin[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i8.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i7 (.D(MixerOutSin_11__N_212[7]), .CK(clk_80mhz), 
            .Q(MixerOutSin[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i7.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i6 (.D(MixerOutSin_11__N_212[6]), .CK(clk_80mhz), 
            .Q(MixerOutSin[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i6.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i5 (.D(MixerOutSin_11__N_212[5]), .CK(clk_80mhz), 
            .Q(MixerOutSin[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i5.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i4 (.D(MixerOutSin_11__N_212[4]), .CK(clk_80mhz), 
            .Q(MixerOutSin[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i4.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i3 (.D(MixerOutSin_11__N_212[3]), .CK(clk_80mhz), 
            .Q(MixerOutSin[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i3.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i2 (.D(MixerOutSin_11__N_212[2]), .CK(clk_80mhz), 
            .Q(MixerOutSin[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i2.GSR = "ENABLED";
    FD1S3AX MixerOutSin_i1 (.D(MixerOutSin_11__N_212[1]), .CK(clk_80mhz), 
            .Q(MixerOutSin[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutSin_i1.GSR = "ENABLED";
    LUT4 MixerOutCos_11__I_0_i7_3_lut (.A(\LOCosine[7] ), .B(MixerOutCos_11__N_250[6]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i6_3_lut (.A(\LOCosine[6] ), .B(MixerOutCos_11__N_250[5]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i11_3_lut (.A(\LOCosine[11] ), .B(MixerOutCos_11__N_250[10]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i5_3_lut (.A(\LOCosine[5] ), .B(MixerOutCos_11__N_250[4]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i4_3_lut (.A(\LOCosine[4] ), .B(MixerOutCos_11__N_250[3]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i3_3_lut (.A(\LOCosine[3] ), .B(MixerOutCos_11__N_250[2]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i1_3_lut (.A(\LOSine[1] ), .B(MixerOutSin_11__N_236[0]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i2_3_lut (.A(\LOCosine[2] ), .B(MixerOutCos_11__N_250[1]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i12_3_lut (.A(\LOCosine[12] ), .B(MixerOutCos_11__N_250[11]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i1_3_lut (.A(\LOCosine[1] ), .B(MixerOutCos_11__N_250[0]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i12_3_lut (.A(\LOSine[12] ), .B(MixerOutSin_11__N_236[11]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i9_3_lut (.A(\LOCosine[9] ), .B(MixerOutCos_11__N_250[8]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutCos_11__I_0_i8_3_lut (.A(\LOCosine[8] ), .B(MixerOutCos_11__N_250[7]), 
         .C(RFInR), .Z(MixerOutCos_11__N_224[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutCos_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i11_3_lut (.A(\LOSine[11] ), .B(MixerOutSin_11__N_236[10]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i10_3_lut (.A(\LOSine[10] ), .B(MixerOutSin_11__N_236[9]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i9_3_lut (.A(\LOSine[9] ), .B(MixerOutSin_11__N_236[8]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i8_3_lut (.A(\LOSine[8] ), .B(MixerOutSin_11__N_236[7]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i7_3_lut (.A(\LOSine[7] ), .B(MixerOutSin_11__N_236[6]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i6_3_lut (.A(\LOSine[6] ), .B(MixerOutSin_11__N_236[5]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i5_3_lut (.A(\LOSine[5] ), .B(MixerOutSin_11__N_236[4]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i5_3_lut.init = 16'hcaca;
    FD1S3AX MixerOutCos_i11 (.D(MixerOutCos_11__N_224[11]), .CK(clk_80mhz), 
            .Q(MixerOutCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=122, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(43[10] 51[6])
    defparam MixerOutCos_i11.GSR = "ENABLED";
    LUT4 MixerOutSin_11__I_0_i4_3_lut (.A(\LOSine[4] ), .B(MixerOutSin_11__N_236[3]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i3_3_lut (.A(\LOSine[3] ), .B(MixerOutSin_11__N_236[2]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 MixerOutSin_11__I_0_i2_3_lut (.A(\LOSine[2] ), .B(MixerOutSin_11__N_236[1]), 
         .C(RFInR), .Z(MixerOutSin_11__N_212[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/Mixer.v(47[14] 50[8])
    defparam MixerOutSin_11__I_0_i2_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module PWM
//

module PWM (\DataInReg[0] , clk_80mhz, \DataInReg_11__N_1856[0] , counter, 
            GND_net, VCC_net, \DataInReg[1] , \DataInReg_11__N_1856[1] , 
            \DataInReg[2] , \DataInReg_11__N_1856[2] , \DataInReg[3] , 
            \DataInReg_11__N_1856[3] , \DataInReg[4] , \DataInReg_11__N_1856[4] , 
            \DataInReg[5] , \DataInReg_11__N_1856[5] , \DataInReg[6] , 
            \DataInReg_11__N_1856[6] , \DataInReg[7] , \DataInReg_11__N_1856[7] , 
            \DataInReg[8] , \DataInReg_11__N_1856[8] , \DataInReg[9] , 
            \DemodOut[9] ) /* synthesis syn_module_defined=1 */ ;
    output \DataInReg[0] ;
    input clk_80mhz;
    input \DataInReg_11__N_1856[0] ;
    output [9:0]counter;
    input GND_net;
    input VCC_net;
    output \DataInReg[1] ;
    input \DataInReg_11__N_1856[1] ;
    output \DataInReg[2] ;
    input \DataInReg_11__N_1856[2] ;
    output \DataInReg[3] ;
    input \DataInReg_11__N_1856[3] ;
    output \DataInReg[4] ;
    input \DataInReg_11__N_1856[4] ;
    output \DataInReg[5] ;
    input \DataInReg_11__N_1856[5] ;
    output \DataInReg[6] ;
    input \DataInReg_11__N_1856[6] ;
    output \DataInReg[7] ;
    input \DataInReg_11__N_1856[7] ;
    output \DataInReg[8] ;
    input \DataInReg_11__N_1856[8] ;
    output \DataInReg[9] ;
    input \DemodOut[9] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(61[23:32])
    
    wire clk_80mhz_enable_1406, n16538;
    wire [9:0]n45;
    
    wire n16537, n16536, n16535, n16534;
    wire [11:0]n3955;
    
    wire n17, n15, n11, n12;
    
    FD1P3AX DataInReg__i1 (.D(\DataInReg_11__N_1856[0] ), .SP(clk_80mhz_enable_1406), 
            .CK(clk_80mhz), .Q(\DataInReg[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(41[8] 53[7])
    defparam DataInReg__i1.GSR = "ENABLED";
    CCU2C counter_1005_add_4_11 (.A0(counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n16538), .S0(n45[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005_add_4_11.INIT0 = 16'haaa0;
    defparam counter_1005_add_4_11.INIT1 = 16'h0000;
    defparam counter_1005_add_4_11.INJECT1_0 = "NO";
    defparam counter_1005_add_4_11.INJECT1_1 = "NO";
    CCU2C counter_1005_add_4_9 (.A0(counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16537), .COUT(n16538), .S0(n45[7]), .S1(n45[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005_add_4_9.INIT0 = 16'haaa0;
    defparam counter_1005_add_4_9.INIT1 = 16'haaa0;
    defparam counter_1005_add_4_9.INJECT1_0 = "NO";
    defparam counter_1005_add_4_9.INJECT1_1 = "NO";
    CCU2C counter_1005_add_4_7 (.A0(counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16536), .COUT(n16537), .S0(n45[5]), .S1(n45[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005_add_4_7.INIT0 = 16'haaa0;
    defparam counter_1005_add_4_7.INIT1 = 16'haaa0;
    defparam counter_1005_add_4_7.INJECT1_0 = "NO";
    defparam counter_1005_add_4_7.INJECT1_1 = "NO";
    CCU2C counter_1005_add_4_5 (.A0(counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16535), .COUT(n16536), .S0(n45[3]), .S1(n45[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005_add_4_5.INIT0 = 16'haaa0;
    defparam counter_1005_add_4_5.INIT1 = 16'haaa0;
    defparam counter_1005_add_4_5.INJECT1_0 = "NO";
    defparam counter_1005_add_4_5.INJECT1_1 = "NO";
    CCU2C counter_1005_add_4_3 (.A0(counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n16534), .COUT(n16535), .S0(n45[1]), .S1(n45[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005_add_4_3.INIT0 = 16'haaa0;
    defparam counter_1005_add_4_3.INIT1 = 16'haaa0;
    defparam counter_1005_add_4_3.INJECT1_0 = "NO";
    defparam counter_1005_add_4_3.INJECT1_1 = "NO";
    CCU2C counter_1005_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n16534), .S1(n45[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005_add_4_1.INIT0 = 16'h0000;
    defparam counter_1005_add_4_1.INIT1 = 16'h555f;
    defparam counter_1005_add_4_1.INJECT1_0 = "NO";
    defparam counter_1005_add_4_1.INJECT1_1 = "NO";
    FD1S3AX counter_1005__i0 (.D(n45[0]), .CK(clk_80mhz), .Q(counter[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005__i0.GSR = "ENABLED";
    FD1P3AX DataInReg__i2 (.D(\DataInReg_11__N_1856[1] ), .SP(clk_80mhz_enable_1406), 
            .CK(clk_80mhz), .Q(\DataInReg[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(41[8] 53[7])
    defparam DataInReg__i2.GSR = "ENABLED";
    FD1P3AX DataInReg__i3 (.D(\DataInReg_11__N_1856[2] ), .SP(clk_80mhz_enable_1406), 
            .CK(clk_80mhz), .Q(\DataInReg[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(41[8] 53[7])
    defparam DataInReg__i3.GSR = "ENABLED";
    FD1P3AX DataInReg__i4 (.D(\DataInReg_11__N_1856[3] ), .SP(clk_80mhz_enable_1406), 
            .CK(clk_80mhz), .Q(\DataInReg[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(41[8] 53[7])
    defparam DataInReg__i4.GSR = "ENABLED";
    FD1P3AX DataInReg__i5 (.D(\DataInReg_11__N_1856[4] ), .SP(clk_80mhz_enable_1406), 
            .CK(clk_80mhz), .Q(\DataInReg[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(41[8] 53[7])
    defparam DataInReg__i5.GSR = "ENABLED";
    FD1P3AX DataInReg__i6 (.D(\DataInReg_11__N_1856[5] ), .SP(clk_80mhz_enable_1406), 
            .CK(clk_80mhz), .Q(\DataInReg[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(41[8] 53[7])
    defparam DataInReg__i6.GSR = "ENABLED";
    FD1P3AX DataInReg__i7 (.D(\DataInReg_11__N_1856[6] ), .SP(clk_80mhz_enable_1406), 
            .CK(clk_80mhz), .Q(\DataInReg[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(41[8] 53[7])
    defparam DataInReg__i7.GSR = "ENABLED";
    FD1P3AX DataInReg__i8 (.D(\DataInReg_11__N_1856[7] ), .SP(clk_80mhz_enable_1406), 
            .CK(clk_80mhz), .Q(\DataInReg[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(41[8] 53[7])
    defparam DataInReg__i8.GSR = "ENABLED";
    FD1P3AX DataInReg__i9 (.D(\DataInReg_11__N_1856[8] ), .SP(clk_80mhz_enable_1406), 
            .CK(clk_80mhz), .Q(\DataInReg[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(41[8] 53[7])
    defparam DataInReg__i9.GSR = "ENABLED";
    FD1P3AX DataInReg__i10 (.D(n3955[9]), .SP(clk_80mhz_enable_1406), .CK(clk_80mhz), 
            .Q(\DataInReg[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=156, LSE_RLINE=160 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(41[8] 53[7])
    defparam DataInReg__i10.GSR = "ENABLED";
    LUT4 i6365_4_lut (.A(n17), .B(n15), .C(n11), .D(n12), .Z(clk_80mhz_enable_1406)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(44[11:23])
    defparam i6365_4_lut.init = 16'h0001;
    LUT4 i7_4_lut (.A(counter[3]), .B(counter[2]), .C(counter[1]), .D(counter[9]), 
         .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(44[11:23])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(counter[6]), .B(counter[4]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(44[11:23])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(counter[0]), .B(counter[5]), .Z(n11)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(44[11:23])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2_2_lut (.A(counter[7]), .B(counter[8]), .Z(n12)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(44[11:23])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1155_1_lut (.A(\DemodOut[9] ), .Z(n3955[9])) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(44[7] 46[10])
    defparam i1155_1_lut.init = 16'h5555;
    FD1S3AX counter_1005__i1 (.D(n45[1]), .CK(clk_80mhz), .Q(counter[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005__i1.GSR = "ENABLED";
    FD1S3AX counter_1005__i2 (.D(n45[2]), .CK(clk_80mhz), .Q(counter[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005__i2.GSR = "ENABLED";
    FD1S3AX counter_1005__i3 (.D(n45[3]), .CK(clk_80mhz), .Q(counter[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005__i3.GSR = "ENABLED";
    FD1S3AX counter_1005__i4 (.D(n45[4]), .CK(clk_80mhz), .Q(counter[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005__i4.GSR = "ENABLED";
    FD1S3AX counter_1005__i5 (.D(n45[5]), .CK(clk_80mhz), .Q(counter[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005__i5.GSR = "ENABLED";
    FD1S3AX counter_1005__i6 (.D(n45[6]), .CK(clk_80mhz), .Q(counter[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005__i6.GSR = "ENABLED";
    FD1S3AX counter_1005__i7 (.D(n45[7]), .CK(clk_80mhz), .Q(counter[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005__i7.GSR = "ENABLED";
    FD1S3AX counter_1005__i8 (.D(n45[8]), .CK(clk_80mhz), .Q(counter[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005__i8.GSR = "ENABLED";
    FD1S3AX counter_1005__i9 (.D(n45[9]), .CK(clk_80mhz), .Q(counter[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/PWM.v(43[18:33])
    defparam counter_1005__i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module SinCos
//

module SinCos (clk_80mhz, VCC_net, GND_net, \phase_accum[57] , \phase_accum[58] , 
            \phase_accum[59] , \phase_accum[60] , \phase_accum[61] , \phase_accum[62] , 
            \phase_accum[63] , \LOSine[1] , \LOSine[2] , \LOSine[3] , 
            \LOSine[4] , \LOSine[5] , \LOSine[6] , \LOSine[7] , \LOSine[8] , 
            \LOSine[9] , \LOSine[10] , \LOSine[11] , \LOSine[12] , \LOCosine[1] , 
            \LOCosine[2] , \LOCosine[3] , \LOCosine[4] , \LOCosine[5] , 
            \LOCosine[6] , \LOCosine[7] , \LOCosine[8] , \LOCosine[9] , 
            \LOCosine[10] , \LOCosine[11] , \LOCosine[12] , \phase_accum[56] ) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk_80mhz;
    input VCC_net;
    input GND_net;
    input \phase_accum[57] ;
    input \phase_accum[58] ;
    input \phase_accum[59] ;
    input \phase_accum[60] ;
    input \phase_accum[61] ;
    input \phase_accum[62] ;
    input \phase_accum[63] ;
    output \LOSine[1] ;
    output \LOSine[2] ;
    output \LOSine[3] ;
    output \LOSine[4] ;
    output \LOSine[5] ;
    output \LOSine[6] ;
    output \LOSine[7] ;
    output \LOSine[8] ;
    output \LOSine[9] ;
    output \LOSine[10] ;
    output \LOSine[11] ;
    output \LOSine[12] ;
    output \LOCosine[1] ;
    output \LOCosine[2] ;
    output \LOCosine[3] ;
    output \LOCosine[4] ;
    output \LOCosine[5] ;
    output \LOCosine[6] ;
    output \LOCosine[7] ;
    output \LOCosine[8] ;
    output \LOCosine[9] ;
    output \LOCosine[10] ;
    output \LOCosine[11] ;
    output \LOCosine[12] ;
    input \phase_accum[56] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(61[23:32])
    
    wire rom_addr0_r_1, rom_addr0_r_1_inv, rom_addr0_r_2, rom_addr0_r_3, 
        rom_addr0_r_4, rom_addr0_r_5, mx_ctrl_r, mx_ctrl_r_1, rom_addr0_r, 
        rom_addr0_r_n, rom_addr0_r_6, rom_dout_11, rom_dout_11_ffin, 
        rom_dout_10, rom_dout_10_ffin, rom_dout_9, rom_dout_9_ffin, 
        rom_dout_8, rom_dout_8_ffin, rom_dout_7, rom_dout_7_ffin, rom_dout_6, 
        rom_dout_6_ffin, rom_dout_5, rom_dout_5_ffin, rom_dout_4, rom_dout_4_ffin, 
        rom_dout_3, rom_dout_3_ffin, rom_dout_2, rom_dout_2_ffin, rom_dout_1, 
        rom_dout_1_ffin, rom_dout, rom_dout_ffin, rom_dout_25, rom_dout_25_ffin, 
        rom_dout_24, rom_dout_24_ffin, rom_dout_23, rom_dout_23_ffin, 
        rom_dout_22, rom_dout_22_ffin, rom_dout_21, rom_dout_21_ffin, 
        rom_dout_20, rom_dout_20_ffin, rom_dout_19, rom_dout_19_ffin, 
        rom_dout_18, rom_dout_18_ffin, rom_dout_17, rom_dout_17_ffin, 
        rom_dout_16, rom_dout_16_ffin, rom_dout_15, rom_dout_15_ffin, 
        rom_dout_14, rom_dout_14_ffin, rom_dout_13, rom_dout_13_ffin, 
        cosromoutsel_i, cosromoutsel, sinromoutsel, sinout_pre_1, sinout_pre_2, 
        sinout_pre_3, sinout_pre_4, sinout_pre_5, sinout_pre_6, sinout_pre_7, 
        sinout_pre_8, sinout_pre_9, sinout_pre_10, sinout_pre_11, sinout_pre_12, 
        cosout_pre_1, cosout_pre_2, cosout_pre_3, cosout_pre_4, cosout_pre_5, 
        cosout_pre_6, cosout_pre_7, cosout_pre_8, cosout_pre_9, cosout_pre_10, 
        cosout_pre_11, cosout_pre_12, rom_addr0_r_inv, co0, rom_addr0_r_n_1, 
        rom_addr0_r_n_2, rom_addr0_r_2_inv, co1, rom_addr0_r_n_3, rom_addr0_r_n_4, 
        rom_addr0_r_4_inv, rom_addr0_r_3_inv, co2, rom_addr0_r_n_5, 
        rom_addr0_r_5_inv, rom_dout_12_ffin, rom_addr0_r_7, rom_addr0_r_8, 
        rom_addr0_r_9, rom_addr0_r_10, rom_addr0_r_11, rom_dout_s_n_1, 
        rom_dout_s_n_2, rom_dout_2_inv, rom_dout_1_inv, co0_1, co1_1, 
        rom_dout_s_n_3, rom_dout_s_n_4, rom_dout_4_inv, rom_dout_3_inv, 
        co2_1, rom_dout_s_n_5, rom_dout_s_n_6, rom_dout_6_inv, rom_dout_5_inv, 
        co3, rom_dout_s_n_7, rom_dout_s_n_8, rom_dout_8_inv, rom_dout_7_inv, 
        co4, rom_dout_s_n_9, rom_dout_s_n_10, rom_dout_10_inv, rom_dout_9_inv, 
        co5, rom_dout_s_n_11, rom_dout_s_n_12, rom_dout_12_inv, rom_dout_11_inv, 
        rom_dout_13_inv, co0_2, rom_dout_c_n_1, rom_dout_c_n_2, rom_dout_15_inv, 
        rom_dout_14_inv, co1_2, rom_dout_c_n_3, rom_dout_c_n_4, rom_dout_17_inv, 
        rom_dout_16_inv, co2_2, rom_dout_c_n_5, rom_dout_c_n_6, rom_dout_19_inv, 
        rom_dout_18_inv, co3_1, rom_dout_c_n_7, rom_dout_c_n_8, rom_dout_21_inv, 
        rom_dout_20_inv, co4_1, rom_dout_c_n_9, rom_dout_c_n_10, rom_dout_23_inv, 
        rom_dout_22_inv, co5_1, rom_dout_c_n_11, rom_dout_c_n_12, rom_dout_25_inv, 
        rom_dout_24_inv, rom_dout_12, rom_dout_inv, func_or_inet, lx_ne0, 
        lx_ne0_inv, out_sel_i, rom_dout_s_1, rom_dout_s_2, rom_dout_s_3, 
        rom_dout_s_4, rom_dout_s_5, rom_dout_s_6, rom_dout_s_7, rom_dout_s_8, 
        rom_dout_s_9, rom_dout_s_10, rom_dout_s_11, rom_dout_s_12, rom_dout_c_1, 
        rom_dout_c_2, rom_dout_c_3, rom_dout_c_4, rom_dout_c_5, rom_dout_c_6, 
        rom_dout_c_7, rom_dout_c_8, rom_dout_c_9, rom_dout_c_10, rom_dout_c_11, 
        rom_dout_c_12, out_sel;
    
    INV INV_29 (.A(rom_addr0_r_1), .Z(rom_addr0_r_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    FD1P3DX FF_61 (.D(\phase_accum[57] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(312[13:88])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(\phase_accum[58] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(315[13:88])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(\phase_accum[59] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(318[13:88])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(\phase_accum[60] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(321[13:88])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(\phase_accum[61] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(324[13:88])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(\phase_accum[62] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(mx_ctrl_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(327[13:84])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(\phase_accum[63] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(mx_ctrl_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(330[13:86])
    defparam FF_55.GSR = "ENABLED";
    MUX21 muxb_57 (.D0(rom_addr0_r), .D1(rom_addr0_r_n), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    FD1P3DX FF_53 (.D(rom_dout_11_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(355[13] 356[25])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rom_dout_10_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(359[13] 360[25])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(rom_dout_9_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(363[13] 364[24])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(rom_dout_8_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(367[13] 368[24])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(rom_dout_7_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(371[13] 372[24])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(rom_dout_6_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(375[13] 376[24])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(rom_dout_5_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(379[13] 380[24])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(rom_dout_4_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(383[13] 384[24])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(rom_dout_3_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(387[13] 388[24])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(rom_dout_2_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(391[13] 392[24])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(rom_dout_1_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(395[13] 396[24])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(rom_dout_ffin), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(rom_dout)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(399[13] 400[22])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(rom_dout_25_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_25)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(403[13] 404[25])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(rom_dout_24_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_24)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(407[13] 408[25])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(rom_dout_23_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(411[13] 412[25])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(rom_dout_22_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(415[13] 416[25])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(rom_dout_21_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(419[13] 420[25])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(rom_dout_20_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(423[13] 424[25])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(rom_dout_19_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(427[13] 428[25])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(rom_dout_18_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(431[13] 432[25])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(rom_dout_17_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(435[13] 436[25])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(rom_dout_16_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(439[13] 440[25])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(rom_dout_15_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(443[13] 444[25])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(rom_dout_14_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(447[13] 448[25])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(rom_dout_13_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(451[13] 452[25])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(cosromoutsel_i), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(cosromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(455[13] 456[26])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(mx_ctrl_r_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(sinromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(459[13] 460[26])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(sinout_pre_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(599[13] 600[21])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(sinout_pre_2), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(603[13] 604[21])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(sinout_pre_3), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(607[13] 608[21])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(sinout_pre_4), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(611[13] 612[21])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(sinout_pre_5), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(615[13] 616[21])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(sinout_pre_6), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(619[13] 620[21])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(sinout_pre_7), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(623[13] 624[21])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(sinout_pre_8), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(627[13] 628[21])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(sinout_pre_9), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(631[13] 632[21])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(sinout_pre_10), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(635[13] 636[22])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(sinout_pre_11), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(639[13] 640[22])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(sinout_pre_12), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOSine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(643[13] 644[22])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(cosout_pre_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(650[13] 651[23])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(cosout_pre_2), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(654[13] 655[23])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(cosout_pre_3), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(658[13] 659[23])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(cosout_pre_4), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(662[13] 663[23])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(cosout_pre_5), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(666[13] 667[23])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(cosout_pre_6), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(670[13] 671[23])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(cosout_pre_7), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(674[13] 675[23])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(cosout_pre_8), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(678[13] 679[23])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(cosout_pre_9), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(682[13] 683[23])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(cosout_pre_10), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(686[13] 687[24])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(cosout_pre_11), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(690[13] 691[24])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(cosout_pre_12), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\LOCosine[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(694[13] 695[24])
    defparam FF_0.GSR = "ENABLED";
    CCU2C neg_rom_addr0_r_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0), .S1(rom_addr0_r_n)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(702[11] 704[71])
    defparam neg_rom_addr0_r_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_0.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_0.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_1 (.A0(rom_addr0_r_1_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_2_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0), .COUT(co1), .S0(rom_addr0_r_n_1), 
          .S1(rom_addr0_r_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(710[11] 713[42])
    defparam neg_rom_addr0_r_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_1.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_2 (.A0(rom_addr0_r_3_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_4_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1), .COUT(co2), .S0(rom_addr0_r_n_3), 
          .S1(rom_addr0_r_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(719[11] 722[42])
    defparam neg_rom_addr0_r_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_2.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_3 (.A0(rom_addr0_r_5_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co2), .S0(rom_addr0_r_n_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(728[11] 730[73])
    defparam neg_rom_addr0_r_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_3.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_3.INJECT1_1 = "NO";
    ROM64X1A triglut_1_0_25 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_12_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_25.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    CCU2C neg_rom_dout_s_n_1 (.A0(rom_dout_1_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_2_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0_1), .COUT(co1_1), .S0(rom_dout_s_n_1), 
          .S1(rom_dout_s_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(874[11] 877[43])
    defparam neg_rom_dout_s_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_1.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_2 (.A0(rom_dout_3_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_4_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1_1), .COUT(co2_1), .S0(rom_dout_s_n_3), 
          .S1(rom_dout_s_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(883[11] 886[43])
    defparam neg_rom_dout_s_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_2.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_3 (.A0(rom_dout_5_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_6_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co2_1), .COUT(co3), .S0(rom_dout_s_n_5), 
          .S1(rom_dout_s_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(892[11] 895[41])
    defparam neg_rom_dout_s_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_3.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_3.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_4 (.A0(rom_dout_7_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_8_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co3), .COUT(co4), .S0(rom_dout_s_n_7), 
          .S1(rom_dout_s_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(901[11] 904[41])
    defparam neg_rom_dout_s_n_4.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_4.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_4.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_4.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_5 (.A0(rom_dout_9_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_10_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co4), .COUT(co5), .S0(rom_dout_s_n_9), 
          .S1(rom_dout_s_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(910[11] 913[42])
    defparam neg_rom_dout_s_n_5.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_5.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_5.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_5.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_6 (.A0(rom_dout_11_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_12_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co5), .S0(rom_dout_s_n_11), .S1(rom_dout_s_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(919[11] 922[42])
    defparam neg_rom_dout_s_n_6.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_6.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_6.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_6.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_13_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(936[11] 938[72])
    defparam neg_rom_dout_c_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_0.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_0.INJECT1_1 = "NO";
    INV INV_30 (.A(rom_addr0_r_2), .Z(rom_addr0_r_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    CCU2C neg_rom_dout_c_n_1 (.A0(rom_dout_14_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_15_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0_2), .COUT(co1_2), .S0(rom_dout_c_n_1), 
          .S1(rom_dout_c_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(944[11] 947[43])
    defparam neg_rom_dout_c_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_1.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_2 (.A0(rom_dout_16_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_17_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1_2), .COUT(co2_2), .S0(rom_dout_c_n_3), 
          .S1(rom_dout_c_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(953[11] 956[43])
    defparam neg_rom_dout_c_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_2.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_3 (.A0(rom_dout_18_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_19_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co2_2), .COUT(co3_1), .S0(rom_dout_c_n_5), 
          .S1(rom_dout_c_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(962[11] 965[43])
    defparam neg_rom_dout_c_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_3.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_3.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_4 (.A0(rom_dout_20_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_21_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co3_1), .COUT(co4_1), .S0(rom_dout_c_n_7), 
          .S1(rom_dout_c_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(971[11] 974[43])
    defparam neg_rom_dout_c_n_4.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_4.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_4.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_4.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_5 (.A0(rom_dout_22_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_23_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co4_1), .COUT(co5_1), .S0(rom_dout_c_n_9), 
          .S1(rom_dout_c_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(980[11] 983[44])
    defparam neg_rom_dout_c_n_5.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_5.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_5.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_5.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_6 (.A0(rom_dout_24_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_25_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co5_1), .S0(rom_dout_c_n_11), .S1(rom_dout_c_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(989[11] 992[44])
    defparam neg_rom_dout_c_n_6.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_6.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_6.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_6.INJECT1_1 = "NO";
    INV INV_31 (.A(rom_addr0_r_3), .Z(rom_addr0_r_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_32 (.A(rom_addr0_r_4), .Z(rom_addr0_r_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_33 (.A(rom_addr0_r_5), .Z(rom_addr0_r_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_28 (.A(rom_addr0_r), .Z(rom_addr0_r_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    XOR2 XOR2_t1 (.A(mx_ctrl_r), .B(mx_ctrl_r_1), .Z(cosromoutsel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(241[10:70])
    INV INV_27 (.A(rom_dout_12), .Z(rom_dout_12_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_26 (.A(rom_dout_11), .Z(rom_dout_11_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_25 (.A(rom_dout_10), .Z(rom_dout_10_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_24 (.A(rom_dout_9), .Z(rom_dout_9_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_23 (.A(rom_dout_8), .Z(rom_dout_8_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_22 (.A(rom_dout_7), .Z(rom_dout_7_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_21 (.A(rom_dout_6), .Z(rom_dout_6_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_20 (.A(rom_dout_5), .Z(rom_dout_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_19 (.A(rom_dout_4), .Z(rom_dout_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_18 (.A(rom_dout_3), .Z(rom_dout_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_17 (.A(rom_dout_2), .Z(rom_dout_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_16 (.A(rom_dout_1), .Z(rom_dout_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_15 (.A(rom_dout), .Z(rom_dout_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_14 (.A(rom_dout_25), .Z(rom_dout_25_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_13 (.A(rom_dout_24), .Z(rom_dout_24_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_12 (.A(rom_dout_23), .Z(rom_dout_23_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_11 (.A(rom_dout_22), .Z(rom_dout_22_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_10 (.A(rom_dout_21), .Z(rom_dout_21_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_9 (.A(rom_dout_20), .Z(rom_dout_20_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_8 (.A(rom_dout_19), .Z(rom_dout_19_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_7 (.A(rom_dout_18), .Z(rom_dout_18_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_6 (.A(rom_dout_17), .Z(rom_dout_17_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_5 (.A(rom_dout_16), .Z(rom_dout_16_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_4 (.A(rom_dout_15), .Z(rom_dout_15_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_3 (.A(rom_dout_14), .Z(rom_dout_14_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    INV INV_2 (.A(rom_dout_13), .Z(rom_dout_13_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    ROM16X1A LUT4_1 (.AD0(rom_addr0_r_9), .AD1(rom_addr0_r_8), .AD2(rom_addr0_r_7), 
            .AD3(rom_addr0_r_6), .DO0(func_or_inet)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam LUT4_1.initval = 16'b1111111111111110;
    ROM16X1A LUT4_0 (.AD0(GND_net), .AD1(rom_addr0_r_11), .AD2(rom_addr0_r_10), 
            .AD3(func_or_inet), .DO0(lx_ne0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam LUT4_0.initval = 16'b1111111111111110;
    INV INV_1 (.A(lx_ne0), .Z(lx_ne0_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    AND2 AND2_t0 (.A(mx_ctrl_r), .B(lx_ne0_inv), .Z(out_sel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(305[10:64])
    FD1P3DX FF_62 (.D(\phase_accum[56] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(309[13:86])
    defparam FF_62.GSR = "ENABLED";
    MUX21 muxb_56 (.D0(rom_addr0_r_1), .D1(rom_addr0_r_n_1), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_55 (.D0(rom_addr0_r_2), .D1(rom_addr0_r_n_2), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_54 (.D0(rom_addr0_r_3), .D1(rom_addr0_r_n_3), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_53 (.D0(rom_addr0_r_4), .D1(rom_addr0_r_n_4), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_52 (.D0(rom_addr0_r_5), .D1(rom_addr0_r_n_5), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    FD1P3DX FF_54 (.D(rom_dout_12_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(351[13] 352[25])
    defparam FF_54.GSR = "ENABLED";
    MUX21 muxb_50 (.D0(rom_dout_1), .D1(rom_dout_s_n_1), .SD(sinromoutsel), 
          .Z(rom_dout_s_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_49 (.D0(rom_dout_2), .D1(rom_dout_s_n_2), .SD(sinromoutsel), 
          .Z(rom_dout_s_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_48 (.D0(rom_dout_3), .D1(rom_dout_s_n_3), .SD(sinromoutsel), 
          .Z(rom_dout_s_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_47 (.D0(rom_dout_4), .D1(rom_dout_s_n_4), .SD(sinromoutsel), 
          .Z(rom_dout_s_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_46 (.D0(rom_dout_5), .D1(rom_dout_s_n_5), .SD(sinromoutsel), 
          .Z(rom_dout_s_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_45 (.D0(rom_dout_6), .D1(rom_dout_s_n_6), .SD(sinromoutsel), 
          .Z(rom_dout_s_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_44 (.D0(rom_dout_7), .D1(rom_dout_s_n_7), .SD(sinromoutsel), 
          .Z(rom_dout_s_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_43 (.D0(rom_dout_8), .D1(rom_dout_s_n_8), .SD(sinromoutsel), 
          .Z(rom_dout_s_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_42 (.D0(rom_dout_9), .D1(rom_dout_s_n_9), .SD(sinromoutsel), 
          .Z(rom_dout_s_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_41 (.D0(rom_dout_10), .D1(rom_dout_s_n_10), .SD(sinromoutsel), 
          .Z(rom_dout_s_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_40 (.D0(rom_dout_11), .D1(rom_dout_s_n_11), .SD(sinromoutsel), 
          .Z(rom_dout_s_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_39 (.D0(rom_dout_12), .D1(rom_dout_s_n_12), .SD(sinromoutsel), 
          .Z(rom_dout_s_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_37 (.D0(rom_dout_14), .D1(rom_dout_c_n_1), .SD(cosromoutsel), 
          .Z(rom_dout_c_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_36 (.D0(rom_dout_15), .D1(rom_dout_c_n_2), .SD(cosromoutsel), 
          .Z(rom_dout_c_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_35 (.D0(rom_dout_16), .D1(rom_dout_c_n_3), .SD(cosromoutsel), 
          .Z(rom_dout_c_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_34 (.D0(rom_dout_17), .D1(rom_dout_c_n_4), .SD(cosromoutsel), 
          .Z(rom_dout_c_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_33 (.D0(rom_dout_18), .D1(rom_dout_c_n_5), .SD(cosromoutsel), 
          .Z(rom_dout_c_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_32 (.D0(rom_dout_19), .D1(rom_dout_c_n_6), .SD(cosromoutsel), 
          .Z(rom_dout_c_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_31 (.D0(rom_dout_20), .D1(rom_dout_c_n_7), .SD(cosromoutsel), 
          .Z(rom_dout_c_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_30 (.D0(rom_dout_21), .D1(rom_dout_c_n_8), .SD(cosromoutsel), 
          .Z(rom_dout_c_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_29 (.D0(rom_dout_22), .D1(rom_dout_c_n_9), .SD(cosromoutsel), 
          .Z(rom_dout_c_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_28 (.D0(rom_dout_23), .D1(rom_dout_c_n_10), .SD(cosromoutsel), 
          .Z(rom_dout_c_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_27 (.D0(rom_dout_24), .D1(rom_dout_c_n_11), .SD(cosromoutsel), 
          .Z(rom_dout_c_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_26 (.D0(rom_dout_25), .D1(rom_dout_c_n_12), .SD(cosromoutsel), 
          .Z(rom_dout_c_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    FD1P3DX FF_26 (.D(out_sel_i), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(out_sel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(541[13:83])
    defparam FF_26.GSR = "ENABLED";
    MUX21 muxb_24 (.D0(rom_dout_s_1), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_23 (.D0(rom_dout_s_2), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_22 (.D0(rom_dout_s_3), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_21 (.D0(rom_dout_s_4), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_20 (.D0(rom_dout_s_5), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_19 (.D0(rom_dout_s_6), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_18 (.D0(rom_dout_s_7), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_17 (.D0(rom_dout_s_8), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_16 (.D0(rom_dout_s_9), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_15 (.D0(rom_dout_s_10), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_14 (.D0(rom_dout_s_11), .D1(VCC_net), .SD(out_sel), .Z(sinout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_13 (.D0(rom_dout_s_12), .D1(mx_ctrl_r_1), .SD(out_sel), 
          .Z(sinout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_11 (.D0(rom_dout_c_1), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_10 (.D0(rom_dout_c_2), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_9 (.D0(rom_dout_c_3), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_8 (.D0(rom_dout_c_4), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_7 (.D0(rom_dout_c_5), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_6 (.D0(rom_dout_c_6), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_5 (.D0(rom_dout_c_7), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_4 (.D0(rom_dout_c_8), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_3 (.D0(rom_dout_c_9), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_2 (.D0(rom_dout_c_10), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_1 (.D0(rom_dout_c_11), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    MUX21 muxb_0 (.D0(rom_dout_c_12), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    ROM64X1A triglut_1_0_24 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_11_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_24.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_23 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_10_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_23.initval = 64'b1111111111111111111111111111111111111111110000000000000000000000;
    ROM64X1A triglut_1_0_22 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_9_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_22.initval = 64'b1111111111111111111111111111100000000000001111111111100000000000;
    ROM64X1A triglut_1_0_21 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_8_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_21.initval = 64'b1111111111111111111100000000011111110000001111110000011111000000;
    ROM64X1A triglut_1_0_20 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_7_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_20.initval = 64'b1111111111111100000011111000011110001110001110001110011100111000;
    ROM64X1A triglut_1_0_19 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_6_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_19.initval = 64'b1111111111000011100011100110011001001101101101001001011010110100;
    ROM64X1A triglut_1_0_18 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_5_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_18.initval = 64'b1111111000110011011010010101010100101001001001101100110001100110;
    ROM64X1A triglut_1_0_17 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_4_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_17.initval = 64'b1111100100101010110011000000000001110011011010110101010110101010;
    ROM64X1A triglut_1_0_16 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_3_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_16.initval = 64'b1110010110011100010101001111111101101010110011100000000011110000;
    ROM64X1A triglut_1_0_15 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_2_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_15.initval = 64'b1101000010100011001111010111110011001100010101100000000011001100;
    ROM64X1A triglut_1_0_14 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_1_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_14.initval = 64'b1111011011100010010110111011101001110011000000100111110010101010;
    ROM64X1A triglut_1_0_13 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_13.initval = 64'b1000100101001010011001010111111001010010011110001001001001111000;
    ROM64X1A triglut_1_0_12 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_25_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_12.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_11 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_24_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_11.initval = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    ROM64X1A triglut_1_0_10 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_23_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_10.initval = 64'b0000000000000000000001111111111111111111111111111111111111111110;
    ROM64X1A triglut_1_0_9 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_22_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_9.initval = 64'b0000000000111111111110000000000000111111111111111111111111111110;
    ROM64X1A triglut_1_0_8 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_21_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_8.initval = 64'b0000011111000001111110000001111111000000000111111111111111111110;
    ROM64X1A triglut_1_0_7 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_20_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_7.initval = 64'b0011100111001110001110001110001111000011111000000111111111111110;
    ROM64X1A triglut_1_0_6 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_19_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_6.initval = 64'b0101101011010010010110110110010011001100111000111000011111111110;
    ROM64X1A triglut_1_0_5 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_18_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_5.initval = 64'b1100110001100110110010010010100101010101001011011001100011111110;
    ROM64X1A triglut_1_0_4 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_17_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_4.initval = 64'b1010101101010101101011011001110000000000011001101010100100111110;
    ROM64X1A triglut_1_0_3 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_16_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_3.initval = 64'b0001111000000000111001101010110111111110010101000111001101001110;
    ROM64X1A triglut_1_0_2 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_15_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_2.initval = 64'b0110011000000000110101000110011001111101011110011000101000010110;
    ROM64X1A triglut_1_0_1 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_14_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_1.initval = 64'b1010101001111100100000011001110010111011101101001000111011011110;
    ROM64X1A triglut_1_0_0 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_13_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(102[11] 109[5])
    defparam triglut_1_0_0.initval = 64'b0011110010010010001111001001010011111101010011001010010100100010;
    CCU2C neg_rom_dout_s_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=5, LSE_LLINE=102, LSE_RLINE=109 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/IP/SinCos/SinCos.v(866[11] 868[72])
    defparam neg_rom_dout_s_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_0.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_0.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PLL
//

module PLL (clk_25mhz_c, clk_80mhz, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk_25mhz_c;
    output clk_80mhz;
    input GND_net;
    
    wire clk_25mhz_c /* synthesis is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(40[22:31])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(61[23:32])
    
    EHXPLLL PLLInst_0 (.CLKI(clk_25mhz_c), .CLKFB(clk_80mhz), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .PHASELOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .CLKOP(clk_80mhz)) /* synthesis FREQUENCY_PIN_CLKOP="83.333333", FREQUENCY_PIN_CLKI="25.000000", ICP_CURRENT="5", LPF_RESISTOR="16", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=8, LSE_RCOL=5, LSE_LLINE=97, LSE_RLINE=100 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(97[8] 100[5])
    defparam PLLInst_0.CLKI_DIV = 3;
    defparam PLLInst_0.CLKFB_DIV = 10;
    defparam PLLInst_0.CLKOP_DIV = 7;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 6;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.CLKOP_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.PLL_LOCK_DELAY = 200;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.REFIN_RESET = "DISABLED";
    defparam PLLInst_0.SYNC_ENABLE = "DISABLED";
    defparam PLLInst_0.INT_LOCK_STICKY = "ENABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module \CIC(WIDTH=72,DECIMATION_RATIO=4096) 
//

module \CIC(WIDTH=72,DECIMATION_RATIO=4096)  (d_tmp, clk_80mhz, d5, d_d_tmp, 
            d2, d2_71__N_490, d3, d3_71__N_562, d4, d4_71__N_634, 
            d5_71__N_706, d6, d6_71__N_1459, d_d6, d7, d7_71__N_1531, 
            d_d7, d8, d8_71__N_1603, d_d8, d9, d9_71__N_1675, d_d9, 
            n19, CIC1_outCos, d1, d1_71__N_418, n22, n8, n37, 
            n11, n10, n13, count, n31, \CICGain[0] , n66, n18, 
            n30, n21, n3, n2, n5, n4, n7, n6, n9, n8_adj_127, 
            n15, n14, \CICGain[1] , \d10[68] , \d10[69] , \d10[67] , 
            n11_adj_128, n10_adj_129, n13_adj_130, n12, n63, n131, 
            \d_out_11__N_1819[2] , n64, n132, \d_out_11__N_1819[3] , 
            n65, n133, \d_out_11__N_1819[4] , n66_adj_131, n134, \d_out_11__N_1819[5] , 
            \d10[66] , n135, \d_out_11__N_1819[6] , n12_adj_132, \d10[67]_adj_133 , 
            n136, \d_out_11__N_1819[7] , n63_adj_134, n131_adj_135, 
            n15_adj_136, n64_adj_137, n132_adj_138, n65_adj_139, n133_adj_140, 
            n134_adj_141, n135_adj_142, n136_adj_143, n36, n25, n24, 
            n25_adj_144, n33, n24_adj_145, n27, n27_adj_146, n26, 
            n32, n14_adj_147, n35, \d10[60] , n26_adj_148, n34, 
            n17, \d10[59] , \d10[61] , \d10[62] , \d10[63] , \d10[64] , 
            \d10[70] , \d10[71] , \d_out_11__N_1819[10] , \d_out_11__N_1819[11] , 
            n20, n29, n16, n37_adj_149, n29_adj_150, n17610, \d10[65] , 
            \d10[68]_adj_151 , n87_adj_252, n28, n31_adj_155, n17630, 
            n19_adj_156, n28_adj_157, n18_adj_158, n21_adj_159, n20_adj_160, 
            n36_adj_161, n30_adj_162, n37_adj_163, n36_adj_164, n3_adj_165, 
            n2_adj_166, n5_adj_167, n4_adj_168, n7_adj_169, n6_adj_170, 
            n9_adj_171, n8_adj_172, n11_adj_173, n10_adj_174, n35_adj_175, 
            n13_adj_176, n12_adj_177, n15_adj_178, n14_adj_179, n17_adj_180, 
            n34_adj_181, n16_adj_182, n19_adj_183, n18_adj_184, n21_adj_185, 
            n20_adj_186, n23, n22_adj_187, n23_adj_188, n25_adj_189, 
            n24_adj_190, n27_adj_191, n26_adj_192, n29_adj_193, n28_adj_194, 
            n3_adj_195, n2_adj_196, n5_adj_197, n31_adj_198, n4_adj_199, 
            n7_adj_200, n6_adj_201, n9_adj_202, n8_adj_203, n30_adj_204, 
            n33_adj_205, n32_adj_206, n35_adj_207, n34_adj_208, n37_adj_209, 
            n36_adj_210, n17_adj_211, n16_adj_212, n11_adj_213, n10_adj_214, 
            n13_adj_215, n12_adj_216, n15_adj_217, n14_adj_218, n17_adj_219, 
            n16_adj_220, n19_adj_221, n18_adj_222, n21_adj_223, n23_adj_224, 
            n22_adj_225, n20_adj_226, n23_adj_227, n22_adj_228, n25_adj_229, 
            n24_adj_230, n27_adj_231, n26_adj_232, n29_adj_233, \d_out_11__N_1819[8] , 
            n28_adj_234, n31_adj_235, n30_adj_236, n118, n120, cout, 
            n115, n117, n112, n114, n109, n111, n33_adj_237, n32_adj_238, 
            n106, n108, n103, n105, n100, n102, n97, n99, n94, 
            n96, n91, n93, n88, n90, n35_adj_239, n85, n87, 
            n82, n84, n79, n81_adj_240, n76, n78_adj_241, n34_adj_242, 
            n33_adj_243, n32_adj_244, n3_adj_245, n2_adj_246, n5_adj_247, 
            n4_adj_248, n7_adj_249, n6_adj_250, n9_adj_251) /* synthesis syn_module_defined=1 */ ;
    output [71:0]d_tmp;
    input clk_80mhz;
    output [71:0]d5;
    output [71:0]d_d_tmp;
    output [71:0]d2;
    input [71:0]d2_71__N_490;
    output [71:0]d3;
    input [71:0]d3_71__N_562;
    output [71:0]d4;
    input [71:0]d4_71__N_634;
    input [71:0]d5_71__N_706;
    output [71:0]d6;
    input [71:0]d6_71__N_1459;
    output [71:0]d_d6;
    output [71:0]d7;
    input [71:0]d7_71__N_1531;
    output [71:0]d_d7;
    output [71:0]d8;
    input [71:0]d8_71__N_1603;
    output [71:0]d_d8;
    output [71:0]d9;
    input [71:0]d9_71__N_1675;
    output [71:0]d_d9;
    output n19;
    output [11:0]CIC1_outCos;
    output [71:0]d1;
    input [71:0]d1_71__N_418;
    output n22;
    output n8;
    output n37;
    output n11;
    output n10;
    output n13;
    output [15:0]count;
    output n31;
    input \CICGain[0] ;
    output n66;
    output n18;
    output n30;
    output n21;
    output n3;
    output n2;
    output n5;
    output n4;
    output n7;
    output n6;
    output n9;
    output n8_adj_127;
    output n15;
    output n14;
    input \CICGain[1] ;
    output \d10[68] ;
    output \d10[69] ;
    output \d10[67] ;
    output n11_adj_128;
    output n10_adj_129;
    output n13_adj_130;
    output n12;
    input n63;
    input n131;
    output \d_out_11__N_1819[2] ;
    input n64;
    input n132;
    output \d_out_11__N_1819[3] ;
    input n65;
    input n133;
    output \d_out_11__N_1819[4] ;
    input n66_adj_131;
    input n134;
    output \d_out_11__N_1819[5] ;
    input \d10[66] ;
    input n135;
    output \d_out_11__N_1819[6] ;
    output n12_adj_132;
    input \d10[67]_adj_133 ;
    input n136;
    output \d_out_11__N_1819[7] ;
    output n63_adj_134;
    input n131_adj_135;
    output n15_adj_136;
    output n64_adj_137;
    input n132_adj_138;
    output n65_adj_139;
    input n133_adj_140;
    input n134_adj_141;
    input n135_adj_142;
    input n136_adj_143;
    output n36;
    output n25;
    output n24;
    output n25_adj_144;
    output n33;
    output n24_adj_145;
    output n27;
    output n27_adj_146;
    output n26;
    output n32;
    output n14_adj_147;
    output n35;
    output \d10[60] ;
    output n26_adj_148;
    output n34;
    output n17;
    output \d10[59] ;
    output \d10[61] ;
    output \d10[62] ;
    output \d10[63] ;
    output \d10[64] ;
    output \d10[70] ;
    output \d10[71] ;
    input \d_out_11__N_1819[10] ;
    input \d_out_11__N_1819[11] ;
    output n20;
    output n29;
    output n16;
    output n37_adj_149;
    output n29_adj_150;
    output n17610;
    input \d10[65] ;
    input \d10[68]_adj_151 ;
    input [15:0]n87_adj_252;
    output n28;
    output n31_adj_155;
    output n17630;
    output n19_adj_156;
    output n28_adj_157;
    output n18_adj_158;
    output n21_adj_159;
    output n20_adj_160;
    output n36_adj_161;
    output n30_adj_162;
    output n37_adj_163;
    output n36_adj_164;
    output n3_adj_165;
    output n2_adj_166;
    output n5_adj_167;
    output n4_adj_168;
    output n7_adj_169;
    output n6_adj_170;
    output n9_adj_171;
    output n8_adj_172;
    output n11_adj_173;
    output n10_adj_174;
    output n35_adj_175;
    output n13_adj_176;
    output n12_adj_177;
    output n15_adj_178;
    output n14_adj_179;
    output n17_adj_180;
    output n34_adj_181;
    output n16_adj_182;
    output n19_adj_183;
    output n18_adj_184;
    output n21_adj_185;
    output n20_adj_186;
    output n23;
    output n22_adj_187;
    output n23_adj_188;
    output n25_adj_189;
    output n24_adj_190;
    output n27_adj_191;
    output n26_adj_192;
    output n29_adj_193;
    output n28_adj_194;
    output n3_adj_195;
    output n2_adj_196;
    output n5_adj_197;
    output n31_adj_198;
    output n4_adj_199;
    output n7_adj_200;
    output n6_adj_201;
    output n9_adj_202;
    output n8_adj_203;
    output n30_adj_204;
    output n33_adj_205;
    output n32_adj_206;
    output n35_adj_207;
    output n34_adj_208;
    output n37_adj_209;
    output n36_adj_210;
    output n17_adj_211;
    output n16_adj_212;
    output n11_adj_213;
    output n10_adj_214;
    output n13_adj_215;
    output n12_adj_216;
    output n15_adj_217;
    output n14_adj_218;
    output n17_adj_219;
    output n16_adj_220;
    output n19_adj_221;
    output n18_adj_222;
    output n21_adj_223;
    output n23_adj_224;
    output n22_adj_225;
    output n20_adj_226;
    output n23_adj_227;
    output n22_adj_228;
    output n25_adj_229;
    output n24_adj_230;
    output n27_adj_231;
    output n26_adj_232;
    output n29_adj_233;
    output \d_out_11__N_1819[8] ;
    output n28_adj_234;
    output n31_adj_235;
    output n30_adj_236;
    input n118;
    input n120;
    input cout;
    input n115;
    input n117;
    input n112;
    input n114;
    input n109;
    input n111;
    output n33_adj_237;
    output n32_adj_238;
    input n106;
    input n108;
    input n103;
    input n105;
    input n100;
    input n102;
    input n97;
    input n99;
    input n94;
    input n96;
    input n91;
    input n93;
    input n88;
    input n90;
    output n35_adj_239;
    input n85;
    input n87;
    input n82;
    input n84;
    input n79;
    input n81_adj_240;
    input n76;
    input n78_adj_241;
    output n34_adj_242;
    output n33_adj_243;
    output n32_adj_244;
    output n3_adj_245;
    output n2_adj_246;
    output n5_adj_247;
    output n4_adj_248;
    output n7_adj_249;
    output n6_adj_250;
    output n9_adj_251;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(61[23:32])
    
    wire clk_80mhz_enable_757, clk_80mhz_enable_797, v_comb;
    wire [71:0]d_out_11__N_1819;
    wire [15:0]count_15__N_1442;
    wire [71:0]d10;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[68:71])
    
    wire n17057, n17584, n17552, n17544, n18105, n17966, n17965, 
        n17969, n17968, n17975, count_15__N_1458, clk_80mhz_enable_847, 
        clk_80mhz_enable_897, clk_80mhz_enable_947, clk_80mhz_enable_997, 
        clk_80mhz_enable_1047, clk_80mhz_enable_1097, clk_80mhz_enable_1147, 
        clk_80mhz_enable_1197, clk_80mhz_enable_1247, clk_80mhz_enable_1297, 
        clk_80mhz_enable_1347, clk_80mhz_enable_1397;
    wire [71:0]d10_71__N_1747;
    
    wire n17974, n17978, n17977, n12708, n17981, n17980, n31_adj_2716, 
        n17511, n17515, n17513, n17574, n17495;
    
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    FD1S3AX d2_i0 (.D(d2_71__N_490[0]), .CK(clk_80mhz), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i0.GSR = "ENABLED";
    FD1S3AX d3_i0 (.D(d3_71__N_562[0]), .CK(clk_80mhz), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_634[0]), .CK(clk_80mhz), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_706[0]), .CK(clk_80mhz), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1459[0]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1531[0]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1603[0]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1675[0]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i55_1_lut (.A(d_d7[54]), .Z(n19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i55_1_lut.init = 16'h5555;
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1819[0]), .SP(clk_80mhz_enable_797), 
            .CK(clk_80mhz), .Q(CIC1_outCos[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_418[0]), .CK(clk_80mhz), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i0.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i52_1_lut (.A(d_d_tmp[51]), .Z(n22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i66_1_lut (.A(d_d_tmp[65]), .Z(n8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i37_1_lut (.A(d_d6[36]), .Z(n37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i63_1_lut (.A(d_d_tmp[62]), .Z(n11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i64_1_lut (.A(d_d_tmp[63]), .Z(n10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i61_1_lut (.A(d_d_tmp[60]), .Z(n13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i61_1_lut.init = 16'h5555;
    FD1S3IX count__i0 (.D(count_15__N_1442[0]), .CK(clk_80mhz), .CD(clk_80mhz_enable_757), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i0.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i43_1_lut (.A(d_d_tmp[42]), .Z(n31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i66_3_lut (.A(d10[65]), .B(d10[66]), .C(\CICGain[0] ), 
         .Z(n66)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i56_1_lut (.A(d_d7[55]), .Z(n18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i44_1_lut (.A(d_d_tmp[43]), .Z(n30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i53_1_lut (.A(d_d7[52]), .Z(n21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i71_1_lut (.A(d_d7[70]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i72_1_lut (.A(d_d7[71]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i69_1_lut (.A(d_d7[68]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i70_1_lut (.A(d_d7[69]), .Z(n4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i67_1_lut (.A(d_d7[66]), .Z(n7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i68_1_lut (.A(d_d7[67]), .Z(n6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 i6326_4_lut_rep_210 (.A(n17057), .B(n17584), .C(n17552), .D(n17544), 
         .Z(n18105)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i6326_4_lut_rep_210.init = 16'h4000;
    LUT4 i6326_4_lut_rep_211 (.A(n17057), .B(n17584), .C(n17552), .D(n17544), 
         .Z(clk_80mhz_enable_757)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i6326_4_lut_rep_211.init = 16'h4000;
    LUT4 sub_27_inv_0_i65_1_lut (.A(d_d7[64]), .Z(n9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i66_1_lut (.A(d_d7[65]), .Z(n8_adj_127)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i59_1_lut (.A(d_d7[58]), .Z(n15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i60_1_lut (.A(d_d7[59]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i210_3_lut_4_lut_then_3_lut (.A(\CICGain[1] ), .B(d10[66]), 
         .C(\d10[68] ), .Z(n17966)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i210_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 shift_right_31_i210_3_lut_4_lut_else_3_lut (.A(\CICGain[1] ), .B(\d10[69] ), 
         .C(\d10[67] ), .Z(n17965)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i210_3_lut_4_lut_else_3_lut.init = 16'he4e4;
    LUT4 sub_27_inv_0_i63_1_lut (.A(d_d7[62]), .Z(n11_adj_128)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i64_1_lut (.A(d_d7[63]), .Z(n10_adj_129)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i61_1_lut (.A(d_d7[60]), .Z(n13_adj_130)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i62_1_lut (.A(d_d7[61]), .Z(n12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i203_3_lut_4_lut (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(n63), .D(n131), .Z(\d_out_11__N_1819[2] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i203_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i204_3_lut_4_lut (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(n64), .D(n132), .Z(\d_out_11__N_1819[3] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i204_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i205_3_lut_4_lut (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(n65), .D(n133), .Z(\d_out_11__N_1819[4] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i205_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i206_3_lut_4_lut (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(n66_adj_131), .D(n134), .Z(\d_out_11__N_1819[5] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i206_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i207_3_lut_4_lut (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(\d10[66] ), .D(n135), .Z(\d_out_11__N_1819[6] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i207_3_lut_4_lut.init = 16'hfe10;
    LUT4 sub_25_inv_0_i62_1_lut (.A(d_d_tmp[61]), .Z(n12_adj_132)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i208_3_lut_4_lut (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(\d10[67]_adj_133 ), .D(n136), .Z(\d_out_11__N_1819[7] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i208_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i209_3_lut_4_lut_then_3_lut (.A(\CICGain[1] ), .B(d10[65]), 
         .C(\d10[67] ), .Z(n17969)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i209_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 shift_right_31_i203_3_lut_4_lut_adj_36 (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(n63_adj_134), .D(n131_adj_135), .Z(d_out_11__N_1819[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i203_3_lut_4_lut_adj_36.init = 16'hfe10;
    LUT4 shift_right_31_i209_3_lut_4_lut_else_3_lut (.A(\CICGain[1] ), .B(\d10[68] ), 
         .C(d10[66]), .Z(n17968)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i209_3_lut_4_lut_else_3_lut.init = 16'he4e4;
    LUT4 sub_25_inv_0_i59_1_lut (.A(d_d_tmp[58]), .Z(n15_adj_136)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i204_3_lut_4_lut_adj_37 (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(n64_adj_137), .D(n132_adj_138), .Z(d_out_11__N_1819[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i204_3_lut_4_lut_adj_37.init = 16'hfe10;
    LUT4 shift_right_31_i205_3_lut_4_lut_adj_38 (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(n65_adj_139), .D(n133_adj_140), .Z(d_out_11__N_1819[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i205_3_lut_4_lut_adj_38.init = 16'hfe10;
    LUT4 shift_right_31_i206_3_lut_4_lut_adj_39 (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(n66), .D(n134_adj_141), .Z(d_out_11__N_1819[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i206_3_lut_4_lut_adj_39.init = 16'hfe10;
    LUT4 shift_right_31_i207_3_lut_4_lut_adj_40 (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(d10[66]), .D(n135_adj_142), .Z(d_out_11__N_1819[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i207_3_lut_4_lut_adj_40.init = 16'hfe10;
    LUT4 shift_right_31_i208_3_lut_4_lut_adj_41 (.A(\CICGain[0] ), .B(\CICGain[1] ), 
         .C(\d10[67] ), .D(n136_adj_143), .Z(d_out_11__N_1819[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i208_3_lut_4_lut_adj_41.init = 16'hfe10;
    LUT4 sub_26_inv_0_i38_1_lut (.A(d_d6[37]), .Z(n36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i49_1_lut (.A(d_d7[48]), .Z(n25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i50_1_lut (.A(d_d7[49]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i49_1_lut (.A(d_d_tmp[48]), .Z(n25_adj_144)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i41_1_lut (.A(d_d_tmp[40]), .Z(n33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i50_1_lut (.A(d_d_tmp[49]), .Z(n24_adj_145)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i47_1_lut (.A(d_d7[46]), .Z(n27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i47_1_lut (.A(d_d_tmp[46]), .Z(n27_adj_146)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i48_1_lut (.A(d_d_tmp[47]), .Z(n26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i42_1_lut (.A(d_d_tmp[41]), .Z(n32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i60_1_lut (.A(d_d_tmp[59]), .Z(n14_adj_147)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i39_1_lut (.A(d_d_tmp[38]), .Z(n35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 i6393_then_3_lut (.A(\CICGain[1] ), .B(\d10[60] ), .C(d10[58]), 
         .Z(n17975)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6393_then_3_lut.init = 16'he4e4;
    LUT4 sub_27_inv_0_i48_1_lut (.A(d_d7[47]), .Z(n26_adj_148)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i40_1_lut (.A(d_d_tmp[39]), .Z(n34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i57_1_lut (.A(d_d_tmp[56]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i57_1_lut.init = 16'h5555;
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(count_15__N_1458), .CK(clk_80mhz), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(clk_80mhz_enable_797), .CK(clk_80mhz), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1S3AX d2_i1 (.D(d2_71__N_490[1]), .CK(clk_80mhz), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i1.GSR = "ENABLED";
    FD1S3AX d2_i2 (.D(d2_71__N_490[2]), .CK(clk_80mhz), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_490[3]), .CK(clk_80mhz), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_490[4]), .CK(clk_80mhz), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_490[5]), .CK(clk_80mhz), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_490[6]), .CK(clk_80mhz), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_490[7]), .CK(clk_80mhz), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_490[8]), .CK(clk_80mhz), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_490[9]), .CK(clk_80mhz), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_490[10]), .CK(clk_80mhz), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_490[11]), .CK(clk_80mhz), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_490[12]), .CK(clk_80mhz), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_490[13]), .CK(clk_80mhz), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_490[14]), .CK(clk_80mhz), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_490[15]), .CK(clk_80mhz), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_490[16]), .CK(clk_80mhz), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_490[17]), .CK(clk_80mhz), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_490[18]), .CK(clk_80mhz), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_490[19]), .CK(clk_80mhz), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_490[20]), .CK(clk_80mhz), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_490[21]), .CK(clk_80mhz), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_490[22]), .CK(clk_80mhz), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_490[23]), .CK(clk_80mhz), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_490[24]), .CK(clk_80mhz), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_490[25]), .CK(clk_80mhz), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_490[26]), .CK(clk_80mhz), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_490[27]), .CK(clk_80mhz), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_490[28]), .CK(clk_80mhz), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_490[29]), .CK(clk_80mhz), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_490[30]), .CK(clk_80mhz), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_490[31]), .CK(clk_80mhz), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_490[32]), .CK(clk_80mhz), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_490[33]), .CK(clk_80mhz), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_490[34]), .CK(clk_80mhz), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_490[35]), .CK(clk_80mhz), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_490[36]), .CK(clk_80mhz), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_490[37]), .CK(clk_80mhz), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_490[38]), .CK(clk_80mhz), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_490[39]), .CK(clk_80mhz), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_490[40]), .CK(clk_80mhz), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_490[41]), .CK(clk_80mhz), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_490[42]), .CK(clk_80mhz), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_490[43]), .CK(clk_80mhz), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_490[44]), .CK(clk_80mhz), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_490[45]), .CK(clk_80mhz), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_490[46]), .CK(clk_80mhz), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_490[47]), .CK(clk_80mhz), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_490[48]), .CK(clk_80mhz), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_490[49]), .CK(clk_80mhz), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_490[50]), .CK(clk_80mhz), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_490[51]), .CK(clk_80mhz), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_490[52]), .CK(clk_80mhz), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_490[53]), .CK(clk_80mhz), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_490[54]), .CK(clk_80mhz), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_490[55]), .CK(clk_80mhz), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_490[56]), .CK(clk_80mhz), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_490[57]), .CK(clk_80mhz), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_490[58]), .CK(clk_80mhz), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_490[59]), .CK(clk_80mhz), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_490[60]), .CK(clk_80mhz), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_490[61]), .CK(clk_80mhz), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_490[62]), .CK(clk_80mhz), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_490[63]), .CK(clk_80mhz), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_490[64]), .CK(clk_80mhz), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_490[65]), .CK(clk_80mhz), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_490[66]), .CK(clk_80mhz), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_490[67]), .CK(clk_80mhz), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_490[68]), .CK(clk_80mhz), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_490[69]), .CK(clk_80mhz), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_490[70]), .CK(clk_80mhz), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_490[71]), .CK(clk_80mhz), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_562[1]), .CK(clk_80mhz), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_562[2]), .CK(clk_80mhz), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_562[3]), .CK(clk_80mhz), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_562[4]), .CK(clk_80mhz), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_562[5]), .CK(clk_80mhz), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_562[6]), .CK(clk_80mhz), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_562[7]), .CK(clk_80mhz), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_562[8]), .CK(clk_80mhz), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_562[9]), .CK(clk_80mhz), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_562[10]), .CK(clk_80mhz), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_562[11]), .CK(clk_80mhz), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_562[12]), .CK(clk_80mhz), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_562[13]), .CK(clk_80mhz), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_562[14]), .CK(clk_80mhz), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_562[15]), .CK(clk_80mhz), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_562[16]), .CK(clk_80mhz), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_562[17]), .CK(clk_80mhz), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_562[18]), .CK(clk_80mhz), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_562[19]), .CK(clk_80mhz), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_562[20]), .CK(clk_80mhz), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_562[21]), .CK(clk_80mhz), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_562[22]), .CK(clk_80mhz), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_562[23]), .CK(clk_80mhz), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_562[24]), .CK(clk_80mhz), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_562[25]), .CK(clk_80mhz), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_562[26]), .CK(clk_80mhz), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_562[27]), .CK(clk_80mhz), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_562[28]), .CK(clk_80mhz), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_562[29]), .CK(clk_80mhz), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_562[30]), .CK(clk_80mhz), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_562[31]), .CK(clk_80mhz), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_562[32]), .CK(clk_80mhz), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_562[33]), .CK(clk_80mhz), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_562[34]), .CK(clk_80mhz), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_562[35]), .CK(clk_80mhz), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_562[36]), .CK(clk_80mhz), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_562[37]), .CK(clk_80mhz), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_562[38]), .CK(clk_80mhz), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_562[39]), .CK(clk_80mhz), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_562[40]), .CK(clk_80mhz), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_562[41]), .CK(clk_80mhz), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_562[42]), .CK(clk_80mhz), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_562[43]), .CK(clk_80mhz), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_562[44]), .CK(clk_80mhz), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_562[45]), .CK(clk_80mhz), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_562[46]), .CK(clk_80mhz), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_562[47]), .CK(clk_80mhz), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_562[48]), .CK(clk_80mhz), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_562[49]), .CK(clk_80mhz), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_562[50]), .CK(clk_80mhz), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_562[51]), .CK(clk_80mhz), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_562[52]), .CK(clk_80mhz), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_562[53]), .CK(clk_80mhz), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_562[54]), .CK(clk_80mhz), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_562[55]), .CK(clk_80mhz), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_562[56]), .CK(clk_80mhz), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_562[57]), .CK(clk_80mhz), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_562[58]), .CK(clk_80mhz), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_562[59]), .CK(clk_80mhz), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_562[60]), .CK(clk_80mhz), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_562[61]), .CK(clk_80mhz), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_562[62]), .CK(clk_80mhz), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_562[63]), .CK(clk_80mhz), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_562[64]), .CK(clk_80mhz), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_562[65]), .CK(clk_80mhz), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_562[66]), .CK(clk_80mhz), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_562[67]), .CK(clk_80mhz), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_562[68]), .CK(clk_80mhz), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_562[69]), .CK(clk_80mhz), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_562[70]), .CK(clk_80mhz), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_562[71]), .CK(clk_80mhz), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_634[1]), .CK(clk_80mhz), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_634[2]), .CK(clk_80mhz), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_634[3]), .CK(clk_80mhz), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_634[4]), .CK(clk_80mhz), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_634[5]), .CK(clk_80mhz), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_634[6]), .CK(clk_80mhz), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_634[7]), .CK(clk_80mhz), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_634[8]), .CK(clk_80mhz), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_634[9]), .CK(clk_80mhz), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_634[10]), .CK(clk_80mhz), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_634[11]), .CK(clk_80mhz), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_634[12]), .CK(clk_80mhz), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_634[13]), .CK(clk_80mhz), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_634[14]), .CK(clk_80mhz), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_634[15]), .CK(clk_80mhz), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_634[16]), .CK(clk_80mhz), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_634[17]), .CK(clk_80mhz), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_634[18]), .CK(clk_80mhz), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_634[19]), .CK(clk_80mhz), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_634[20]), .CK(clk_80mhz), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_634[21]), .CK(clk_80mhz), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_634[22]), .CK(clk_80mhz), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_634[23]), .CK(clk_80mhz), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_634[24]), .CK(clk_80mhz), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_634[25]), .CK(clk_80mhz), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_634[26]), .CK(clk_80mhz), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_634[27]), .CK(clk_80mhz), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_634[28]), .CK(clk_80mhz), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_634[29]), .CK(clk_80mhz), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_634[30]), .CK(clk_80mhz), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_634[31]), .CK(clk_80mhz), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_634[32]), .CK(clk_80mhz), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_634[33]), .CK(clk_80mhz), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_634[34]), .CK(clk_80mhz), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_634[35]), .CK(clk_80mhz), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_634[36]), .CK(clk_80mhz), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_634[37]), .CK(clk_80mhz), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_634[38]), .CK(clk_80mhz), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_634[39]), .CK(clk_80mhz), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_634[40]), .CK(clk_80mhz), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_634[41]), .CK(clk_80mhz), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_634[42]), .CK(clk_80mhz), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_634[43]), .CK(clk_80mhz), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_634[44]), .CK(clk_80mhz), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_634[45]), .CK(clk_80mhz), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_634[46]), .CK(clk_80mhz), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_634[47]), .CK(clk_80mhz), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_634[48]), .CK(clk_80mhz), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_634[49]), .CK(clk_80mhz), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_634[50]), .CK(clk_80mhz), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_634[51]), .CK(clk_80mhz), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_634[52]), .CK(clk_80mhz), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_634[53]), .CK(clk_80mhz), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_634[54]), .CK(clk_80mhz), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_634[55]), .CK(clk_80mhz), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_634[56]), .CK(clk_80mhz), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_634[57]), .CK(clk_80mhz), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_634[58]), .CK(clk_80mhz), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_634[59]), .CK(clk_80mhz), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_634[60]), .CK(clk_80mhz), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_634[61]), .CK(clk_80mhz), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_634[62]), .CK(clk_80mhz), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_634[63]), .CK(clk_80mhz), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_634[64]), .CK(clk_80mhz), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_634[65]), .CK(clk_80mhz), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_634[66]), .CK(clk_80mhz), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_634[67]), .CK(clk_80mhz), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_634[68]), .CK(clk_80mhz), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_634[69]), .CK(clk_80mhz), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_634[70]), .CK(clk_80mhz), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_634[71]), .CK(clk_80mhz), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_706[1]), .CK(clk_80mhz), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_706[2]), .CK(clk_80mhz), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_706[3]), .CK(clk_80mhz), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_706[4]), .CK(clk_80mhz), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_706[5]), .CK(clk_80mhz), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_706[6]), .CK(clk_80mhz), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_706[7]), .CK(clk_80mhz), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_706[8]), .CK(clk_80mhz), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_706[9]), .CK(clk_80mhz), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_706[10]), .CK(clk_80mhz), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_706[11]), .CK(clk_80mhz), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_706[12]), .CK(clk_80mhz), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_706[13]), .CK(clk_80mhz), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_706[14]), .CK(clk_80mhz), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_706[15]), .CK(clk_80mhz), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_706[16]), .CK(clk_80mhz), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_706[17]), .CK(clk_80mhz), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_706[18]), .CK(clk_80mhz), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_706[19]), .CK(clk_80mhz), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_706[20]), .CK(clk_80mhz), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_706[21]), .CK(clk_80mhz), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_706[22]), .CK(clk_80mhz), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_706[23]), .CK(clk_80mhz), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_706[24]), .CK(clk_80mhz), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_706[25]), .CK(clk_80mhz), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_706[26]), .CK(clk_80mhz), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_706[27]), .CK(clk_80mhz), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_706[28]), .CK(clk_80mhz), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_706[29]), .CK(clk_80mhz), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_706[30]), .CK(clk_80mhz), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_706[31]), .CK(clk_80mhz), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_706[32]), .CK(clk_80mhz), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_706[33]), .CK(clk_80mhz), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_706[34]), .CK(clk_80mhz), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_706[35]), .CK(clk_80mhz), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_706[36]), .CK(clk_80mhz), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_706[37]), .CK(clk_80mhz), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_706[38]), .CK(clk_80mhz), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_706[39]), .CK(clk_80mhz), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_706[40]), .CK(clk_80mhz), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_706[41]), .CK(clk_80mhz), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_706[42]), .CK(clk_80mhz), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_706[43]), .CK(clk_80mhz), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_706[44]), .CK(clk_80mhz), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_706[45]), .CK(clk_80mhz), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_706[46]), .CK(clk_80mhz), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_706[47]), .CK(clk_80mhz), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_706[48]), .CK(clk_80mhz), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_706[49]), .CK(clk_80mhz), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_706[50]), .CK(clk_80mhz), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_706[51]), .CK(clk_80mhz), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_706[52]), .CK(clk_80mhz), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_706[53]), .CK(clk_80mhz), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_706[54]), .CK(clk_80mhz), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_706[55]), .CK(clk_80mhz), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_706[56]), .CK(clk_80mhz), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_706[57]), .CK(clk_80mhz), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_706[58]), .CK(clk_80mhz), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_706[59]), .CK(clk_80mhz), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_706[60]), .CK(clk_80mhz), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_706[61]), .CK(clk_80mhz), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_706[62]), .CK(clk_80mhz), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_706[63]), .CK(clk_80mhz), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_706[64]), .CK(clk_80mhz), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_706[65]), .CK(clk_80mhz), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_706[66]), .CK(clk_80mhz), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_706[67]), .CK(clk_80mhz), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_706[68]), .CK(clk_80mhz), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_706[69]), .CK(clk_80mhz), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_706[70]), .CK(clk_80mhz), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_706[71]), .CK(clk_80mhz), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1459[1]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1459[2]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1459[3]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1459[4]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1459[5]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1459[6]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1459[7]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1459[8]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1459[9]), .SP(clk_80mhz_enable_847), .CK(clk_80mhz), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1459[10]), .SP(clk_80mhz_enable_847), 
            .CK(clk_80mhz), .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1459[11]), .SP(clk_80mhz_enable_847), 
            .CK(clk_80mhz), .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1459[12]), .SP(clk_80mhz_enable_847), 
            .CK(clk_80mhz), .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1459[13]), .SP(clk_80mhz_enable_847), 
            .CK(clk_80mhz), .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1459[14]), .SP(clk_80mhz_enable_847), 
            .CK(clk_80mhz), .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1459[15]), .SP(clk_80mhz_enable_847), 
            .CK(clk_80mhz), .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1459[16]), .SP(clk_80mhz_enable_847), 
            .CK(clk_80mhz), .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1459[17]), .SP(clk_80mhz_enable_847), 
            .CK(clk_80mhz), .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1459[18]), .SP(clk_80mhz_enable_847), 
            .CK(clk_80mhz), .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1459[19]), .SP(clk_80mhz_enable_847), 
            .CK(clk_80mhz), .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1459[20]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1459[21]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1459[22]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1459[23]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1459[24]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1459[25]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1459[26]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1459[27]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1459[28]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1459[29]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1459[30]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1459[31]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1459[32]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1459[33]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1459[34]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1459[35]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1459[36]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1459[37]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1459[38]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1459[39]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1459[40]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1459[41]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1459[42]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1459[43]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1459[44]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1459[45]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1459[46]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1459[47]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1459[48]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1459[49]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1459[50]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1459[51]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1459[52]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1459[53]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1459[54]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1459[55]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1459[56]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1459[57]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1459[58]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1459[59]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1459[60]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1459[61]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1459[62]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1459[63]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1459[64]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1459[65]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1459[66]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1459[67]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1459[68]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1459[69]), .SP(clk_80mhz_enable_897), 
            .CK(clk_80mhz), .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1459[70]), .SP(clk_80mhz_enable_947), 
            .CK(clk_80mhz), .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1459[71]), .SP(clk_80mhz_enable_947), 
            .CK(clk_80mhz), .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(clk_80mhz_enable_947), .CK(clk_80mhz), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1531[1]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1531[2]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1531[3]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1531[4]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1531[5]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1531[6]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1531[7]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1531[8]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1531[9]), .SP(clk_80mhz_enable_997), .CK(clk_80mhz), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1531[10]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1531[11]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1531[12]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1531[13]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1531[14]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1531[15]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1531[16]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1531[17]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1531[18]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1531[19]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1531[20]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1531[21]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1531[22]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1531[23]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1531[24]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1531[25]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1531[26]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1531[27]), .SP(clk_80mhz_enable_997), 
            .CK(clk_80mhz), .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1531[28]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1531[29]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1531[30]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1531[31]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1531[32]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1531[33]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1531[34]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1531[35]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1531[36]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1531[37]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1531[38]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1531[39]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1531[40]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1531[41]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1531[42]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1531[43]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1531[44]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1531[45]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1531[46]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1531[47]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1531[48]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1531[49]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1531[50]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1531[51]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1531[52]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1531[53]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1531[54]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1531[55]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1531[56]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1531[57]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1531[58]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1531[59]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1531[60]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1531[61]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1531[62]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1531[63]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1531[64]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1531[65]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1531[66]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1531[67]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1531[68]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1531[69]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1531[70]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1531[71]), .SP(clk_80mhz_enable_1047), 
            .CK(clk_80mhz), .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(clk_80mhz_enable_1047), .CK(clk_80mhz), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(clk_80mhz_enable_1047), .CK(clk_80mhz), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(clk_80mhz_enable_1047), .CK(clk_80mhz), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(clk_80mhz_enable_1047), .CK(clk_80mhz), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(clk_80mhz_enable_1047), .CK(clk_80mhz), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(clk_80mhz_enable_1047), .CK(clk_80mhz), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(clk_80mhz_enable_1097), .CK(clk_80mhz), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(clk_80mhz_enable_1147), .CK(clk_80mhz), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1603[1]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1603[2]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1603[3]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1603[4]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1603[5]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1603[6]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1603[7]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1603[8]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1603[9]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1603[10]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1603[11]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1603[12]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1603[13]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1603[14]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1603[15]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1603[16]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1603[17]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1603[18]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1603[19]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1603[20]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1603[21]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1603[22]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1603[23]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1603[24]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1603[25]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1603[26]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1603[27]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1603[28]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1603[29]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1603[30]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1603[31]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1603[32]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1603[33]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1603[34]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1603[35]), .SP(clk_80mhz_enable_1147), 
            .CK(clk_80mhz), .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1603[36]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1603[37]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1603[38]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1603[39]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1603[40]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1603[41]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1603[42]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1603[43]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1603[44]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1603[45]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1603[46]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1603[47]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1603[48]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1603[49]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1603[50]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1603[51]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1603[52]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1603[53]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1603[54]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1603[55]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1603[56]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1603[57]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1603[58]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1603[59]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1603[60]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1603[61]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1603[62]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1603[63]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1603[64]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1603[65]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1603[66]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1603[67]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1603[68]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1603[69]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1603[70]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1603[71]), .SP(clk_80mhz_enable_1197), 
            .CK(clk_80mhz), .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(clk_80mhz_enable_1197), .CK(clk_80mhz), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(clk_80mhz_enable_1247), .CK(clk_80mhz), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(clk_80mhz_enable_1297), .CK(clk_80mhz), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(clk_80mhz_enable_1297), .CK(clk_80mhz), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(clk_80mhz_enable_1297), .CK(clk_80mhz), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(clk_80mhz_enable_1297), .CK(clk_80mhz), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(clk_80mhz_enable_1297), .CK(clk_80mhz), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(clk_80mhz_enable_1297), .CK(clk_80mhz), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(clk_80mhz_enable_1297), .CK(clk_80mhz), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1675[1]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1675[2]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1675[3]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1675[4]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1675[5]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1675[6]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1675[7]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1675[8]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1675[9]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1675[10]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1675[11]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1675[12]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1675[13]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1675[14]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1675[15]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1675[16]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1675[17]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1675[18]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1675[19]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1675[20]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1675[21]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1675[22]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1675[23]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1675[24]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1675[25]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1675[26]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1675[27]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1675[28]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1675[29]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1675[30]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1675[31]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1675[32]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1675[33]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1675[34]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1675[35]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1675[36]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1675[37]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1675[38]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1675[39]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1675[40]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1675[41]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1675[42]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1675[43]), .SP(clk_80mhz_enable_1297), 
            .CK(clk_80mhz), .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1675[44]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1675[45]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1675[46]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1675[47]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1675[48]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1675[49]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1675[50]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1675[51]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1675[52]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1675[53]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1675[54]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1675[55]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1675[56]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1675[57]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1675[58]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1675[59]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1675[60]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1675[61]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1675[62]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1675[63]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1675[64]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1675[65]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1675[66]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1675[67]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1675[68]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1675[69]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1675[70]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1675[71]), .SP(clk_80mhz_enable_1347), 
            .CK(clk_80mhz), .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(clk_80mhz_enable_1347), .CK(clk_80mhz), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(clk_80mhz_enable_1397), .CK(clk_80mhz), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1747[57]), .SP(clk_80mhz_enable_1397), 
            .CK(clk_80mhz), .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1747[58]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1747[59]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1747[60]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1747[61]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[61] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1747[62]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[62] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1747[63]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[63] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1747[64]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[64] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1747[65]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1747[66]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1747[67]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[67] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1747[68]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[68] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1747[69]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[69] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1747[70]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[70] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1747[71]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[71] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1819[1]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(d_out_11__N_1819[2]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(d_out_11__N_1819[3]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(d_out_11__N_1819[4]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(d_out_11__N_1819[5]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(d_out_11__N_1819[6]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(d_out_11__N_1819[7]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(d_out_11__N_1819[8]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(d_out_11__N_1819[9]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(\d_out_11__N_1819[10] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(\d_out_11__N_1819[11] ), .SP(v_comb), .CK(clk_80mhz), 
            .Q(CIC1_outCos[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_418[1]), .CK(clk_80mhz), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_418[2]), .CK(clk_80mhz), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_418[3]), .CK(clk_80mhz), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_418[4]), .CK(clk_80mhz), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_418[5]), .CK(clk_80mhz), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_418[6]), .CK(clk_80mhz), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_418[7]), .CK(clk_80mhz), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_418[8]), .CK(clk_80mhz), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_418[9]), .CK(clk_80mhz), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_418[10]), .CK(clk_80mhz), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_418[11]), .CK(clk_80mhz), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_418[12]), .CK(clk_80mhz), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_418[13]), .CK(clk_80mhz), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_418[14]), .CK(clk_80mhz), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_418[15]), .CK(clk_80mhz), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_418[16]), .CK(clk_80mhz), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_418[17]), .CK(clk_80mhz), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_418[18]), .CK(clk_80mhz), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_418[19]), .CK(clk_80mhz), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_418[20]), .CK(clk_80mhz), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_418[21]), .CK(clk_80mhz), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_418[22]), .CK(clk_80mhz), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_418[23]), .CK(clk_80mhz), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_418[24]), .CK(clk_80mhz), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_418[25]), .CK(clk_80mhz), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_418[26]), .CK(clk_80mhz), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_418[27]), .CK(clk_80mhz), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_418[28]), .CK(clk_80mhz), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_418[29]), .CK(clk_80mhz), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_418[30]), .CK(clk_80mhz), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_418[31]), .CK(clk_80mhz), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_418[32]), .CK(clk_80mhz), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_418[33]), .CK(clk_80mhz), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_418[34]), .CK(clk_80mhz), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_418[35]), .CK(clk_80mhz), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_418[36]), .CK(clk_80mhz), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_418[37]), .CK(clk_80mhz), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_418[38]), .CK(clk_80mhz), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_418[39]), .CK(clk_80mhz), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_418[40]), .CK(clk_80mhz), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_418[41]), .CK(clk_80mhz), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_418[42]), .CK(clk_80mhz), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_418[43]), .CK(clk_80mhz), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_418[44]), .CK(clk_80mhz), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_418[45]), .CK(clk_80mhz), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_418[46]), .CK(clk_80mhz), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_418[47]), .CK(clk_80mhz), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_418[48]), .CK(clk_80mhz), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_418[49]), .CK(clk_80mhz), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_418[50]), .CK(clk_80mhz), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_418[51]), .CK(clk_80mhz), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_418[52]), .CK(clk_80mhz), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_418[53]), .CK(clk_80mhz), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_418[54]), .CK(clk_80mhz), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_418[55]), .CK(clk_80mhz), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_418[56]), .CK(clk_80mhz), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_418[57]), .CK(clk_80mhz), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_418[58]), .CK(clk_80mhz), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_418[59]), .CK(clk_80mhz), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_418[60]), .CK(clk_80mhz), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_418[61]), .CK(clk_80mhz), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_418[62]), .CK(clk_80mhz), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_418[63]), .CK(clk_80mhz), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_418[64]), .CK(clk_80mhz), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_418[65]), .CK(clk_80mhz), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_418[66]), .CK(clk_80mhz), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_418[67]), .CK(clk_80mhz), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_418[68]), .CK(clk_80mhz), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_418[69]), .CK(clk_80mhz), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_418[70]), .CK(clk_80mhz), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_418[71]), .CK(clk_80mhz), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i71.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i54_1_lut (.A(d_d7[53]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i45_1_lut (.A(d_d7[44]), .Z(n29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i58_1_lut (.A(d_d_tmp[57]), .Z(n16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i37_1_lut (.A(d_d_tmp[36]), .Z(n37_adj_149)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i45_1_lut (.A(d_d_tmp[44]), .Z(n29_adj_150)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 i6393_else_3_lut (.A(n17610), .B(\CICGain[1] ), .C(\d10[59] ), 
         .Z(n17974)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6393_else_3_lut.init = 16'he2e2;
    LUT4 shift_right_31_i209_3_lut_4_lut_then_3_lut_adj_42 (.A(\CICGain[1] ), 
         .B(\d10[65] ), .C(\d10[67]_adj_133 ), .Z(n17978)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i209_3_lut_4_lut_then_3_lut_adj_42.init = 16'hd8d8;
    LUT4 shift_right_31_i209_3_lut_4_lut_else_3_lut_adj_43 (.A(\CICGain[1] ), 
         .B(\d10[68]_adj_151 ), .C(\d10[66] ), .Z(n17977)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i209_3_lut_4_lut_else_3_lut_adj_43.init = 16'he4e4;
    FD1S3IX count__i2 (.D(n87_adj_252[2]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n87_adj_252[3]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n87_adj_252[4]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n87_adj_252[5]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n87_adj_252[6]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n87_adj_252[7]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n87_adj_252[8]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n87_adj_252[9]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n87_adj_252[10]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1442[11]), .CK(clk_80mhz), .CD(count_15__N_1458), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n87_adj_252[12]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n87_adj_252[13]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n87_adj_252[14]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n87_adj_252[15]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i15.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i46_1_lut (.A(d_d7[45]), .Z(n28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i43_1_lut (.A(d_d7[42]), .Z(n31_adj_155)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 i6390_then_3_lut (.A(\CICGain[1] ), .B(\d10[59] ), .C(d10[57]), 
         .Z(n17981)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6390_then_3_lut.init = 16'he4e4;
    LUT4 i6390_else_3_lut (.A(n17630), .B(\CICGain[1] ), .C(d10[58]), 
         .Z(n17980)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6390_else_3_lut.init = 16'he2e2;
    LUT4 sub_25_inv_0_i55_1_lut (.A(d_d_tmp[54]), .Z(n19_adj_156)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i46_1_lut (.A(d_d_tmp[45]), .Z(n28_adj_157)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i56_1_lut (.A(d_d_tmp[55]), .Z(n18_adj_158)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i53_1_lut (.A(d_d_tmp[52]), .Z(n21_adj_159)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i54_1_lut (.A(d_d_tmp[53]), .Z(n20_adj_160)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i61_rep_43_3_lut (.A(\d10[60] ), .B(\d10[61] ), 
         .C(\CICGain[0] ), .Z(n17630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i61_rep_43_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i38_1_lut (.A(d_d_tmp[37]), .Z(n36_adj_161)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i44_1_lut (.A(d_d7[43]), .Z(n30_adj_162)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 i3119_2_lut (.A(n87_adj_252[0]), .B(n31_adj_2716), .Z(count_15__N_1442[0])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(78[18] 81[12])
    defparam i3119_2_lut.init = 16'hbbbb;
    LUT4 sub_27_inv_0_i37_1_lut (.A(d_d7[36]), .Z(n37_adj_163)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i38_1_lut (.A(d_d7[37]), .Z(n36_adj_164)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i71_1_lut (.A(d_d8[70]), .Z(n3_adj_165)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 i1_4_lut (.A(n17511), .B(n17057), .C(n17515), .D(n17513), .Z(n31_adj_2716)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 sub_28_inv_0_i72_1_lut (.A(d_d8[71]), .Z(n2_adj_166)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i69_1_lut (.A(d_d8[68]), .Z(n5_adj_167)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i70_1_lut (.A(d_d8[69]), .Z(n4_adj_168)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i67_1_lut (.A(d_d8[66]), .Z(n7_adj_169)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i68_1_lut (.A(d_d8[67]), .Z(n6_adj_170)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i65_1_lut (.A(d_d8[64]), .Z(n9_adj_171)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i66_1_lut (.A(d_d8[65]), .Z(n8_adj_172)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i63_1_lut (.A(d_d8[62]), .Z(n11_adj_173)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i64_1_lut (.A(d_d8[63]), .Z(n10_adj_174)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i39_1_lut (.A(d_d7[38]), .Z(n35_adj_175)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i61_1_lut (.A(d_d8[60]), .Z(n13_adj_176)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i62_1_lut (.A(d_d8[61]), .Z(n12_adj_177)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i59_1_lut (.A(d_d8[58]), .Z(n15_adj_178)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i60_1_lut (.A(d_d8[59]), .Z(n14_adj_179)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i57_1_lut (.A(d_d8[56]), .Z(n17_adj_180)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i40_1_lut (.A(d_d7[39]), .Z(n34_adj_181)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i58_1_lut (.A(d_d8[57]), .Z(n16_adj_182)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i55_1_lut (.A(d_d8[54]), .Z(n19_adj_183)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i56_1_lut (.A(d_d8[55]), .Z(n18_adj_184)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i53_1_lut (.A(d_d8[52]), .Z(n21_adj_185)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i54_1_lut (.A(d_d8[53]), .Z(n20_adj_186)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i51_1_lut (.A(d_d8[50]), .Z(n23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i52_1_lut (.A(d_d8[51]), .Z(n22_adj_187)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i51_1_lut (.A(d_d_tmp[50]), .Z(n23_adj_188)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i49_1_lut (.A(d_d8[48]), .Z(n25_adj_189)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i50_1_lut (.A(d_d8[49]), .Z(n24_adj_190)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i47_1_lut (.A(d_d8[46]), .Z(n27_adj_191)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i48_1_lut (.A(d_d8[47]), .Z(n26_adj_192)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i45_1_lut (.A(d_d8[44]), .Z(n29_adj_193)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 i1_3_lut (.A(count[8]), .B(count[1]), .C(count[9]), .Z(n17511)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_44 (.A(count[10]), .B(count[6]), .C(count[7]), .D(count[5]), 
         .Z(n17515)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i1_4_lut_adj_44.init = 16'hfffe;
    LUT4 sub_28_inv_0_i46_1_lut (.A(d_d8[45]), .Z(n28_adj_194)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_45 (.A(count[2]), .B(count[4]), .C(count[0]), .D(count[3]), 
         .Z(n17513)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i1_4_lut_adj_45.init = 16'hfffe;
    LUT4 sub_26_inv_0_i71_1_lut (.A(d_d6[70]), .Z(n3_adj_195)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i72_1_lut (.A(d_d6[71]), .Z(n2_adj_196)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i69_1_lut (.A(d_d6[68]), .Z(n5_adj_197)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i43_1_lut (.A(d_d8[42]), .Z(n31_adj_198)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i70_1_lut (.A(d_d6[69]), .Z(n4_adj_199)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i67_1_lut (.A(d_d6[66]), .Z(n7_adj_200)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i68_1_lut (.A(d_d6[67]), .Z(n6_adj_201)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i65_1_lut (.A(d_d6[64]), .Z(n9_adj_202)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i66_1_lut (.A(d_d6[65]), .Z(n8_adj_203)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i44_1_lut (.A(d_d8[43]), .Z(n30_adj_204)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i41_1_lut (.A(d_d8[40]), .Z(n33_adj_205)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i42_1_lut (.A(d_d8[41]), .Z(n32_adj_206)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i39_1_lut (.A(d_d8[38]), .Z(n35_adj_207)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i40_1_lut (.A(d_d8[39]), .Z(n34_adj_208)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i37_1_lut (.A(d_d8[36]), .Z(n37_adj_209)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i38_1_lut (.A(d_d8[37]), .Z(n36_adj_210)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i57_1_lut (.A(d_d7[56]), .Z(n17_adj_211)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i58_1_lut (.A(d_d7[57]), .Z(n16_adj_212)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i63_1_lut (.A(d_d6[62]), .Z(n11_adj_213)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i64_1_lut (.A(d_d6[63]), .Z(n10_adj_214)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i61_1_lut (.A(d_d6[60]), .Z(n13_adj_215)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i62_1_lut (.A(d_d6[61]), .Z(n12_adj_216)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i59_1_lut (.A(d_d6[58]), .Z(n15_adj_217)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 i6326_4_lut (.A(n17057), .B(n17584), .C(n17552), .D(n17544), 
         .Z(count_15__N_1458)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i6326_4_lut.init = 16'h4000;
    LUT4 sub_26_inv_0_i60_1_lut (.A(d_d6[59]), .Z(n14_adj_218)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 i6258_2_lut (.A(count[5]), .B(count[8]), .Z(n17552)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6258_2_lut.init = 16'h8888;
    LUT4 sub_26_inv_0_i57_1_lut (.A(d_d6[56]), .Z(n17_adj_219)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i58_1_lut (.A(d_d6[57]), .Z(n16_adj_220)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i55_1_lut (.A(d_d6[54]), .Z(n19_adj_221)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i56_1_lut (.A(d_d6[55]), .Z(n18_adj_222)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 i6250_2_lut (.A(count[0]), .B(count[3]), .Z(n17544)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6250_2_lut.init = 16'h8888;
    LUT4 sub_26_inv_0_i53_1_lut (.A(d_d6[52]), .Z(n21_adj_223)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i51_1_lut (.A(d_d7[50]), .Z(n23_adj_224)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i52_1_lut (.A(d_d7[51]), .Z(n22_adj_225)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i54_1_lut (.A(d_d6[53]), .Z(n20_adj_226)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i51_1_lut (.A(d_d6[50]), .Z(n23_adj_227)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i52_1_lut (.A(d_d6[51]), .Z(n22_adj_228)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 i6280_4_lut (.A(count[2]), .B(count[4]), .C(count[1]), .D(count[6]), 
         .Z(n17574)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6280_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_46 (.A(count[12]), .B(count[11]), .C(n17495), .D(count[15]), 
         .Z(n17057)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_46.init = 16'hfffb;
    LUT4 i1_2_lut (.A(count[14]), .B(count[13]), .Z(n17495)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 sub_26_inv_0_i49_1_lut (.A(d_d6[48]), .Z(n25_adj_229)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i50_1_lut (.A(d_d6[49]), .Z(n24_adj_230)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i47_1_lut (.A(d_d6[46]), .Z(n27_adj_231)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 i6290_4_lut (.A(count[7]), .B(n17574), .C(count[9]), .D(count[10]), 
         .Z(n17584)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6290_4_lut.init = 16'h8000;
    LUT4 sub_26_inv_0_i48_1_lut (.A(d_d6[47]), .Z(n26_adj_232)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i48_1_lut.init = 16'h5555;
    PFUMX i6433 (.BLUT(n17980), .ALUT(n17981), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[0]));
    LUT4 sub_26_inv_0_i45_1_lut (.A(d_d6[44]), .Z(n29_adj_233)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i45_1_lut.init = 16'h5555;
    PFUMX i6431 (.BLUT(n17977), .ALUT(n17978), .C0(\CICGain[0] ), .Z(\d_out_11__N_1819[8] ));
    LUT4 sub_26_inv_0_i46_1_lut (.A(d_d6[45]), .Z(n28_adj_234)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i43_1_lut (.A(d_d6[42]), .Z(n31_adj_235)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i43_1_lut.init = 16'h5555;
    PFUMX i6429 (.BLUT(n17974), .ALUT(n17975), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[1]));
    LUT4 sub_26_inv_0_i44_1_lut (.A(d_d6[43]), .Z(n30_adj_236)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i44_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_225 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1397)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_225.GSR = "ENABLED";
    LUT4 mux_1249_i2_3_lut (.A(n118), .B(n120), .C(cout), .Z(d10_71__N_1747[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i2_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_224 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1347)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_224.GSR = "ENABLED";
    PFUMX i6425 (.BLUT(n17968), .ALUT(n17969), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[8]));
    LUT4 mux_1249_i3_3_lut (.A(n115), .B(n117), .C(cout), .Z(d10_71__N_1747[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i3_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_223 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1297)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_223.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_222 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1247)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_222.GSR = "ENABLED";
    LUT4 mux_1249_i4_3_lut (.A(n112), .B(n114), .C(cout), .Z(d10_71__N_1747[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i4_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_221 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1197)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_221.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_220 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1147)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_220.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_219 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1097)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_219.GSR = "ENABLED";
    LUT4 mux_1249_i5_3_lut (.A(n109), .B(n111), .C(cout), .Z(d10_71__N_1747[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i5_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i41_1_lut (.A(d_d6[40]), .Z(n33_adj_237)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i41_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_218 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1047)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_218.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i42_1_lut (.A(d_d6[41]), .Z(n32_adj_238)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i42_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_217 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_997)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_217.GSR = "ENABLED";
    LUT4 mux_1249_i6_3_lut (.A(n106), .B(n108), .C(cout), .Z(d10_71__N_1747[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1249_i7_3_lut (.A(n103), .B(n105), .C(cout), .Z(d10_71__N_1747[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1249_i8_3_lut (.A(n100), .B(n102), .C(cout), .Z(d10_71__N_1747[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i8_3_lut.init = 16'hcaca;
    FD1S3IX count__i1 (.D(n87_adj_252[1]), .CK(clk_80mhz), .CD(n12708), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i1.GSR = "ENABLED";
    LUT4 mux_1249_i9_3_lut (.A(n97), .B(n99), .C(cout), .Z(d10_71__N_1747[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1249_i10_3_lut (.A(n94), .B(n96), .C(cout), .Z(d10_71__N_1747[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i10_3_lut.init = 16'hcaca;
    PFUMX i6423 (.BLUT(n17965), .ALUT(n17966), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[9]));
    LUT4 mux_1249_i11_3_lut (.A(n91), .B(n93), .C(cout), .Z(d10_71__N_1747[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1249_i12_3_lut (.A(n88), .B(n90), .C(cout), .Z(d10_71__N_1747[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i12_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i39_1_lut (.A(d_d6[38]), .Z(n35_adj_239)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 mux_1249_i13_3_lut (.A(n85), .B(n87), .C(cout), .Z(d10_71__N_1747[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1249_i14_3_lut (.A(n82), .B(n84), .C(cout), .Z(d10_71__N_1747[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i14_3_lut.init = 16'hcaca;
    FD1S3AX v_comb_66_rep_216 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_947)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_216.GSR = "ENABLED";
    LUT4 mux_1249_i15_3_lut (.A(n79), .B(n81_adj_240), .C(cout), .Z(d10_71__N_1747[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1249_i16_3_lut (.A(n76), .B(n78_adj_241), .C(cout), .Z(d10_71__N_1747[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1249_i16_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i40_1_lut (.A(d_d6[39]), .Z(n34_adj_242)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 i6346_2_lut (.A(n31_adj_2716), .B(n18105), .Z(n12708)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam i6346_2_lut.init = 16'hdddd;
    LUT4 shift_right_31_i62_rep_23_3_lut (.A(\d10[61] ), .B(\d10[62] ), 
         .C(\CICGain[0] ), .Z(n17610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i62_rep_23_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i41_1_lut (.A(d_d7[40]), .Z(n33_adj_243)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i42_1_lut (.A(d_d7[41]), .Z(n32_adj_244)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 i3169_2_lut (.A(n87_adj_252[11]), .B(n31_adj_2716), .Z(count_15__N_1442[11])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(78[18] 81[12])
    defparam i3169_2_lut.init = 16'hbbbb;
    LUT4 sub_25_inv_0_i71_1_lut (.A(d_d_tmp[70]), .Z(n3_adj_245)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i71_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_215 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_897)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_215.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i72_1_lut (.A(d_d_tmp[71]), .Z(n2_adj_246)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i63_3_lut (.A(\d10[62] ), .B(\d10[63] ), .C(\CICGain[0] ), 
         .Z(n63_adj_134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i69_1_lut (.A(d_d_tmp[68]), .Z(n5_adj_247)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i69_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_214 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_847)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_214.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_213 (.D(clk_80mhz_enable_757), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_797)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=148, LSE_RLINE=154 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_213.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i70_1_lut (.A(d_d_tmp[69]), .Z(n4_adj_248)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i64_3_lut (.A(\d10[63] ), .B(\d10[64] ), .C(\CICGain[0] ), 
         .Z(n64_adj_137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i67_1_lut (.A(d_d_tmp[66]), .Z(n7_adj_249)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i68_1_lut (.A(d_d_tmp[67]), .Z(n6_adj_250)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i65_1_lut (.A(d_d_tmp[64]), .Z(n9_adj_251)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i65_3_lut (.A(\d10[64] ), .B(d10[65]), .C(\CICGain[0] ), 
         .Z(n65_adj_139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module nco_sig
//

module nco_sig (\phase_accum[63] , sinGen_c) /* synthesis syn_module_defined=1 */ ;
    input \phase_accum[63] ;
    output sinGen_c;
    
    
    LUT4 phase_accum_63__I_0_13_1_lut (.A(\phase_accum[63] ), .Z(sinGen_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/NCO.v(34[22:66])
    defparam phase_accum_63__I_0_13_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module AMDemodulator
//

module AMDemodulator (\DataInReg_11__N_1856[0] , CIC1_out_clkSin, CIC1_outCos, 
            MultResult2, \d_out_d_11__N_1880[17] , d_out_d_11__N_1879, 
            \d_out_d_11__N_1878[17] , d_out_d_11__N_1877, \d_out_d_11__N_1876[17] , 
            d_out_d_11__N_1875, MultDataB, MultResult1, VCC_net, GND_net, 
            \DataInReg_11__N_1856[1] , \DataInReg_11__N_1856[2] , \DataInReg_11__N_1856[3] , 
            \DataInReg_11__N_1856[4] , \DataInReg_11__N_1856[5] , \DataInReg_11__N_1856[6] , 
            \DataInReg_11__N_1856[7] , \DataInReg_11__N_1856[8] , \DemodOut[9] , 
            \d_out_d_11__N_2383[17] , \d_out_d_11__N_2401[17] , \d_out_d_11__N_1892[17] , 
            \ISquare[31] , n213, \d_out_d_11__N_1874[17] , d_out_d_11__N_1873, 
            \d_out_d_11__N_1888[17] , \d_out_d_11__N_1890[17] , \d_out_d_11__N_1886[17] , 
            \d_out_d_11__N_1884[17] , \d_out_d_11__N_1882[17] ) /* synthesis syn_module_defined=1 */ ;
    output \DataInReg_11__N_1856[0] ;
    input CIC1_out_clkSin;
    input [11:0]CIC1_outCos;
    output [23:0]MultResult2;
    input \d_out_d_11__N_1880[17] ;
    output d_out_d_11__N_1879;
    input \d_out_d_11__N_1878[17] ;
    output d_out_d_11__N_1877;
    input \d_out_d_11__N_1876[17] ;
    output d_out_d_11__N_1875;
    input [11:0]MultDataB;
    output [23:0]MultResult1;
    input VCC_net;
    input GND_net;
    output \DataInReg_11__N_1856[1] ;
    output \DataInReg_11__N_1856[2] ;
    output \DataInReg_11__N_1856[3] ;
    output \DataInReg_11__N_1856[4] ;
    output \DataInReg_11__N_1856[5] ;
    output \DataInReg_11__N_1856[6] ;
    output \DataInReg_11__N_1856[7] ;
    output \DataInReg_11__N_1856[8] ;
    output \DemodOut[9] ;
    input \d_out_d_11__N_2383[17] ;
    input \d_out_d_11__N_2401[17] ;
    input \d_out_d_11__N_1892[17] ;
    input \ISquare[31] ;
    output n213;
    input \d_out_d_11__N_1874[17] ;
    output d_out_d_11__N_1873;
    input \d_out_d_11__N_1888[17] ;
    input \d_out_d_11__N_1890[17] ;
    input \d_out_d_11__N_1886[17] ;
    input \d_out_d_11__N_1884[17] ;
    input \d_out_d_11__N_1882[17] ;
    
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(74[23:38])
    wire [15:0]d_out_d;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(30[28:35])
    wire [12:0]n27;
    wire [25:0]n83;
    wire [17:0]d_out_d_11__N_1894;
    
    wire d_out_d_11__N_1891, d_out_d_11__N_1889, d_out_d_11__N_1887, d_out_d_11__N_1885, 
        d_out_d_11__N_1883, d_out_d_11__N_1881;
    
    FD1S3AX d_out_i1 (.D(d_out_d[0]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i1.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i1 (.D(CIC1_outCos[0]), .CK(CIC1_out_clkSin), 
            .Q(n27[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i1.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i0 (.D(n83[0]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i0.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i1 (.D(d_out_d_11__N_1894[17]), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i1.GSR = "ENABLED";
    LUT4 d_out_d_11__I_4_1_lut (.A(\d_out_d_11__N_1880[17] ), .Z(d_out_d_11__N_1879)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_4_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_3_1_lut (.A(\d_out_d_11__N_1878[17] ), .Z(d_out_d_11__N_1877)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_3_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_2_1_lut (.A(\d_out_d_11__N_1876[17] ), .Z(d_out_d_11__N_1875)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_2_1_lut.init = 16'h5555;
    MULT18X18D MultResult1_e3 (.A17(MultDataB[11]), .A16(MultDataB[11]), 
            .A15(MultDataB[11]), .A14(MultDataB[11]), .A13(MultDataB[11]), 
            .A12(MultDataB[11]), .A11(MultDataB[11]), .A10(MultDataB[10]), 
            .A9(MultDataB[9]), .A8(MultDataB[8]), .A7(MultDataB[7]), .A6(MultDataB[6]), 
            .A5(MultDataB[5]), .A4(MultDataB[4]), .A3(MultDataB[3]), .A2(MultDataB[2]), 
            .A1(MultDataB[1]), .A0(MultDataB[0]), .B17(MultDataB[11]), 
            .B16(MultDataB[11]), .B15(MultDataB[11]), .B14(MultDataB[11]), 
            .B13(MultDataB[11]), .B12(MultDataB[11]), .B11(MultDataB[11]), 
            .B10(MultDataB[10]), .B9(MultDataB[9]), .B8(MultDataB[8]), 
            .B7(MultDataB[7]), .B6(MultDataB[6]), .B5(MultDataB[5]), .B4(MultDataB[4]), 
            .B3(MultDataB[3]), .B2(MultDataB[2]), .B1(MultDataB[1]), .B0(MultDataB[0]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(CIC1_out_clkSin), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(VCC_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .P23(MultResult1[23]), 
            .P22(MultResult1[22]), .P21(MultResult1[21]), .P20(MultResult1[20]), 
            .P19(MultResult1[19]), .P18(MultResult1[18]), .P17(MultResult1[17]), 
            .P16(MultResult1[16]), .P15(MultResult1[15]), .P14(MultResult1[14]), 
            .P13(MultResult1[13]), .P12(MultResult1[12]), .P11(MultResult1[11]), 
            .P10(MultResult1[10]), .P9(MultResult1[9]), .P8(MultResult1[8]), 
            .P7(MultResult1[7]), .P6(MultResult1[6]), .P5(MultResult1[5]), 
            .P4(MultResult1[4]), .P3(MultResult1[3]), .P2(MultResult1[2]), 
            .P1(MultResult1[1]), .P0(MultResult1[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(86[20:39])
    defparam MultResult1_e3.REG_INPUTA_CLK = "CLK3";
    defparam MultResult1_e3.REG_INPUTA_CE = "CE3";
    defparam MultResult1_e3.REG_INPUTA_RST = "RST3";
    defparam MultResult1_e3.REG_INPUTB_CLK = "CLK3";
    defparam MultResult1_e3.REG_INPUTB_CE = "CE3";
    defparam MultResult1_e3.REG_INPUTB_RST = "RST3";
    defparam MultResult1_e3.REG_INPUTC_CLK = "NONE";
    defparam MultResult1_e3.REG_INPUTC_CE = "CE0";
    defparam MultResult1_e3.REG_INPUTC_RST = "RST0";
    defparam MultResult1_e3.REG_PIPELINE_CLK = "NONE";
    defparam MultResult1_e3.REG_PIPELINE_CE = "CE0";
    defparam MultResult1_e3.REG_PIPELINE_RST = "RST0";
    defparam MultResult1_e3.REG_OUTPUT_CLK = "CLK3";
    defparam MultResult1_e3.REG_OUTPUT_CE = "CE3";
    defparam MultResult1_e3.REG_OUTPUT_RST = "RST3";
    defparam MultResult1_e3.CLK0_DIV = "ENABLED";
    defparam MultResult1_e3.CLK1_DIV = "ENABLED";
    defparam MultResult1_e3.CLK2_DIV = "ENABLED";
    defparam MultResult1_e3.CLK3_DIV = "ENABLED";
    defparam MultResult1_e3.HIGHSPEED_CLK = "NONE";
    defparam MultResult1_e3.GSR = "ENABLED";
    defparam MultResult1_e3.CAS_MATCH_REG = "FALSE";
    defparam MultResult1_e3.SOURCEB_MODE = "B_SHIFT";
    defparam MultResult1_e3.MULT_BYPASS = "DISABLED";
    defparam MultResult1_e3.RESETMODE = "ASYNC";
    MULT18X18D MultResult2_res2_mult_2 (.A17(n27[12]), .A16(n27[12]), .A15(n27[12]), 
            .A14(n27[12]), .A13(n27[12]), .A12(n27[12]), .A11(n27[12]), 
            .A10(n27[10]), .A9(n27[9]), .A8(n27[8]), .A7(n27[7]), .A6(n27[6]), 
            .A5(n27[5]), .A4(n27[4]), .A3(n27[3]), .A2(n27[2]), .A1(n27[1]), 
            .A0(n27[0]), .B17(n27[12]), .B16(n27[12]), .B15(n27[12]), 
            .B14(n27[12]), .B13(n27[12]), .B12(n27[12]), .B11(n27[12]), 
            .B10(n27[10]), .B9(n27[9]), .B8(n27[8]), .B7(n27[7]), .B6(n27[6]), 
            .B5(n27[5]), .B4(n27[4]), .B3(n27[3]), .B2(n27[2]), .B1(n27[1]), 
            .B0(n27[0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), 
            .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .P23(n83[23]), 
            .P22(n83[22]), .P21(n83[21]), .P20(n83[20]), .P19(n83[19]), 
            .P18(n83[18]), .P17(n83[17]), .P16(n83[16]), .P15(n83[15]), 
            .P14(n83[14]), .P13(n83[13]), .P12(n83[12]), .P11(n83[11]), 
            .P10(n83[10]), .P9(n83[9]), .P8(n83[8]), .P7(n83[7]), .P6(n83[6]), 
            .P5(n83[5]), .P4(n83[4]), .P3(n83[3]), .P2(n83[2]), .P1(n83[1]), 
            .P0(n83[0]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_mult_2.REG_INPUTA_CLK = "NONE";
    defparam MultResult2_res2_mult_2.REG_INPUTA_CE = "CE0";
    defparam MultResult2_res2_mult_2.REG_INPUTA_RST = "RST0";
    defparam MultResult2_res2_mult_2.REG_INPUTB_CLK = "NONE";
    defparam MultResult2_res2_mult_2.REG_INPUTB_CE = "CE0";
    defparam MultResult2_res2_mult_2.REG_INPUTB_RST = "RST0";
    defparam MultResult2_res2_mult_2.REG_INPUTC_CLK = "NONE";
    defparam MultResult2_res2_mult_2.REG_INPUTC_CE = "CE0";
    defparam MultResult2_res2_mult_2.REG_INPUTC_RST = "RST0";
    defparam MultResult2_res2_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam MultResult2_res2_mult_2.REG_PIPELINE_CE = "CE0";
    defparam MultResult2_res2_mult_2.REG_PIPELINE_RST = "RST0";
    defparam MultResult2_res2_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam MultResult2_res2_mult_2.REG_OUTPUT_CE = "CE0";
    defparam MultResult2_res2_mult_2.REG_OUTPUT_RST = "RST0";
    defparam MultResult2_res2_mult_2.CLK0_DIV = "ENABLED";
    defparam MultResult2_res2_mult_2.CLK1_DIV = "ENABLED";
    defparam MultResult2_res2_mult_2.CLK2_DIV = "ENABLED";
    defparam MultResult2_res2_mult_2.CLK3_DIV = "ENABLED";
    defparam MultResult2_res2_mult_2.HIGHSPEED_CLK = "NONE";
    defparam MultResult2_res2_mult_2.GSR = "ENABLED";
    defparam MultResult2_res2_mult_2.CAS_MATCH_REG = "FALSE";
    defparam MultResult2_res2_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam MultResult2_res2_mult_2.MULT_BYPASS = "DISABLED";
    defparam MultResult2_res2_mult_2.RESETMODE = "SYNC";
    FD1S3AX d_out_i2 (.D(d_out_d[1]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i2.GSR = "ENABLED";
    FD1S3AX d_out_i3 (.D(d_out_d[2]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i3.GSR = "ENABLED";
    FD1S3AX d_out_i4 (.D(d_out_d[3]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i4.GSR = "ENABLED";
    FD1S3AX d_out_i5 (.D(d_out_d[4]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i5.GSR = "ENABLED";
    FD1S3AX d_out_i6 (.D(d_out_d[5]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i6.GSR = "ENABLED";
    FD1S3AX d_out_i7 (.D(d_out_d[6]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i7.GSR = "ENABLED";
    FD1S3AX d_out_i8 (.D(d_out_d[7]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i8.GSR = "ENABLED";
    FD1S3AX d_out_i9 (.D(d_out_d[8]), .CK(CIC1_out_clkSin), .Q(\DataInReg_11__N_1856[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i9.GSR = "ENABLED";
    FD1S3AX d_out_i10 (.D(d_out_d[9]), .CK(CIC1_out_clkSin), .Q(\DemodOut[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_i10.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i2 (.D(CIC1_outCos[1]), .CK(CIC1_out_clkSin), 
            .Q(n27[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i2.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i3 (.D(CIC1_outCos[2]), .CK(CIC1_out_clkSin), 
            .Q(n27[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i3.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i4 (.D(CIC1_outCos[3]), .CK(CIC1_out_clkSin), 
            .Q(n27[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i4.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i5 (.D(CIC1_outCos[4]), .CK(CIC1_out_clkSin), 
            .Q(n27[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i5.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i6 (.D(CIC1_outCos[5]), .CK(CIC1_out_clkSin), 
            .Q(n27[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i6.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i7 (.D(CIC1_outCos[6]), .CK(CIC1_out_clkSin), 
            .Q(n27[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i7.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i8 (.D(CIC1_outCos[7]), .CK(CIC1_out_clkSin), 
            .Q(n27[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i8.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i9 (.D(CIC1_outCos[8]), .CK(CIC1_out_clkSin), 
            .Q(n27[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i9.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i10 (.D(CIC1_outCos[9]), .CK(CIC1_out_clkSin), 
            .Q(n27[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i10.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i11 (.D(CIC1_outCos[10]), .CK(CIC1_out_clkSin), 
            .Q(n27[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i11.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e1__i12 (.D(CIC1_outCos[11]), .CK(CIC1_out_clkSin), 
            .Q(n27[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e1__i12.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i1 (.D(n83[1]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i1.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i2 (.D(n83[2]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i2.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i3 (.D(n83[3]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i3.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i4 (.D(n83[4]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i4.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i5 (.D(n83[5]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i5.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i6 (.D(n83[6]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i6.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i7 (.D(n83[7]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i7.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i8 (.D(n83[8]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i8.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i9 (.D(n83[9]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i9.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i10 (.D(n83[10]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i10.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i11 (.D(n83[11]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i11.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i12 (.D(n83[12]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i12.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i13 (.D(n83[13]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i13.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i14 (.D(n83[14]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i14.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i15 (.D(n83[15]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i15.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i16 (.D(n83[16]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i16.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i17 (.D(n83[17]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i17.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i18 (.D(n83[18]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i18.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i19 (.D(n83[19]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i19.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i20 (.D(n83[20]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i20.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i21 (.D(n83[21]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i21.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i22 (.D(n83[22]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i22.GSR = "ENABLED";
    FD1S3AX MultResult2_res2_e3_i0_i23 (.D(n83[23]), .CK(CIC1_out_clkSin), 
            .Q(MultResult2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=18, LSE_RCOL=5, LSE_LLINE=171, LSE_RLINE=176 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(87[20:39])
    defparam MultResult2_res2_e3_i0_i23.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i2 (.D(d_out_d_11__N_1891), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[1]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i2.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i3 (.D(d_out_d_11__N_1889), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[2]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i3.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i4 (.D(d_out_d_11__N_1887), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[3]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i4.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i5 (.D(d_out_d_11__N_1885), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[4]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i5.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i6 (.D(d_out_d_11__N_1883), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[5]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i6.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i7 (.D(d_out_d_11__N_1881), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[6]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i7.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i8 (.D(d_out_d_11__N_1879), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[7]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i8.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i9 (.D(d_out_d_11__N_1877), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[8]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i9.GSR = "ENABLED";
    FD1S3AX d_out_d__0_i10 (.D(d_out_d_11__N_1875), .CK(CIC1_out_clkSin), 
            .Q(d_out_d[9]));   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(79[10] 97[6])
    defparam d_out_d__0_i10.GSR = "ENABLED";
    LUT4 mux_81_i1_3_lut (.A(\d_out_d_11__N_2383[17] ), .B(\d_out_d_11__N_2401[17] ), 
         .C(\d_out_d_11__N_1892[17] ), .Z(d_out_d_11__N_1894[17])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(70[11:28])
    defparam mux_81_i1_3_lut.init = 16'h3535;
    LUT4 i1344_1_lut (.A(\ISquare[31] ), .Z(n213)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1344_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_1_1_lut (.A(\d_out_d_11__N_1874[17] ), .Z(d_out_d_11__N_1873)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_1_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_8_1_lut (.A(\d_out_d_11__N_1888[17] ), .Z(d_out_d_11__N_1887)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_8_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_10_1_lut (.A(\d_out_d_11__N_1892[17] ), .Z(d_out_d_11__N_1891)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_10_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_9_1_lut (.A(\d_out_d_11__N_1890[17] ), .Z(d_out_d_11__N_1889)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_9_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_7_1_lut (.A(\d_out_d_11__N_1886[17] ), .Z(d_out_d_11__N_1885)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_7_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_6_1_lut (.A(\d_out_d_11__N_1884[17] ), .Z(d_out_d_11__N_1883)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_6_1_lut.init = 16'h5555;
    LUT4 d_out_d_11__I_5_1_lut (.A(\d_out_d_11__N_1882[17] ), .Z(d_out_d_11__N_1881)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/AMDemod.v(71[23:29])
    defparam d_out_d_11__I_5_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module \CIC(WIDTH=72,DECIMATION_RATIO=4096)_U0 
//

module \CIC(WIDTH=72,DECIMATION_RATIO=4096)_U0  (d_tmp, clk_80mhz, d5, 
            d_d_tmp, d2, d2_71__N_490, d_d8, n11, d3, d3_71__N_562, 
            d4, d4_71__N_634, d5_71__N_706, d6, d6_71__N_1459, d_d6, 
            CIC1_out_clkSin, d7, d7_71__N_1531, d_d7, d8, d8_71__N_1603, 
            d9, d9_71__N_1675, d_d9, n26, MultDataB, d1, d1_71__N_418, 
            count, n29, n10, n13, n12, n15, \CICGain[1] , n18, 
            n21, n20, n23, n22, n25, n24, n27, n26_adj_1, n29_adj_2, 
            n28, n31, n30, n33, n118, n120, cout, n115, n117, 
            n112, n114, n32, n35, n109, n111, n34, n106, n108, 
            n37, n103, n105, n36, n3, n2, n100, n102, n97, 
            n99, n5, n4, n94, n96, n91, n93, n88, n90, n7, 
            n85, n87, n82, n84, n79, n81, n76, n78, n14, n6, 
            n8, \d10[68] , \d10[66] , \d10[67] , n28_adj_3, n31_adj_4, 
            n11_adj_5, n9, \d10[65] , \d_out_11__N_1819[2] , \d_out_11__N_1819[3] , 
            \d_out_11__N_1819[4] , \d_out_11__N_1819[5] , \d_out_11__N_1819[6] , 
            \d_out_11__N_1819[7] , \d_out_11__N_1819[8] , n87_adj_126, 
            \CICGain[0] , n30_adj_9, n63_adj_10, n65, n135, n64, 
            n134, n133, n8_adj_11, n132, n66_adj_12, n136, n11_adj_13, 
            n10_adj_14, n66_adj_15, \d10[64] , n136_adj_16, n65_adj_17, 
            \d10[63] , n135_adj_18, n63_adj_19, \d10[61] , n133_adj_20, 
            n13_adj_21, \d10[68]_adj_22 , \d10[69] , \d10[71] , \d10[70] , 
            n64_adj_23, \d10[62] , n134_adj_24, n17, n16, n19, n18_adj_25, 
            n21_adj_26, n20_adj_27, n23_adj_28, n22_adj_29, n17610, 
            \d10[60] , n132_adj_30, n17630, \d10[59] , n131, n12_adj_31, 
            n3_adj_32, n2_adj_33, n10_adj_34, n13_adj_35, n12_adj_36, 
            n15_adj_37, n14_adj_38, n17_adj_39, n16_adj_40, n19_adj_41, 
            n131_adj_42, \d10[67]_adj_43 , n18_adj_44, n21_adj_45, n20_adj_46, 
            n23_adj_47, n22_adj_48, n25_adj_49, n24_adj_50, n25_adj_51, 
            n24_adj_52, n27_adj_53, n26_adj_54, n29_adj_55, n28_adj_56, 
            n31_adj_57, n30_adj_58, n33_adj_59, n32_adj_60, n27_adj_61, 
            n35_adj_62, n34_adj_63, n37_adj_64, n36_adj_65, n15_adj_66, 
            n14_adj_67, n17_adj_68, n16_adj_69, n5_adj_70, n4_adj_71, 
            n33_adj_72, n7_adj_73, n32_adj_74, n35_adj_75, n34_adj_76, 
            n6_adj_77, n9_adj_78, n8_adj_79, n11_adj_80, n37_adj_81, 
            n10_adj_82, n36_adj_83, n13_adj_84, n3_adj_85, n2_adj_86, 
            n5_adj_87, n12_adj_88, n4_adj_89, n7_adj_90, n15_adj_91, 
            n14_adj_92, n6_adj_93, n17_adj_94, n19_adj_95, n18_adj_96, 
            n9_adj_97, n16_adj_98, \d_out_11__N_1819[10] , n19_adj_99, 
            n21_adj_100, n20_adj_101, \d_out_11__N_1819[11] , n23_adj_102, 
            n22_adj_103, n25_adj_104, n24_adj_105, n27_adj_106, n26_adj_107, 
            n29_adj_108, n28_adj_109, n31_adj_110, n30_adj_111, n33_adj_112, 
            n32_adj_113, n35_adj_114, n34_adj_115, n37_adj_116, n36_adj_117, 
            n3_adj_118, n2_adj_119, n5_adj_120, n4_adj_121, n7_adj_122, 
            n6_adj_123, n9_adj_124, n8_adj_125) /* synthesis syn_module_defined=1 */ ;
    output [71:0]d_tmp;
    input clk_80mhz;
    output [71:0]d5;
    output [71:0]d_d_tmp;
    output [71:0]d2;
    input [71:0]d2_71__N_490;
    output [71:0]d_d8;
    output n11;
    output [71:0]d3;
    input [71:0]d3_71__N_562;
    output [71:0]d4;
    input [71:0]d4_71__N_634;
    input [71:0]d5_71__N_706;
    output [71:0]d6;
    input [71:0]d6_71__N_1459;
    output [71:0]d_d6;
    output CIC1_out_clkSin;
    output [71:0]d7;
    input [71:0]d7_71__N_1531;
    output [71:0]d_d7;
    output [71:0]d8;
    input [71:0]d8_71__N_1603;
    output [71:0]d9;
    input [71:0]d9_71__N_1675;
    output [71:0]d_d9;
    output n26;
    output [11:0]MultDataB;
    output [71:0]d1;
    input [71:0]d1_71__N_418;
    output [15:0]count;
    output n29;
    output n10;
    output n13;
    output n12;
    output n15;
    input \CICGain[1] ;
    output n18;
    output n21;
    output n20;
    output n23;
    output n22;
    output n25;
    output n24;
    output n27;
    output n26_adj_1;
    output n29_adj_2;
    output n28;
    output n31;
    output n30;
    output n33;
    input n118;
    input n120;
    input cout;
    input n115;
    input n117;
    input n112;
    input n114;
    output n32;
    output n35;
    input n109;
    input n111;
    output n34;
    input n106;
    input n108;
    output n37;
    input n103;
    input n105;
    output n36;
    output n3;
    output n2;
    input n100;
    input n102;
    input n97;
    input n99;
    output n5;
    output n4;
    input n94;
    input n96;
    input n91;
    input n93;
    input n88;
    input n90;
    output n7;
    input n85;
    input n87;
    input n82;
    input n84;
    input n79;
    input n81;
    input n76;
    input n78;
    output n14;
    output n6;
    output n8;
    output \d10[68] ;
    output \d10[66] ;
    output \d10[67] ;
    output n28_adj_3;
    output n31_adj_4;
    output n11_adj_5;
    output n9;
    output \d10[65] ;
    input \d_out_11__N_1819[2] ;
    input \d_out_11__N_1819[3] ;
    input \d_out_11__N_1819[4] ;
    input \d_out_11__N_1819[5] ;
    input \d_out_11__N_1819[6] ;
    input \d_out_11__N_1819[7] ;
    input \d_out_11__N_1819[8] ;
    input [15:0]n87_adj_126;
    input \CICGain[0] ;
    output n30_adj_9;
    output n63_adj_10;
    output n65;
    output n135;
    output n64;
    output n134;
    output n133;
    output n8_adj_11;
    output n132;
    output n66_adj_12;
    output n136;
    output n11_adj_13;
    output n10_adj_14;
    input n66_adj_15;
    input \d10[64] ;
    output n136_adj_16;
    input n65_adj_17;
    input \d10[63] ;
    output n135_adj_18;
    input n63_adj_19;
    input \d10[61] ;
    output n133_adj_20;
    output n13_adj_21;
    input \d10[68]_adj_22 ;
    input \d10[69] ;
    input \d10[71] ;
    input \d10[70] ;
    input n64_adj_23;
    input \d10[62] ;
    output n134_adj_24;
    output n17;
    output n16;
    output n19;
    output n18_adj_25;
    output n21_adj_26;
    output n20_adj_27;
    output n23_adj_28;
    output n22_adj_29;
    input n17610;
    input \d10[60] ;
    output n132_adj_30;
    input n17630;
    input \d10[59] ;
    output n131;
    output n12_adj_31;
    output n3_adj_32;
    output n2_adj_33;
    output n10_adj_34;
    output n13_adj_35;
    output n12_adj_36;
    output n15_adj_37;
    output n14_adj_38;
    output n17_adj_39;
    output n16_adj_40;
    output n19_adj_41;
    output n131_adj_42;
    input \d10[67]_adj_43 ;
    output n18_adj_44;
    output n21_adj_45;
    output n20_adj_46;
    output n23_adj_47;
    output n22_adj_48;
    output n25_adj_49;
    output n24_adj_50;
    output n25_adj_51;
    output n24_adj_52;
    output n27_adj_53;
    output n26_adj_54;
    output n29_adj_55;
    output n28_adj_56;
    output n31_adj_57;
    output n30_adj_58;
    output n33_adj_59;
    output n32_adj_60;
    output n27_adj_61;
    output n35_adj_62;
    output n34_adj_63;
    output n37_adj_64;
    output n36_adj_65;
    output n15_adj_66;
    output n14_adj_67;
    output n17_adj_68;
    output n16_adj_69;
    output n5_adj_70;
    output n4_adj_71;
    output n33_adj_72;
    output n7_adj_73;
    output n32_adj_74;
    output n35_adj_75;
    output n34_adj_76;
    output n6_adj_77;
    output n9_adj_78;
    output n8_adj_79;
    output n11_adj_80;
    output n37_adj_81;
    output n10_adj_82;
    output n36_adj_83;
    output n13_adj_84;
    output n3_adj_85;
    output n2_adj_86;
    output n5_adj_87;
    output n12_adj_88;
    output n4_adj_89;
    output n7_adj_90;
    output n15_adj_91;
    output n14_adj_92;
    output n6_adj_93;
    output n17_adj_94;
    output n19_adj_95;
    output n18_adj_96;
    output n9_adj_97;
    output n16_adj_98;
    output \d_out_11__N_1819[10] ;
    output n19_adj_99;
    output n21_adj_100;
    output n20_adj_101;
    output \d_out_11__N_1819[11] ;
    output n23_adj_102;
    output n22_adj_103;
    output n25_adj_104;
    output n24_adj_105;
    output n27_adj_106;
    output n26_adj_107;
    output n29_adj_108;
    output n28_adj_109;
    output n31_adj_110;
    output n30_adj_111;
    output n33_adj_112;
    output n32_adj_113;
    output n35_adj_114;
    output n34_adj_115;
    output n37_adj_116;
    output n36_adj_117;
    output n3_adj_118;
    output n2_adj_119;
    output n5_adj_120;
    output n4_adj_121;
    output n7_adj_122;
    output n6_adj_123;
    output n9_adj_124;
    output n8_adj_125;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(61[23:32])
    wire CIC1_out_clkSin /* synthesis SET_AS_NETWORK=CIC1_out_clkSin, is_clock=1 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/top.v(74[23:38])
    
    wire clk_80mhz_enable_129, clk_80mhz_enable_65, d_clk_tmp, n12681, 
        v_comb, clk_80mhz_enable_11;
    wire [71:0]d_out_11__N_1819;
    wire [15:0]count_15__N_1442;
    
    wire n17459, n17054, n17463, n17461, n31_c;
    wire [71:0]d10;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(54[68:71])
    
    wire n17957, n17655, n17956, n17963, n17636, n17962, n17586, 
        n17562, n17554, d_clk_tmp_N_1831, n17580;
    wire [71:0]d10_71__N_1747;
    
    wire clk_80mhz_enable_706, n17469, n18089, n17972, n17628, n17971, 
        clk_80mhz_enable_149, clk_80mhz_enable_199, clk_80mhz_enable_249, 
        clk_80mhz_enable_299, clk_80mhz_enable_349, clk_80mhz_enable_399, 
        clk_80mhz_enable_449, clk_80mhz_enable_499, clk_80mhz_enable_549, 
        clk_80mhz_enable_599, clk_80mhz_enable_649, clk_80mhz_enable_699, 
        clk_80mhz_enable_700, clk_80mhz_enable_701, clk_80mhz_enable_702, 
        clk_80mhz_enable_703, clk_80mhz_enable_704, clk_80mhz_enable_705, 
        clk_80mhz_enable_707, clk_80mhz_enable_708, clk_80mhz_enable_709, 
        clk_80mhz_enable_710, n12697, n17984, n17983, n17987, n17986, 
        n17990, n17989, n17993, n17992;
    
    FD1P3AX d_tmp_i0_i0 (.D(d5[0]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i0 (.D(d_tmp[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i0.GSR = "ENABLED";
    FD1S3AX d2_i0 (.D(d2_71__N_490[0]), .CK(clk_80mhz), .Q(d2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i0.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i63_1_lut (.A(d_d8[62]), .Z(n11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i63_1_lut.init = 16'h5555;
    FD1S3AX d3_i0 (.D(d3_71__N_562[0]), .CK(clk_80mhz), .Q(d3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i0.GSR = "ENABLED";
    FD1S3AX d4_i0 (.D(d4_71__N_634[0]), .CK(clk_80mhz), .Q(d4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i0.GSR = "ENABLED";
    FD1S3AX d5_i0 (.D(d5_71__N_706[0]), .CK(clk_80mhz), .Q(d5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i0.GSR = "ENABLED";
    FD1P3AX d6_i0_i0 (.D(d6_71__N_1459[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i0 (.D(d6[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i0.GSR = "ENABLED";
    FD1S3JX d_clk_tmp_65 (.D(n12681), .CK(clk_80mhz), .PD(clk_80mhz_enable_129), 
            .Q(d_clk_tmp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_clk_tmp_65.GSR = "ENABLED";
    FD1S3AX v_comb_66 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), .Q(v_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66.GSR = "ENABLED";
    FD1S3AX d_clk_67 (.D(d_clk_tmp), .CK(clk_80mhz), .Q(CIC1_out_clkSin)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_clk_67.GSR = "ENABLED";
    FD1P3AX d7_i0_i0 (.D(d7_71__N_1531[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i0 (.D(d7[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX d8_i0_i0 (.D(d8_71__N_1603[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i0 (.D(d8[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX d9_i0_i0 (.D(d9_71__N_1675[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i0.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i0 (.D(d9[0]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i0.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i48_1_lut (.A(d_d8[47]), .Z(n26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i48_1_lut.init = 16'h5555;
    FD1P3AX d_out_i0_i0 (.D(d_out_11__N_1819[0]), .SP(clk_80mhz_enable_11), 
            .CK(clk_80mhz), .Q(MultDataB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i0.GSR = "ENABLED";
    FD1S3AX d1_i0 (.D(d1_71__N_418[0]), .CK(clk_80mhz), .Q(d1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i0.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_15__N_1442[0]), .CK(clk_80mhz), .CD(clk_80mhz_enable_129), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i0.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i45_1_lut (.A(d_d8[44]), .Z(n29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i64_1_lut (.A(d_d8[63]), .Z(n10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 i1_4_lut (.A(n17459), .B(n17054), .C(n17463), .D(n17461), .Z(n31_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 sub_28_inv_0_i61_1_lut (.A(d_d8[60]), .Z(n13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i62_1_lut (.A(d_d8[61]), .Z(n12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i59_1_lut (.A(d_d8[58]), .Z(n15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 i6381_then_3_lut (.A(\CICGain[1] ), .B(d10[59]), .C(d10[57]), 
         .Z(n17957)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6381_then_3_lut.init = 16'he4e4;
    LUT4 sub_26_inv_0_i56_1_lut (.A(d_d6[55]), .Z(n18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 i6381_else_3_lut (.A(n17655), .B(\CICGain[1] ), .C(d10[58]), 
         .Z(n17956)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6381_else_3_lut.init = 16'he2e2;
    LUT4 sub_26_inv_0_i53_1_lut (.A(d_d6[52]), .Z(n21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i54_1_lut (.A(d_d6[53]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 i6404_then_3_lut (.A(\CICGain[1] ), .B(d10[60]), .C(d10[58]), 
         .Z(n17963)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6404_then_3_lut.init = 16'he4e4;
    LUT4 i6404_else_3_lut (.A(n17636), .B(\CICGain[1] ), .C(d10[59]), 
         .Z(n17962)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6404_else_3_lut.init = 16'he2e2;
    LUT4 sub_26_inv_0_i51_1_lut (.A(d_d6[50]), .Z(n23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i52_1_lut (.A(d_d6[51]), .Z(n22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i49_1_lut (.A(d_d6[48]), .Z(n25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i50_1_lut (.A(d_d6[49]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i47_1_lut (.A(d_d6[46]), .Z(n27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i48_1_lut (.A(d_d6[47]), .Z(n26_adj_1)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i45_1_lut (.A(d_d6[44]), .Z(n29_adj_2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 i6329_4_lut (.A(n17054), .B(n17586), .C(n17562), .D(n17554), 
         .Z(d_clk_tmp_N_1831)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i6329_4_lut.init = 16'h4000;
    LUT4 sub_26_inv_0_i46_1_lut (.A(d_d6[45]), .Z(n28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i43_1_lut (.A(d_d6[42]), .Z(n31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i44_1_lut (.A(d_d6[43]), .Z(n30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 i6292_4_lut (.A(count[7]), .B(n17580), .C(count[0]), .D(count[10]), 
         .Z(n17586)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6292_4_lut.init = 16'h8000;
    LUT4 sub_26_inv_0_i41_1_lut (.A(d_d6[40]), .Z(n33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 mux_1250_i2_3_lut (.A(n118), .B(n120), .C(cout), .Z(d10_71__N_1747[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i3_3_lut (.A(n115), .B(n117), .C(cout), .Z(d10_71__N_1747[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i4_3_lut (.A(n112), .B(n114), .C(cout), .Z(d10_71__N_1747[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i4_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i42_1_lut (.A(d_d6[41]), .Z(n32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i39_1_lut (.A(d_d6[38]), .Z(n35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 mux_1250_i5_3_lut (.A(n109), .B(n111), .C(cout), .Z(d10_71__N_1747[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i5_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i40_1_lut (.A(d_d6[39]), .Z(n34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 mux_1250_i6_3_lut (.A(n106), .B(n108), .C(cout), .Z(d10_71__N_1747[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i6_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i37_1_lut (.A(d_d6[36]), .Z(n37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 i6268_2_lut (.A(count[6]), .B(count[4]), .Z(n17562)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6268_2_lut.init = 16'h8888;
    LUT4 mux_1250_i7_3_lut (.A(n103), .B(n105), .C(cout), .Z(d10_71__N_1747[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i7_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i38_1_lut (.A(d_d6[37]), .Z(n36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i71_1_lut (.A(d_d_tmp[70]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i72_1_lut (.A(d_d_tmp[71]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 mux_1250_i8_3_lut (.A(n100), .B(n102), .C(cout), .Z(d10_71__N_1747[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i8_3_lut.init = 16'hcaca;
    LUT4 i6260_2_lut (.A(count[1]), .B(count[3]), .Z(n17554)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6260_2_lut.init = 16'h8888;
    LUT4 i6286_4_lut (.A(count[5]), .B(count[2]), .C(count[9]), .D(count[8]), 
         .Z(n17580)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6286_4_lut.init = 16'h8000;
    LUT4 mux_1250_i9_3_lut (.A(n97), .B(n99), .C(cout), .Z(d10_71__N_1747[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i9_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i69_1_lut (.A(d_d_tmp[68]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i69_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_189 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_706)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_189.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i70_1_lut (.A(d_d_tmp[69]), .Z(n4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_25 (.A(count[12]), .B(count[11]), .C(n17469), .D(count[15]), 
         .Z(n17054)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_25.init = 16'hfffb;
    LUT4 mux_1250_i10_3_lut (.A(n94), .B(n96), .C(cout), .Z(d10_71__N_1747[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i11_3_lut (.A(n91), .B(n93), .C(cout), .Z(d10_71__N_1747[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i12_3_lut (.A(n88), .B(n90), .C(cout), .Z(d10_71__N_1747[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i12_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i67_1_lut (.A(d_d_tmp[66]), .Z(n7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 i1_2_lut (.A(count[14]), .B(count[13]), .Z(n17469)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 mux_1250_i13_3_lut (.A(n85), .B(n87), .C(cout), .Z(d10_71__N_1747[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i14_3_lut (.A(n82), .B(n84), .C(cout), .Z(d10_71__N_1747[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i15_3_lut (.A(n79), .B(n81), .C(cout), .Z(d10_71__N_1747[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1250_i16_3_lut (.A(n76), .B(n78), .C(cout), .Z(d10_71__N_1747[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(99[25:34])
    defparam mux_1250_i16_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i60_1_lut (.A(d_d8[59]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 i6329_4_lut_rep_194 (.A(n17054), .B(n17586), .C(n17562), .D(n17554), 
         .Z(n18089)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i6329_4_lut_rep_194.init = 16'h4000;
    LUT4 sub_25_inv_0_i68_1_lut (.A(d_d_tmp[67]), .Z(n6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i66_1_lut (.A(d_d7[65]), .Z(n8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 i6397_then_3_lut (.A(\CICGain[1] ), .B(\d10[68] ), .C(\d10[66] ), 
         .Z(n17972)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i6397_then_3_lut.init = 16'he4e4;
    LUT4 i6397_else_3_lut (.A(n17628), .B(\CICGain[1] ), .C(\d10[67] ), 
         .Z(n17971)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i6397_else_3_lut.init = 16'he2e2;
    FD1P3AX d_d_tmp_i0_i71 (.D(d_tmp[71]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i70 (.D(d_tmp[70]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i69 (.D(d_tmp[69]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i68 (.D(d_tmp[68]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i67 (.D(d_tmp[67]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i66 (.D(d_tmp[66]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i65 (.D(d_tmp[65]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i64 (.D(d_tmp[64]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i63 (.D(d_tmp[63]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i62 (.D(d_tmp[62]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i61 (.D(d_tmp[61]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i60 (.D(d_tmp[60]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i59 (.D(d_tmp[59]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i58 (.D(d_tmp[58]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i57 (.D(d_tmp[57]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i56 (.D(d_tmp[56]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i55 (.D(d_tmp[55]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i54 (.D(d_tmp[54]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i53 (.D(d_tmp[53]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i52 (.D(d_tmp[52]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i51 (.D(d_tmp[51]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i50 (.D(d_tmp[50]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i49 (.D(d_tmp[49]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i48 (.D(d_tmp[48]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i47 (.D(d_tmp[47]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i46 (.D(d_tmp[46]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i45 (.D(d_tmp[45]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i44 (.D(d_tmp[44]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i43 (.D(d_tmp[43]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i42 (.D(d_tmp[42]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i41 (.D(d_tmp[41]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i40 (.D(d_tmp[40]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i39 (.D(d_tmp[39]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i38 (.D(d_tmp[38]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i37 (.D(d_tmp[37]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i36 (.D(d_tmp[36]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i35 (.D(d_tmp[35]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i34 (.D(d_tmp[34]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i33 (.D(d_tmp[33]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i32 (.D(d_tmp[32]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i31 (.D(d_tmp[31]), .SP(clk_80mhz_enable_65), .CK(clk_80mhz), 
            .Q(d_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i30 (.D(d_tmp[30]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i29 (.D(d_tmp[29]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i28 (.D(d_tmp[28]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i27 (.D(d_tmp[27]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i26 (.D(d_tmp[26]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i25 (.D(d_tmp[25]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i24 (.D(d_tmp[24]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i23 (.D(d_tmp[23]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i22 (.D(d_tmp[22]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i21 (.D(d_tmp[21]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i20 (.D(d_tmp[20]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i19 (.D(d_tmp[19]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i18 (.D(d_tmp[18]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i17 (.D(d_tmp[17]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i16 (.D(d_tmp[16]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i15 (.D(d_tmp[15]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i14 (.D(d_tmp[14]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i13 (.D(d_tmp[13]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i12 (.D(d_tmp[12]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i11 (.D(d_tmp[11]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i10 (.D(d_tmp[10]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i9 (.D(d_tmp[9]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i8 (.D(d_tmp[8]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i7 (.D(d_tmp[7]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i6 (.D(d_tmp[6]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i5 (.D(d_tmp[5]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i4 (.D(d_tmp[4]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i3 (.D(d_tmp[3]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i2 (.D(d_tmp[2]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d_tmp_i0_i1 (.D(d_tmp[1]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i71 (.D(d5[71]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i70 (.D(d5[70]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i69 (.D(d5[69]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i68 (.D(d5[68]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i67 (.D(d5[67]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i66 (.D(d5[66]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i65 (.D(d5[65]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i64 (.D(d5[64]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i63 (.D(d5[63]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i62 (.D(d5[62]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i61 (.D(d5[61]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i60 (.D(d5[60]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i59 (.D(d5[59]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i58 (.D(d5[58]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i57 (.D(d5[57]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i56 (.D(d5[56]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i55 (.D(d5[55]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i54 (.D(d5[54]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i53 (.D(d5[53]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i52 (.D(d5[52]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i51 (.D(d5[51]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i50 (.D(d5[50]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i49 (.D(d5[49]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i48 (.D(d5[48]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i47 (.D(d5[47]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i46 (.D(d5[46]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i45 (.D(d5[45]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i44 (.D(d5[44]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i43 (.D(d5[43]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i42 (.D(d5[42]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i41 (.D(d5[41]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i40 (.D(d5[40]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i39 (.D(d5[39]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i38 (.D(d5[38]), .SP(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i37 (.D(d5[37]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i36 (.D(d5[36]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i35 (.D(d5[35]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i34 (.D(d5[34]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i33 (.D(d5[33]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i32 (.D(d5[32]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i31 (.D(d5[31]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i30 (.D(d5[30]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i29 (.D(d5[29]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i28 (.D(d5[28]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i27 (.D(d5[27]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i26 (.D(d5[26]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i25 (.D(d5[25]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i24 (.D(d5[24]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i23 (.D(d5[23]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i22 (.D(d5[22]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i21 (.D(d5[21]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i20 (.D(d5[20]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i19 (.D(d5[19]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i18 (.D(d5[18]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i17 (.D(d5[17]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i16 (.D(d5[16]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i15 (.D(d5[15]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i14 (.D(d5[14]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i13 (.D(d5[13]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i12 (.D(d5[12]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i11 (.D(d5[11]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i10 (.D(d5[10]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i9 (.D(d5[9]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i8 (.D(d5[8]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i7 (.D(d5[7]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i6 (.D(d5[6]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i5 (.D(d5[5]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i4 (.D(d5[4]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i3 (.D(d5[3]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i2 (.D(d5[2]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX d_tmp_i0_i1 (.D(d5[1]), .SP(d_clk_tmp_N_1831), .CK(clk_80mhz), 
            .Q(d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d_tmp_i0_i1.GSR = "ENABLED";
    FD1S3AX d2_i1 (.D(d2_71__N_490[1]), .CK(clk_80mhz), .Q(d2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i1.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i46_1_lut (.A(d_d8[45]), .Z(n28_adj_3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i43_1_lut (.A(d_d8[42]), .Z(n31_adj_4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i63_1_lut (.A(d_d7[62]), .Z(n11_adj_5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i65_1_lut (.A(d_d_tmp[64]), .Z(n9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i65_1_lut.init = 16'h5555;
    FD1S3AX d2_i2 (.D(d2_71__N_490[2]), .CK(clk_80mhz), .Q(d2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i2.GSR = "ENABLED";
    FD1S3AX d2_i3 (.D(d2_71__N_490[3]), .CK(clk_80mhz), .Q(d2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i3.GSR = "ENABLED";
    FD1S3AX d2_i4 (.D(d2_71__N_490[4]), .CK(clk_80mhz), .Q(d2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i4.GSR = "ENABLED";
    FD1S3AX d2_i5 (.D(d2_71__N_490[5]), .CK(clk_80mhz), .Q(d2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i5.GSR = "ENABLED";
    FD1S3AX d2_i6 (.D(d2_71__N_490[6]), .CK(clk_80mhz), .Q(d2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i6.GSR = "ENABLED";
    FD1S3AX d2_i7 (.D(d2_71__N_490[7]), .CK(clk_80mhz), .Q(d2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i7.GSR = "ENABLED";
    FD1S3AX d2_i8 (.D(d2_71__N_490[8]), .CK(clk_80mhz), .Q(d2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i8.GSR = "ENABLED";
    FD1S3AX d2_i9 (.D(d2_71__N_490[9]), .CK(clk_80mhz), .Q(d2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i9.GSR = "ENABLED";
    FD1S3AX d2_i10 (.D(d2_71__N_490[10]), .CK(clk_80mhz), .Q(d2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i10.GSR = "ENABLED";
    FD1S3AX d2_i11 (.D(d2_71__N_490[11]), .CK(clk_80mhz), .Q(d2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i11.GSR = "ENABLED";
    FD1S3AX d2_i12 (.D(d2_71__N_490[12]), .CK(clk_80mhz), .Q(d2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i12.GSR = "ENABLED";
    FD1S3AX d2_i13 (.D(d2_71__N_490[13]), .CK(clk_80mhz), .Q(d2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i13.GSR = "ENABLED";
    FD1S3AX d2_i14 (.D(d2_71__N_490[14]), .CK(clk_80mhz), .Q(d2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i14.GSR = "ENABLED";
    FD1S3AX d2_i15 (.D(d2_71__N_490[15]), .CK(clk_80mhz), .Q(d2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i15.GSR = "ENABLED";
    FD1S3AX d2_i16 (.D(d2_71__N_490[16]), .CK(clk_80mhz), .Q(d2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i16.GSR = "ENABLED";
    FD1S3AX d2_i17 (.D(d2_71__N_490[17]), .CK(clk_80mhz), .Q(d2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i17.GSR = "ENABLED";
    FD1S3AX d2_i18 (.D(d2_71__N_490[18]), .CK(clk_80mhz), .Q(d2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i18.GSR = "ENABLED";
    FD1S3AX d2_i19 (.D(d2_71__N_490[19]), .CK(clk_80mhz), .Q(d2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i19.GSR = "ENABLED";
    FD1S3AX d2_i20 (.D(d2_71__N_490[20]), .CK(clk_80mhz), .Q(d2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i20.GSR = "ENABLED";
    FD1S3AX d2_i21 (.D(d2_71__N_490[21]), .CK(clk_80mhz), .Q(d2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i21.GSR = "ENABLED";
    FD1S3AX d2_i22 (.D(d2_71__N_490[22]), .CK(clk_80mhz), .Q(d2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i22.GSR = "ENABLED";
    FD1S3AX d2_i23 (.D(d2_71__N_490[23]), .CK(clk_80mhz), .Q(d2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i23.GSR = "ENABLED";
    FD1S3AX d2_i24 (.D(d2_71__N_490[24]), .CK(clk_80mhz), .Q(d2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i24.GSR = "ENABLED";
    FD1S3AX d2_i25 (.D(d2_71__N_490[25]), .CK(clk_80mhz), .Q(d2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i25.GSR = "ENABLED";
    FD1S3AX d2_i26 (.D(d2_71__N_490[26]), .CK(clk_80mhz), .Q(d2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i26.GSR = "ENABLED";
    FD1S3AX d2_i27 (.D(d2_71__N_490[27]), .CK(clk_80mhz), .Q(d2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i27.GSR = "ENABLED";
    FD1S3AX d2_i28 (.D(d2_71__N_490[28]), .CK(clk_80mhz), .Q(d2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i28.GSR = "ENABLED";
    FD1S3AX d2_i29 (.D(d2_71__N_490[29]), .CK(clk_80mhz), .Q(d2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i29.GSR = "ENABLED";
    FD1S3AX d2_i30 (.D(d2_71__N_490[30]), .CK(clk_80mhz), .Q(d2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i30.GSR = "ENABLED";
    FD1S3AX d2_i31 (.D(d2_71__N_490[31]), .CK(clk_80mhz), .Q(d2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i31.GSR = "ENABLED";
    FD1S3AX d2_i32 (.D(d2_71__N_490[32]), .CK(clk_80mhz), .Q(d2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i32.GSR = "ENABLED";
    FD1S3AX d2_i33 (.D(d2_71__N_490[33]), .CK(clk_80mhz), .Q(d2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i33.GSR = "ENABLED";
    FD1S3AX d2_i34 (.D(d2_71__N_490[34]), .CK(clk_80mhz), .Q(d2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i34.GSR = "ENABLED";
    FD1S3AX d2_i35 (.D(d2_71__N_490[35]), .CK(clk_80mhz), .Q(d2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i35.GSR = "ENABLED";
    FD1S3AX d2_i36 (.D(d2_71__N_490[36]), .CK(clk_80mhz), .Q(d2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i36.GSR = "ENABLED";
    FD1S3AX d2_i37 (.D(d2_71__N_490[37]), .CK(clk_80mhz), .Q(d2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i37.GSR = "ENABLED";
    FD1S3AX d2_i38 (.D(d2_71__N_490[38]), .CK(clk_80mhz), .Q(d2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i38.GSR = "ENABLED";
    FD1S3AX d2_i39 (.D(d2_71__N_490[39]), .CK(clk_80mhz), .Q(d2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i39.GSR = "ENABLED";
    FD1S3AX d2_i40 (.D(d2_71__N_490[40]), .CK(clk_80mhz), .Q(d2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i40.GSR = "ENABLED";
    FD1S3AX d2_i41 (.D(d2_71__N_490[41]), .CK(clk_80mhz), .Q(d2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i41.GSR = "ENABLED";
    FD1S3AX d2_i42 (.D(d2_71__N_490[42]), .CK(clk_80mhz), .Q(d2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i42.GSR = "ENABLED";
    FD1S3AX d2_i43 (.D(d2_71__N_490[43]), .CK(clk_80mhz), .Q(d2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i43.GSR = "ENABLED";
    FD1S3AX d2_i44 (.D(d2_71__N_490[44]), .CK(clk_80mhz), .Q(d2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i44.GSR = "ENABLED";
    FD1S3AX d2_i45 (.D(d2_71__N_490[45]), .CK(clk_80mhz), .Q(d2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i45.GSR = "ENABLED";
    FD1S3AX d2_i46 (.D(d2_71__N_490[46]), .CK(clk_80mhz), .Q(d2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i46.GSR = "ENABLED";
    FD1S3AX d2_i47 (.D(d2_71__N_490[47]), .CK(clk_80mhz), .Q(d2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i47.GSR = "ENABLED";
    FD1S3AX d2_i48 (.D(d2_71__N_490[48]), .CK(clk_80mhz), .Q(d2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i48.GSR = "ENABLED";
    FD1S3AX d2_i49 (.D(d2_71__N_490[49]), .CK(clk_80mhz), .Q(d2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i49.GSR = "ENABLED";
    FD1S3AX d2_i50 (.D(d2_71__N_490[50]), .CK(clk_80mhz), .Q(d2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i50.GSR = "ENABLED";
    FD1S3AX d2_i51 (.D(d2_71__N_490[51]), .CK(clk_80mhz), .Q(d2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i51.GSR = "ENABLED";
    FD1S3AX d2_i52 (.D(d2_71__N_490[52]), .CK(clk_80mhz), .Q(d2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i52.GSR = "ENABLED";
    FD1S3AX d2_i53 (.D(d2_71__N_490[53]), .CK(clk_80mhz), .Q(d2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i53.GSR = "ENABLED";
    FD1S3AX d2_i54 (.D(d2_71__N_490[54]), .CK(clk_80mhz), .Q(d2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i54.GSR = "ENABLED";
    FD1S3AX d2_i55 (.D(d2_71__N_490[55]), .CK(clk_80mhz), .Q(d2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i55.GSR = "ENABLED";
    FD1S3AX d2_i56 (.D(d2_71__N_490[56]), .CK(clk_80mhz), .Q(d2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i56.GSR = "ENABLED";
    FD1S3AX d2_i57 (.D(d2_71__N_490[57]), .CK(clk_80mhz), .Q(d2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i57.GSR = "ENABLED";
    FD1S3AX d2_i58 (.D(d2_71__N_490[58]), .CK(clk_80mhz), .Q(d2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i58.GSR = "ENABLED";
    FD1S3AX d2_i59 (.D(d2_71__N_490[59]), .CK(clk_80mhz), .Q(d2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i59.GSR = "ENABLED";
    FD1S3AX d2_i60 (.D(d2_71__N_490[60]), .CK(clk_80mhz), .Q(d2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i60.GSR = "ENABLED";
    FD1S3AX d2_i61 (.D(d2_71__N_490[61]), .CK(clk_80mhz), .Q(d2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i61.GSR = "ENABLED";
    FD1S3AX d2_i62 (.D(d2_71__N_490[62]), .CK(clk_80mhz), .Q(d2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i62.GSR = "ENABLED";
    FD1S3AX d2_i63 (.D(d2_71__N_490[63]), .CK(clk_80mhz), .Q(d2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i63.GSR = "ENABLED";
    FD1S3AX d2_i64 (.D(d2_71__N_490[64]), .CK(clk_80mhz), .Q(d2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i64.GSR = "ENABLED";
    FD1S3AX d2_i65 (.D(d2_71__N_490[65]), .CK(clk_80mhz), .Q(d2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i65.GSR = "ENABLED";
    FD1S3AX d2_i66 (.D(d2_71__N_490[66]), .CK(clk_80mhz), .Q(d2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i66.GSR = "ENABLED";
    FD1S3AX d2_i67 (.D(d2_71__N_490[67]), .CK(clk_80mhz), .Q(d2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i67.GSR = "ENABLED";
    FD1S3AX d2_i68 (.D(d2_71__N_490[68]), .CK(clk_80mhz), .Q(d2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i68.GSR = "ENABLED";
    FD1S3AX d2_i69 (.D(d2_71__N_490[69]), .CK(clk_80mhz), .Q(d2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i69.GSR = "ENABLED";
    FD1S3AX d2_i70 (.D(d2_71__N_490[70]), .CK(clk_80mhz), .Q(d2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i70.GSR = "ENABLED";
    FD1S3AX d2_i71 (.D(d2_71__N_490[71]), .CK(clk_80mhz), .Q(d2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d2_i71.GSR = "ENABLED";
    FD1S3AX d3_i1 (.D(d3_71__N_562[1]), .CK(clk_80mhz), .Q(d3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i1.GSR = "ENABLED";
    FD1S3AX d3_i2 (.D(d3_71__N_562[2]), .CK(clk_80mhz), .Q(d3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i2.GSR = "ENABLED";
    FD1S3AX d3_i3 (.D(d3_71__N_562[3]), .CK(clk_80mhz), .Q(d3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i3.GSR = "ENABLED";
    FD1S3AX d3_i4 (.D(d3_71__N_562[4]), .CK(clk_80mhz), .Q(d3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i4.GSR = "ENABLED";
    FD1S3AX d3_i5 (.D(d3_71__N_562[5]), .CK(clk_80mhz), .Q(d3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i5.GSR = "ENABLED";
    FD1S3AX d3_i6 (.D(d3_71__N_562[6]), .CK(clk_80mhz), .Q(d3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i6.GSR = "ENABLED";
    FD1S3AX d3_i7 (.D(d3_71__N_562[7]), .CK(clk_80mhz), .Q(d3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i7.GSR = "ENABLED";
    FD1S3AX d3_i8 (.D(d3_71__N_562[8]), .CK(clk_80mhz), .Q(d3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i8.GSR = "ENABLED";
    FD1S3AX d3_i9 (.D(d3_71__N_562[9]), .CK(clk_80mhz), .Q(d3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i9.GSR = "ENABLED";
    FD1S3AX d3_i10 (.D(d3_71__N_562[10]), .CK(clk_80mhz), .Q(d3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i10.GSR = "ENABLED";
    FD1S3AX d3_i11 (.D(d3_71__N_562[11]), .CK(clk_80mhz), .Q(d3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i11.GSR = "ENABLED";
    FD1S3AX d3_i12 (.D(d3_71__N_562[12]), .CK(clk_80mhz), .Q(d3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i12.GSR = "ENABLED";
    FD1S3AX d3_i13 (.D(d3_71__N_562[13]), .CK(clk_80mhz), .Q(d3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i13.GSR = "ENABLED";
    FD1S3AX d3_i14 (.D(d3_71__N_562[14]), .CK(clk_80mhz), .Q(d3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i14.GSR = "ENABLED";
    FD1S3AX d3_i15 (.D(d3_71__N_562[15]), .CK(clk_80mhz), .Q(d3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i15.GSR = "ENABLED";
    FD1S3AX d3_i16 (.D(d3_71__N_562[16]), .CK(clk_80mhz), .Q(d3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i16.GSR = "ENABLED";
    FD1S3AX d3_i17 (.D(d3_71__N_562[17]), .CK(clk_80mhz), .Q(d3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i17.GSR = "ENABLED";
    FD1S3AX d3_i18 (.D(d3_71__N_562[18]), .CK(clk_80mhz), .Q(d3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i18.GSR = "ENABLED";
    FD1S3AX d3_i19 (.D(d3_71__N_562[19]), .CK(clk_80mhz), .Q(d3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i19.GSR = "ENABLED";
    FD1S3AX d3_i20 (.D(d3_71__N_562[20]), .CK(clk_80mhz), .Q(d3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i20.GSR = "ENABLED";
    FD1S3AX d3_i21 (.D(d3_71__N_562[21]), .CK(clk_80mhz), .Q(d3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i21.GSR = "ENABLED";
    FD1S3AX d3_i22 (.D(d3_71__N_562[22]), .CK(clk_80mhz), .Q(d3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i22.GSR = "ENABLED";
    FD1S3AX d3_i23 (.D(d3_71__N_562[23]), .CK(clk_80mhz), .Q(d3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i23.GSR = "ENABLED";
    FD1S3AX d3_i24 (.D(d3_71__N_562[24]), .CK(clk_80mhz), .Q(d3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i24.GSR = "ENABLED";
    FD1S3AX d3_i25 (.D(d3_71__N_562[25]), .CK(clk_80mhz), .Q(d3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i25.GSR = "ENABLED";
    FD1S3AX d3_i26 (.D(d3_71__N_562[26]), .CK(clk_80mhz), .Q(d3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i26.GSR = "ENABLED";
    FD1S3AX d3_i27 (.D(d3_71__N_562[27]), .CK(clk_80mhz), .Q(d3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i27.GSR = "ENABLED";
    FD1S3AX d3_i28 (.D(d3_71__N_562[28]), .CK(clk_80mhz), .Q(d3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i28.GSR = "ENABLED";
    FD1S3AX d3_i29 (.D(d3_71__N_562[29]), .CK(clk_80mhz), .Q(d3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i29.GSR = "ENABLED";
    FD1S3AX d3_i30 (.D(d3_71__N_562[30]), .CK(clk_80mhz), .Q(d3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i30.GSR = "ENABLED";
    FD1S3AX d3_i31 (.D(d3_71__N_562[31]), .CK(clk_80mhz), .Q(d3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i31.GSR = "ENABLED";
    FD1S3AX d3_i32 (.D(d3_71__N_562[32]), .CK(clk_80mhz), .Q(d3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i32.GSR = "ENABLED";
    FD1S3AX d3_i33 (.D(d3_71__N_562[33]), .CK(clk_80mhz), .Q(d3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i33.GSR = "ENABLED";
    FD1S3AX d3_i34 (.D(d3_71__N_562[34]), .CK(clk_80mhz), .Q(d3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i34.GSR = "ENABLED";
    FD1S3AX d3_i35 (.D(d3_71__N_562[35]), .CK(clk_80mhz), .Q(d3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i35.GSR = "ENABLED";
    FD1S3AX d3_i36 (.D(d3_71__N_562[36]), .CK(clk_80mhz), .Q(d3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i36.GSR = "ENABLED";
    FD1S3AX d3_i37 (.D(d3_71__N_562[37]), .CK(clk_80mhz), .Q(d3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i37.GSR = "ENABLED";
    FD1S3AX d3_i38 (.D(d3_71__N_562[38]), .CK(clk_80mhz), .Q(d3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i38.GSR = "ENABLED";
    FD1S3AX d3_i39 (.D(d3_71__N_562[39]), .CK(clk_80mhz), .Q(d3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i39.GSR = "ENABLED";
    FD1S3AX d3_i40 (.D(d3_71__N_562[40]), .CK(clk_80mhz), .Q(d3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i40.GSR = "ENABLED";
    FD1S3AX d3_i41 (.D(d3_71__N_562[41]), .CK(clk_80mhz), .Q(d3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i41.GSR = "ENABLED";
    FD1S3AX d3_i42 (.D(d3_71__N_562[42]), .CK(clk_80mhz), .Q(d3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i42.GSR = "ENABLED";
    FD1S3AX d3_i43 (.D(d3_71__N_562[43]), .CK(clk_80mhz), .Q(d3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i43.GSR = "ENABLED";
    FD1S3AX d3_i44 (.D(d3_71__N_562[44]), .CK(clk_80mhz), .Q(d3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i44.GSR = "ENABLED";
    FD1S3AX d3_i45 (.D(d3_71__N_562[45]), .CK(clk_80mhz), .Q(d3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i45.GSR = "ENABLED";
    FD1S3AX d3_i46 (.D(d3_71__N_562[46]), .CK(clk_80mhz), .Q(d3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i46.GSR = "ENABLED";
    FD1S3AX d3_i47 (.D(d3_71__N_562[47]), .CK(clk_80mhz), .Q(d3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i47.GSR = "ENABLED";
    FD1S3AX d3_i48 (.D(d3_71__N_562[48]), .CK(clk_80mhz), .Q(d3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i48.GSR = "ENABLED";
    FD1S3AX d3_i49 (.D(d3_71__N_562[49]), .CK(clk_80mhz), .Q(d3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i49.GSR = "ENABLED";
    FD1S3AX d3_i50 (.D(d3_71__N_562[50]), .CK(clk_80mhz), .Q(d3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i50.GSR = "ENABLED";
    FD1S3AX d3_i51 (.D(d3_71__N_562[51]), .CK(clk_80mhz), .Q(d3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i51.GSR = "ENABLED";
    FD1S3AX d3_i52 (.D(d3_71__N_562[52]), .CK(clk_80mhz), .Q(d3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i52.GSR = "ENABLED";
    FD1S3AX d3_i53 (.D(d3_71__N_562[53]), .CK(clk_80mhz), .Q(d3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i53.GSR = "ENABLED";
    FD1S3AX d3_i54 (.D(d3_71__N_562[54]), .CK(clk_80mhz), .Q(d3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i54.GSR = "ENABLED";
    FD1S3AX d3_i55 (.D(d3_71__N_562[55]), .CK(clk_80mhz), .Q(d3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i55.GSR = "ENABLED";
    FD1S3AX d3_i56 (.D(d3_71__N_562[56]), .CK(clk_80mhz), .Q(d3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i56.GSR = "ENABLED";
    FD1S3AX d3_i57 (.D(d3_71__N_562[57]), .CK(clk_80mhz), .Q(d3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i57.GSR = "ENABLED";
    FD1S3AX d3_i58 (.D(d3_71__N_562[58]), .CK(clk_80mhz), .Q(d3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i58.GSR = "ENABLED";
    FD1S3AX d3_i59 (.D(d3_71__N_562[59]), .CK(clk_80mhz), .Q(d3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i59.GSR = "ENABLED";
    FD1S3AX d3_i60 (.D(d3_71__N_562[60]), .CK(clk_80mhz), .Q(d3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i60.GSR = "ENABLED";
    FD1S3AX d3_i61 (.D(d3_71__N_562[61]), .CK(clk_80mhz), .Q(d3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i61.GSR = "ENABLED";
    FD1S3AX d3_i62 (.D(d3_71__N_562[62]), .CK(clk_80mhz), .Q(d3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i62.GSR = "ENABLED";
    FD1S3AX d3_i63 (.D(d3_71__N_562[63]), .CK(clk_80mhz), .Q(d3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i63.GSR = "ENABLED";
    FD1S3AX d3_i64 (.D(d3_71__N_562[64]), .CK(clk_80mhz), .Q(d3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i64.GSR = "ENABLED";
    FD1S3AX d3_i65 (.D(d3_71__N_562[65]), .CK(clk_80mhz), .Q(d3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i65.GSR = "ENABLED";
    FD1S3AX d3_i66 (.D(d3_71__N_562[66]), .CK(clk_80mhz), .Q(d3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i66.GSR = "ENABLED";
    FD1S3AX d3_i67 (.D(d3_71__N_562[67]), .CK(clk_80mhz), .Q(d3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i67.GSR = "ENABLED";
    FD1S3AX d3_i68 (.D(d3_71__N_562[68]), .CK(clk_80mhz), .Q(d3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i68.GSR = "ENABLED";
    FD1S3AX d3_i69 (.D(d3_71__N_562[69]), .CK(clk_80mhz), .Q(d3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i69.GSR = "ENABLED";
    FD1S3AX d3_i70 (.D(d3_71__N_562[70]), .CK(clk_80mhz), .Q(d3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i70.GSR = "ENABLED";
    FD1S3AX d3_i71 (.D(d3_71__N_562[71]), .CK(clk_80mhz), .Q(d3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d3_i71.GSR = "ENABLED";
    FD1S3AX d4_i1 (.D(d4_71__N_634[1]), .CK(clk_80mhz), .Q(d4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i1.GSR = "ENABLED";
    FD1S3AX d4_i2 (.D(d4_71__N_634[2]), .CK(clk_80mhz), .Q(d4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i2.GSR = "ENABLED";
    FD1S3AX d4_i3 (.D(d4_71__N_634[3]), .CK(clk_80mhz), .Q(d4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i3.GSR = "ENABLED";
    FD1S3AX d4_i4 (.D(d4_71__N_634[4]), .CK(clk_80mhz), .Q(d4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i4.GSR = "ENABLED";
    FD1S3AX d4_i5 (.D(d4_71__N_634[5]), .CK(clk_80mhz), .Q(d4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i5.GSR = "ENABLED";
    FD1S3AX d4_i6 (.D(d4_71__N_634[6]), .CK(clk_80mhz), .Q(d4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i6.GSR = "ENABLED";
    FD1S3AX d4_i7 (.D(d4_71__N_634[7]), .CK(clk_80mhz), .Q(d4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i7.GSR = "ENABLED";
    FD1S3AX d4_i8 (.D(d4_71__N_634[8]), .CK(clk_80mhz), .Q(d4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i8.GSR = "ENABLED";
    FD1S3AX d4_i9 (.D(d4_71__N_634[9]), .CK(clk_80mhz), .Q(d4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i9.GSR = "ENABLED";
    FD1S3AX d4_i10 (.D(d4_71__N_634[10]), .CK(clk_80mhz), .Q(d4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i10.GSR = "ENABLED";
    FD1S3AX d4_i11 (.D(d4_71__N_634[11]), .CK(clk_80mhz), .Q(d4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i11.GSR = "ENABLED";
    FD1S3AX d4_i12 (.D(d4_71__N_634[12]), .CK(clk_80mhz), .Q(d4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i12.GSR = "ENABLED";
    FD1S3AX d4_i13 (.D(d4_71__N_634[13]), .CK(clk_80mhz), .Q(d4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i13.GSR = "ENABLED";
    FD1S3AX d4_i14 (.D(d4_71__N_634[14]), .CK(clk_80mhz), .Q(d4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i14.GSR = "ENABLED";
    FD1S3AX d4_i15 (.D(d4_71__N_634[15]), .CK(clk_80mhz), .Q(d4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i15.GSR = "ENABLED";
    FD1S3AX d4_i16 (.D(d4_71__N_634[16]), .CK(clk_80mhz), .Q(d4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i16.GSR = "ENABLED";
    FD1S3AX d4_i17 (.D(d4_71__N_634[17]), .CK(clk_80mhz), .Q(d4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i17.GSR = "ENABLED";
    FD1S3AX d4_i18 (.D(d4_71__N_634[18]), .CK(clk_80mhz), .Q(d4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i18.GSR = "ENABLED";
    FD1S3AX d4_i19 (.D(d4_71__N_634[19]), .CK(clk_80mhz), .Q(d4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i19.GSR = "ENABLED";
    FD1S3AX d4_i20 (.D(d4_71__N_634[20]), .CK(clk_80mhz), .Q(d4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i20.GSR = "ENABLED";
    FD1S3AX d4_i21 (.D(d4_71__N_634[21]), .CK(clk_80mhz), .Q(d4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i21.GSR = "ENABLED";
    FD1S3AX d4_i22 (.D(d4_71__N_634[22]), .CK(clk_80mhz), .Q(d4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i22.GSR = "ENABLED";
    FD1S3AX d4_i23 (.D(d4_71__N_634[23]), .CK(clk_80mhz), .Q(d4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i23.GSR = "ENABLED";
    FD1S3AX d4_i24 (.D(d4_71__N_634[24]), .CK(clk_80mhz), .Q(d4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i24.GSR = "ENABLED";
    FD1S3AX d4_i25 (.D(d4_71__N_634[25]), .CK(clk_80mhz), .Q(d4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i25.GSR = "ENABLED";
    FD1S3AX d4_i26 (.D(d4_71__N_634[26]), .CK(clk_80mhz), .Q(d4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i26.GSR = "ENABLED";
    FD1S3AX d4_i27 (.D(d4_71__N_634[27]), .CK(clk_80mhz), .Q(d4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i27.GSR = "ENABLED";
    FD1S3AX d4_i28 (.D(d4_71__N_634[28]), .CK(clk_80mhz), .Q(d4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i28.GSR = "ENABLED";
    FD1S3AX d4_i29 (.D(d4_71__N_634[29]), .CK(clk_80mhz), .Q(d4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i29.GSR = "ENABLED";
    FD1S3AX d4_i30 (.D(d4_71__N_634[30]), .CK(clk_80mhz), .Q(d4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i30.GSR = "ENABLED";
    FD1S3AX d4_i31 (.D(d4_71__N_634[31]), .CK(clk_80mhz), .Q(d4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i31.GSR = "ENABLED";
    FD1S3AX d4_i32 (.D(d4_71__N_634[32]), .CK(clk_80mhz), .Q(d4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i32.GSR = "ENABLED";
    FD1S3AX d4_i33 (.D(d4_71__N_634[33]), .CK(clk_80mhz), .Q(d4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i33.GSR = "ENABLED";
    FD1S3AX d4_i34 (.D(d4_71__N_634[34]), .CK(clk_80mhz), .Q(d4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i34.GSR = "ENABLED";
    FD1S3AX d4_i35 (.D(d4_71__N_634[35]), .CK(clk_80mhz), .Q(d4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i35.GSR = "ENABLED";
    FD1S3AX d4_i36 (.D(d4_71__N_634[36]), .CK(clk_80mhz), .Q(d4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i36.GSR = "ENABLED";
    FD1S3AX d4_i37 (.D(d4_71__N_634[37]), .CK(clk_80mhz), .Q(d4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i37.GSR = "ENABLED";
    FD1S3AX d4_i38 (.D(d4_71__N_634[38]), .CK(clk_80mhz), .Q(d4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i38.GSR = "ENABLED";
    FD1S3AX d4_i39 (.D(d4_71__N_634[39]), .CK(clk_80mhz), .Q(d4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i39.GSR = "ENABLED";
    FD1S3AX d4_i40 (.D(d4_71__N_634[40]), .CK(clk_80mhz), .Q(d4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i40.GSR = "ENABLED";
    FD1S3AX d4_i41 (.D(d4_71__N_634[41]), .CK(clk_80mhz), .Q(d4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i41.GSR = "ENABLED";
    FD1S3AX d4_i42 (.D(d4_71__N_634[42]), .CK(clk_80mhz), .Q(d4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i42.GSR = "ENABLED";
    FD1S3AX d4_i43 (.D(d4_71__N_634[43]), .CK(clk_80mhz), .Q(d4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i43.GSR = "ENABLED";
    FD1S3AX d4_i44 (.D(d4_71__N_634[44]), .CK(clk_80mhz), .Q(d4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i44.GSR = "ENABLED";
    FD1S3AX d4_i45 (.D(d4_71__N_634[45]), .CK(clk_80mhz), .Q(d4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i45.GSR = "ENABLED";
    FD1S3AX d4_i46 (.D(d4_71__N_634[46]), .CK(clk_80mhz), .Q(d4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i46.GSR = "ENABLED";
    FD1S3AX d4_i47 (.D(d4_71__N_634[47]), .CK(clk_80mhz), .Q(d4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i47.GSR = "ENABLED";
    FD1S3AX d4_i48 (.D(d4_71__N_634[48]), .CK(clk_80mhz), .Q(d4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i48.GSR = "ENABLED";
    FD1S3AX d4_i49 (.D(d4_71__N_634[49]), .CK(clk_80mhz), .Q(d4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i49.GSR = "ENABLED";
    FD1S3AX d4_i50 (.D(d4_71__N_634[50]), .CK(clk_80mhz), .Q(d4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i50.GSR = "ENABLED";
    FD1S3AX d4_i51 (.D(d4_71__N_634[51]), .CK(clk_80mhz), .Q(d4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i51.GSR = "ENABLED";
    FD1S3AX d4_i52 (.D(d4_71__N_634[52]), .CK(clk_80mhz), .Q(d4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i52.GSR = "ENABLED";
    FD1S3AX d4_i53 (.D(d4_71__N_634[53]), .CK(clk_80mhz), .Q(d4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i53.GSR = "ENABLED";
    FD1S3AX d4_i54 (.D(d4_71__N_634[54]), .CK(clk_80mhz), .Q(d4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i54.GSR = "ENABLED";
    FD1S3AX d4_i55 (.D(d4_71__N_634[55]), .CK(clk_80mhz), .Q(d4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i55.GSR = "ENABLED";
    FD1S3AX d4_i56 (.D(d4_71__N_634[56]), .CK(clk_80mhz), .Q(d4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i56.GSR = "ENABLED";
    FD1S3AX d4_i57 (.D(d4_71__N_634[57]), .CK(clk_80mhz), .Q(d4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i57.GSR = "ENABLED";
    FD1S3AX d4_i58 (.D(d4_71__N_634[58]), .CK(clk_80mhz), .Q(d4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i58.GSR = "ENABLED";
    FD1S3AX d4_i59 (.D(d4_71__N_634[59]), .CK(clk_80mhz), .Q(d4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i59.GSR = "ENABLED";
    FD1S3AX d4_i60 (.D(d4_71__N_634[60]), .CK(clk_80mhz), .Q(d4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i60.GSR = "ENABLED";
    FD1S3AX d4_i61 (.D(d4_71__N_634[61]), .CK(clk_80mhz), .Q(d4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i61.GSR = "ENABLED";
    FD1S3AX d4_i62 (.D(d4_71__N_634[62]), .CK(clk_80mhz), .Q(d4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i62.GSR = "ENABLED";
    FD1S3AX d4_i63 (.D(d4_71__N_634[63]), .CK(clk_80mhz), .Q(d4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i63.GSR = "ENABLED";
    FD1S3AX d4_i64 (.D(d4_71__N_634[64]), .CK(clk_80mhz), .Q(d4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i64.GSR = "ENABLED";
    FD1S3AX d4_i65 (.D(d4_71__N_634[65]), .CK(clk_80mhz), .Q(d4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i65.GSR = "ENABLED";
    FD1S3AX d4_i66 (.D(d4_71__N_634[66]), .CK(clk_80mhz), .Q(d4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i66.GSR = "ENABLED";
    FD1S3AX d4_i67 (.D(d4_71__N_634[67]), .CK(clk_80mhz), .Q(d4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i67.GSR = "ENABLED";
    FD1S3AX d4_i68 (.D(d4_71__N_634[68]), .CK(clk_80mhz), .Q(d4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i68.GSR = "ENABLED";
    FD1S3AX d4_i69 (.D(d4_71__N_634[69]), .CK(clk_80mhz), .Q(d4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i69.GSR = "ENABLED";
    FD1S3AX d4_i70 (.D(d4_71__N_634[70]), .CK(clk_80mhz), .Q(d4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i70.GSR = "ENABLED";
    FD1S3AX d4_i71 (.D(d4_71__N_634[71]), .CK(clk_80mhz), .Q(d4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d4_i71.GSR = "ENABLED";
    FD1S3AX d5_i1 (.D(d5_71__N_706[1]), .CK(clk_80mhz), .Q(d5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i1.GSR = "ENABLED";
    FD1S3AX d5_i2 (.D(d5_71__N_706[2]), .CK(clk_80mhz), .Q(d5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i2.GSR = "ENABLED";
    FD1S3AX d5_i3 (.D(d5_71__N_706[3]), .CK(clk_80mhz), .Q(d5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i3.GSR = "ENABLED";
    FD1S3AX d5_i4 (.D(d5_71__N_706[4]), .CK(clk_80mhz), .Q(d5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i4.GSR = "ENABLED";
    FD1S3AX d5_i5 (.D(d5_71__N_706[5]), .CK(clk_80mhz), .Q(d5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i5.GSR = "ENABLED";
    FD1S3AX d5_i6 (.D(d5_71__N_706[6]), .CK(clk_80mhz), .Q(d5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i6.GSR = "ENABLED";
    FD1S3AX d5_i7 (.D(d5_71__N_706[7]), .CK(clk_80mhz), .Q(d5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i7.GSR = "ENABLED";
    FD1S3AX d5_i8 (.D(d5_71__N_706[8]), .CK(clk_80mhz), .Q(d5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i8.GSR = "ENABLED";
    FD1S3AX d5_i9 (.D(d5_71__N_706[9]), .CK(clk_80mhz), .Q(d5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i9.GSR = "ENABLED";
    FD1S3AX d5_i10 (.D(d5_71__N_706[10]), .CK(clk_80mhz), .Q(d5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i10.GSR = "ENABLED";
    FD1S3AX d5_i11 (.D(d5_71__N_706[11]), .CK(clk_80mhz), .Q(d5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i11.GSR = "ENABLED";
    FD1S3AX d5_i12 (.D(d5_71__N_706[12]), .CK(clk_80mhz), .Q(d5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i12.GSR = "ENABLED";
    FD1S3AX d5_i13 (.D(d5_71__N_706[13]), .CK(clk_80mhz), .Q(d5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i13.GSR = "ENABLED";
    FD1S3AX d5_i14 (.D(d5_71__N_706[14]), .CK(clk_80mhz), .Q(d5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i14.GSR = "ENABLED";
    FD1S3AX d5_i15 (.D(d5_71__N_706[15]), .CK(clk_80mhz), .Q(d5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i15.GSR = "ENABLED";
    FD1S3AX d5_i16 (.D(d5_71__N_706[16]), .CK(clk_80mhz), .Q(d5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i16.GSR = "ENABLED";
    FD1S3AX d5_i17 (.D(d5_71__N_706[17]), .CK(clk_80mhz), .Q(d5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i17.GSR = "ENABLED";
    FD1S3AX d5_i18 (.D(d5_71__N_706[18]), .CK(clk_80mhz), .Q(d5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i18.GSR = "ENABLED";
    FD1S3AX d5_i19 (.D(d5_71__N_706[19]), .CK(clk_80mhz), .Q(d5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i19.GSR = "ENABLED";
    FD1S3AX d5_i20 (.D(d5_71__N_706[20]), .CK(clk_80mhz), .Q(d5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i20.GSR = "ENABLED";
    FD1S3AX d5_i21 (.D(d5_71__N_706[21]), .CK(clk_80mhz), .Q(d5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i21.GSR = "ENABLED";
    FD1S3AX d5_i22 (.D(d5_71__N_706[22]), .CK(clk_80mhz), .Q(d5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i22.GSR = "ENABLED";
    FD1S3AX d5_i23 (.D(d5_71__N_706[23]), .CK(clk_80mhz), .Q(d5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i23.GSR = "ENABLED";
    FD1S3AX d5_i24 (.D(d5_71__N_706[24]), .CK(clk_80mhz), .Q(d5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i24.GSR = "ENABLED";
    FD1S3AX d5_i25 (.D(d5_71__N_706[25]), .CK(clk_80mhz), .Q(d5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i25.GSR = "ENABLED";
    FD1S3AX d5_i26 (.D(d5_71__N_706[26]), .CK(clk_80mhz), .Q(d5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i26.GSR = "ENABLED";
    FD1S3AX d5_i27 (.D(d5_71__N_706[27]), .CK(clk_80mhz), .Q(d5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i27.GSR = "ENABLED";
    FD1S3AX d5_i28 (.D(d5_71__N_706[28]), .CK(clk_80mhz), .Q(d5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i28.GSR = "ENABLED";
    FD1S3AX d5_i29 (.D(d5_71__N_706[29]), .CK(clk_80mhz), .Q(d5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i29.GSR = "ENABLED";
    FD1S3AX d5_i30 (.D(d5_71__N_706[30]), .CK(clk_80mhz), .Q(d5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i30.GSR = "ENABLED";
    FD1S3AX d5_i31 (.D(d5_71__N_706[31]), .CK(clk_80mhz), .Q(d5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i31.GSR = "ENABLED";
    FD1S3AX d5_i32 (.D(d5_71__N_706[32]), .CK(clk_80mhz), .Q(d5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i32.GSR = "ENABLED";
    FD1S3AX d5_i33 (.D(d5_71__N_706[33]), .CK(clk_80mhz), .Q(d5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i33.GSR = "ENABLED";
    FD1S3AX d5_i34 (.D(d5_71__N_706[34]), .CK(clk_80mhz), .Q(d5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i34.GSR = "ENABLED";
    FD1S3AX d5_i35 (.D(d5_71__N_706[35]), .CK(clk_80mhz), .Q(d5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i35.GSR = "ENABLED";
    FD1S3AX d5_i36 (.D(d5_71__N_706[36]), .CK(clk_80mhz), .Q(d5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i36.GSR = "ENABLED";
    FD1S3AX d5_i37 (.D(d5_71__N_706[37]), .CK(clk_80mhz), .Q(d5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i37.GSR = "ENABLED";
    FD1S3AX d5_i38 (.D(d5_71__N_706[38]), .CK(clk_80mhz), .Q(d5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i38.GSR = "ENABLED";
    FD1S3AX d5_i39 (.D(d5_71__N_706[39]), .CK(clk_80mhz), .Q(d5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i39.GSR = "ENABLED";
    FD1S3AX d5_i40 (.D(d5_71__N_706[40]), .CK(clk_80mhz), .Q(d5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i40.GSR = "ENABLED";
    FD1S3AX d5_i41 (.D(d5_71__N_706[41]), .CK(clk_80mhz), .Q(d5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i41.GSR = "ENABLED";
    FD1S3AX d5_i42 (.D(d5_71__N_706[42]), .CK(clk_80mhz), .Q(d5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i42.GSR = "ENABLED";
    FD1S3AX d5_i43 (.D(d5_71__N_706[43]), .CK(clk_80mhz), .Q(d5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i43.GSR = "ENABLED";
    FD1S3AX d5_i44 (.D(d5_71__N_706[44]), .CK(clk_80mhz), .Q(d5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i44.GSR = "ENABLED";
    FD1S3AX d5_i45 (.D(d5_71__N_706[45]), .CK(clk_80mhz), .Q(d5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i45.GSR = "ENABLED";
    FD1S3AX d5_i46 (.D(d5_71__N_706[46]), .CK(clk_80mhz), .Q(d5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i46.GSR = "ENABLED";
    FD1S3AX d5_i47 (.D(d5_71__N_706[47]), .CK(clk_80mhz), .Q(d5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i47.GSR = "ENABLED";
    FD1S3AX d5_i48 (.D(d5_71__N_706[48]), .CK(clk_80mhz), .Q(d5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i48.GSR = "ENABLED";
    FD1S3AX d5_i49 (.D(d5_71__N_706[49]), .CK(clk_80mhz), .Q(d5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i49.GSR = "ENABLED";
    FD1S3AX d5_i50 (.D(d5_71__N_706[50]), .CK(clk_80mhz), .Q(d5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i50.GSR = "ENABLED";
    FD1S3AX d5_i51 (.D(d5_71__N_706[51]), .CK(clk_80mhz), .Q(d5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i51.GSR = "ENABLED";
    FD1S3AX d5_i52 (.D(d5_71__N_706[52]), .CK(clk_80mhz), .Q(d5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i52.GSR = "ENABLED";
    FD1S3AX d5_i53 (.D(d5_71__N_706[53]), .CK(clk_80mhz), .Q(d5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i53.GSR = "ENABLED";
    FD1S3AX d5_i54 (.D(d5_71__N_706[54]), .CK(clk_80mhz), .Q(d5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i54.GSR = "ENABLED";
    FD1S3AX d5_i55 (.D(d5_71__N_706[55]), .CK(clk_80mhz), .Q(d5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i55.GSR = "ENABLED";
    FD1S3AX d5_i56 (.D(d5_71__N_706[56]), .CK(clk_80mhz), .Q(d5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i56.GSR = "ENABLED";
    FD1S3AX d5_i57 (.D(d5_71__N_706[57]), .CK(clk_80mhz), .Q(d5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i57.GSR = "ENABLED";
    FD1S3AX d5_i58 (.D(d5_71__N_706[58]), .CK(clk_80mhz), .Q(d5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i58.GSR = "ENABLED";
    FD1S3AX d5_i59 (.D(d5_71__N_706[59]), .CK(clk_80mhz), .Q(d5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i59.GSR = "ENABLED";
    FD1S3AX d5_i60 (.D(d5_71__N_706[60]), .CK(clk_80mhz), .Q(d5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i60.GSR = "ENABLED";
    FD1S3AX d5_i61 (.D(d5_71__N_706[61]), .CK(clk_80mhz), .Q(d5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i61.GSR = "ENABLED";
    FD1S3AX d5_i62 (.D(d5_71__N_706[62]), .CK(clk_80mhz), .Q(d5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i62.GSR = "ENABLED";
    FD1S3AX d5_i63 (.D(d5_71__N_706[63]), .CK(clk_80mhz), .Q(d5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i63.GSR = "ENABLED";
    FD1S3AX d5_i64 (.D(d5_71__N_706[64]), .CK(clk_80mhz), .Q(d5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i64.GSR = "ENABLED";
    FD1S3AX d5_i65 (.D(d5_71__N_706[65]), .CK(clk_80mhz), .Q(d5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i65.GSR = "ENABLED";
    FD1S3AX d5_i66 (.D(d5_71__N_706[66]), .CK(clk_80mhz), .Q(d5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i66.GSR = "ENABLED";
    FD1S3AX d5_i67 (.D(d5_71__N_706[67]), .CK(clk_80mhz), .Q(d5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i67.GSR = "ENABLED";
    FD1S3AX d5_i68 (.D(d5_71__N_706[68]), .CK(clk_80mhz), .Q(d5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i68.GSR = "ENABLED";
    FD1S3AX d5_i69 (.D(d5_71__N_706[69]), .CK(clk_80mhz), .Q(d5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i69.GSR = "ENABLED";
    FD1S3AX d5_i70 (.D(d5_71__N_706[70]), .CK(clk_80mhz), .Q(d5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i70.GSR = "ENABLED";
    FD1S3AX d5_i71 (.D(d5_71__N_706[71]), .CK(clk_80mhz), .Q(d5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d5_i71.GSR = "ENABLED";
    FD1P3AX d6_i0_i1 (.D(d6_71__N_1459[1]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d6_i0_i2 (.D(d6_71__N_1459[2]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d6_i0_i3 (.D(d6_71__N_1459[3]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d6_i0_i4 (.D(d6_71__N_1459[4]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d6_i0_i5 (.D(d6_71__N_1459[5]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d6_i0_i6 (.D(d6_71__N_1459[6]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d6_i0_i7 (.D(d6_71__N_1459[7]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d6_i0_i8 (.D(d6_71__N_1459[8]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d6_i0_i9 (.D(d6_71__N_1459[9]), .SP(clk_80mhz_enable_149), .CK(clk_80mhz), 
            .Q(d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d6_i0_i10 (.D(d6_71__N_1459[10]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d6_i0_i11 (.D(d6_71__N_1459[11]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d6_i0_i12 (.D(d6_71__N_1459[12]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d6_i0_i13 (.D(d6_71__N_1459[13]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d6_i0_i14 (.D(d6_71__N_1459[14]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d6_i0_i15 (.D(d6_71__N_1459[15]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d6_i0_i16 (.D(d6_71__N_1459[16]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d6_i0_i17 (.D(d6_71__N_1459[17]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d6_i0_i18 (.D(d6_71__N_1459[18]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d6_i0_i19 (.D(d6_71__N_1459[19]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d6_i0_i20 (.D(d6_71__N_1459[20]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d6_i0_i21 (.D(d6_71__N_1459[21]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d6_i0_i22 (.D(d6_71__N_1459[22]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d6_i0_i23 (.D(d6_71__N_1459[23]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d6_i0_i24 (.D(d6_71__N_1459[24]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d6_i0_i25 (.D(d6_71__N_1459[25]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d6_i0_i26 (.D(d6_71__N_1459[26]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d6_i0_i27 (.D(d6_71__N_1459[27]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d6_i0_i28 (.D(d6_71__N_1459[28]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d6_i0_i29 (.D(d6_71__N_1459[29]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d6_i0_i30 (.D(d6_71__N_1459[30]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d6_i0_i31 (.D(d6_71__N_1459[31]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d6_i0_i32 (.D(d6_71__N_1459[32]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d6_i0_i33 (.D(d6_71__N_1459[33]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d6_i0_i34 (.D(d6_71__N_1459[34]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d6_i0_i35 (.D(d6_71__N_1459[35]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d6_i0_i36 (.D(d6_71__N_1459[36]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d6_i0_i37 (.D(d6_71__N_1459[37]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d6_i0_i38 (.D(d6_71__N_1459[38]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d6_i0_i39 (.D(d6_71__N_1459[39]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d6_i0_i40 (.D(d6_71__N_1459[40]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d6_i0_i41 (.D(d6_71__N_1459[41]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d6_i0_i42 (.D(d6_71__N_1459[42]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d6_i0_i43 (.D(d6_71__N_1459[43]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d6_i0_i44 (.D(d6_71__N_1459[44]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d6_i0_i45 (.D(d6_71__N_1459[45]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d6_i0_i46 (.D(d6_71__N_1459[46]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d6_i0_i47 (.D(d6_71__N_1459[47]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d6_i0_i48 (.D(d6_71__N_1459[48]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d6_i0_i49 (.D(d6_71__N_1459[49]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d6_i0_i50 (.D(d6_71__N_1459[50]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d6_i0_i51 (.D(d6_71__N_1459[51]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d6_i0_i52 (.D(d6_71__N_1459[52]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d6_i0_i53 (.D(d6_71__N_1459[53]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d6_i0_i54 (.D(d6_71__N_1459[54]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d6_i0_i55 (.D(d6_71__N_1459[55]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d6_i0_i56 (.D(d6_71__N_1459[56]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d6_i0_i57 (.D(d6_71__N_1459[57]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d6_i0_i58 (.D(d6_71__N_1459[58]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d6_i0_i59 (.D(d6_71__N_1459[59]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d6_i0_i60 (.D(d6_71__N_1459[60]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d6_i0_i61 (.D(d6_71__N_1459[61]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d6_i0_i62 (.D(d6_71__N_1459[62]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d6_i0_i63 (.D(d6_71__N_1459[63]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d6_i0_i64 (.D(d6_71__N_1459[64]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d6_i0_i65 (.D(d6_71__N_1459[65]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d6_i0_i66 (.D(d6_71__N_1459[66]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d6_i0_i67 (.D(d6_71__N_1459[67]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d6_i0_i68 (.D(d6_71__N_1459[68]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d6_i0_i69 (.D(d6_71__N_1459[69]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d6_i0_i70 (.D(d6_71__N_1459[70]), .SP(clk_80mhz_enable_199), 
            .CK(clk_80mhz), .Q(d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d6_i0_i71 (.D(d6_71__N_1459[71]), .SP(clk_80mhz_enable_249), 
            .CK(clk_80mhz), .Q(d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i1 (.D(d6[1]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i2 (.D(d6[2]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i3 (.D(d6[3]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i4 (.D(d6[4]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i5 (.D(d6[5]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i6 (.D(d6[6]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i7 (.D(d6[7]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i8 (.D(d6[8]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i9 (.D(d6[9]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i10 (.D(d6[10]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i11 (.D(d6[11]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i12 (.D(d6[12]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i13 (.D(d6[13]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i14 (.D(d6[14]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i15 (.D(d6[15]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i16 (.D(d6[16]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i17 (.D(d6[17]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i18 (.D(d6[18]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i19 (.D(d6[19]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i20 (.D(d6[20]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i21 (.D(d6[21]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i22 (.D(d6[22]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i23 (.D(d6[23]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i24 (.D(d6[24]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i25 (.D(d6[25]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i26 (.D(d6[26]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i27 (.D(d6[27]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i28 (.D(d6[28]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i29 (.D(d6[29]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i30 (.D(d6[30]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i31 (.D(d6[31]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i32 (.D(d6[32]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i33 (.D(d6[33]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i34 (.D(d6[34]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i35 (.D(d6[35]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i36 (.D(d6[36]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i37 (.D(d6[37]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i38 (.D(d6[38]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i39 (.D(d6[39]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i40 (.D(d6[40]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i41 (.D(d6[41]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i42 (.D(d6[42]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i43 (.D(d6[43]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i44 (.D(d6[44]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i45 (.D(d6[45]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i46 (.D(d6[46]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i47 (.D(d6[47]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i48 (.D(d6[48]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i49 (.D(d6[49]), .SP(clk_80mhz_enable_249), .CK(clk_80mhz), 
            .Q(d_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i50 (.D(d6[50]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i51 (.D(d6[51]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i52 (.D(d6[52]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i53 (.D(d6[53]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i54 (.D(d6[54]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i55 (.D(d6[55]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i56 (.D(d6[56]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i57 (.D(d6[57]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i58 (.D(d6[58]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i59 (.D(d6[59]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i60 (.D(d6[60]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i61 (.D(d6[61]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i62 (.D(d6[62]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i63 (.D(d6[63]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i64 (.D(d6[64]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i65 (.D(d6[65]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i66 (.D(d6[66]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i67 (.D(d6[67]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i68 (.D(d6[68]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i69 (.D(d6[69]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i70 (.D(d6[70]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d6_i0_i71 (.D(d6[71]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX d7_i0_i1 (.D(d7_71__N_1531[1]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d7_i0_i2 (.D(d7_71__N_1531[2]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d7_i0_i3 (.D(d7_71__N_1531[3]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d7_i0_i4 (.D(d7_71__N_1531[4]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d7_i0_i5 (.D(d7_71__N_1531[5]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d7_i0_i6 (.D(d7_71__N_1531[6]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d7_i0_i7 (.D(d7_71__N_1531[7]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d7_i0_i8 (.D(d7_71__N_1531[8]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d7_i0_i9 (.D(d7_71__N_1531[9]), .SP(clk_80mhz_enable_299), .CK(clk_80mhz), 
            .Q(d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d7_i0_i10 (.D(d7_71__N_1531[10]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d7_i0_i11 (.D(d7_71__N_1531[11]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d7_i0_i12 (.D(d7_71__N_1531[12]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d7_i0_i13 (.D(d7_71__N_1531[13]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d7_i0_i14 (.D(d7_71__N_1531[14]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d7_i0_i15 (.D(d7_71__N_1531[15]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d7_i0_i16 (.D(d7_71__N_1531[16]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d7_i0_i17 (.D(d7_71__N_1531[17]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d7_i0_i18 (.D(d7_71__N_1531[18]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d7_i0_i19 (.D(d7_71__N_1531[19]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d7_i0_i20 (.D(d7_71__N_1531[20]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d7_i0_i21 (.D(d7_71__N_1531[21]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d7_i0_i22 (.D(d7_71__N_1531[22]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d7_i0_i23 (.D(d7_71__N_1531[23]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d7_i0_i24 (.D(d7_71__N_1531[24]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d7_i0_i25 (.D(d7_71__N_1531[25]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d7_i0_i26 (.D(d7_71__N_1531[26]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d7_i0_i27 (.D(d7_71__N_1531[27]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d7_i0_i28 (.D(d7_71__N_1531[28]), .SP(clk_80mhz_enable_299), 
            .CK(clk_80mhz), .Q(d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d7_i0_i29 (.D(d7_71__N_1531[29]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d7_i0_i30 (.D(d7_71__N_1531[30]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d7_i0_i31 (.D(d7_71__N_1531[31]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d7_i0_i32 (.D(d7_71__N_1531[32]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d7_i0_i33 (.D(d7_71__N_1531[33]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d7_i0_i34 (.D(d7_71__N_1531[34]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d7_i0_i35 (.D(d7_71__N_1531[35]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d7_i0_i36 (.D(d7_71__N_1531[36]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d7_i0_i37 (.D(d7_71__N_1531[37]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d7_i0_i38 (.D(d7_71__N_1531[38]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d7_i0_i39 (.D(d7_71__N_1531[39]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d7_i0_i40 (.D(d7_71__N_1531[40]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d7_i0_i41 (.D(d7_71__N_1531[41]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d7_i0_i42 (.D(d7_71__N_1531[42]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d7_i0_i43 (.D(d7_71__N_1531[43]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d7_i0_i44 (.D(d7_71__N_1531[44]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d7_i0_i45 (.D(d7_71__N_1531[45]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d7_i0_i46 (.D(d7_71__N_1531[46]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d7_i0_i47 (.D(d7_71__N_1531[47]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d7_i0_i48 (.D(d7_71__N_1531[48]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d7_i0_i49 (.D(d7_71__N_1531[49]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d7_i0_i50 (.D(d7_71__N_1531[50]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d7_i0_i51 (.D(d7_71__N_1531[51]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d7_i0_i52 (.D(d7_71__N_1531[52]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d7_i0_i53 (.D(d7_71__N_1531[53]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d7_i0_i54 (.D(d7_71__N_1531[54]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d7_i0_i55 (.D(d7_71__N_1531[55]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d7_i0_i56 (.D(d7_71__N_1531[56]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d7_i0_i57 (.D(d7_71__N_1531[57]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d7_i0_i58 (.D(d7_71__N_1531[58]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d7_i0_i59 (.D(d7_71__N_1531[59]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d7_i0_i60 (.D(d7_71__N_1531[60]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d7_i0_i61 (.D(d7_71__N_1531[61]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d7_i0_i62 (.D(d7_71__N_1531[62]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d7_i0_i63 (.D(d7_71__N_1531[63]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d7_i0_i64 (.D(d7_71__N_1531[64]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d7_i0_i65 (.D(d7_71__N_1531[65]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d7_i0_i66 (.D(d7_71__N_1531[66]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d7_i0_i67 (.D(d7_71__N_1531[67]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d7_i0_i68 (.D(d7_71__N_1531[68]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d7_i0_i69 (.D(d7_71__N_1531[69]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d7_i0_i70 (.D(d7_71__N_1531[70]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d7_i0_i71 (.D(d7_71__N_1531[71]), .SP(clk_80mhz_enable_349), 
            .CK(clk_80mhz), .Q(d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i1 (.D(d7[1]), .SP(clk_80mhz_enable_349), .CK(clk_80mhz), 
            .Q(d_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i2 (.D(d7[2]), .SP(clk_80mhz_enable_349), .CK(clk_80mhz), 
            .Q(d_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i3 (.D(d7[3]), .SP(clk_80mhz_enable_349), .CK(clk_80mhz), 
            .Q(d_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i4 (.D(d7[4]), .SP(clk_80mhz_enable_349), .CK(clk_80mhz), 
            .Q(d_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i5 (.D(d7[5]), .SP(clk_80mhz_enable_349), .CK(clk_80mhz), 
            .Q(d_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i6 (.D(d7[6]), .SP(clk_80mhz_enable_349), .CK(clk_80mhz), 
            .Q(d_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i7 (.D(d7[7]), .SP(clk_80mhz_enable_349), .CK(clk_80mhz), 
            .Q(d_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i8 (.D(d7[8]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i9 (.D(d7[9]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i10 (.D(d7[10]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i11 (.D(d7[11]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i12 (.D(d7[12]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i13 (.D(d7[13]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i14 (.D(d7[14]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i15 (.D(d7[15]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i16 (.D(d7[16]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i17 (.D(d7[17]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i18 (.D(d7[18]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i19 (.D(d7[19]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i20 (.D(d7[20]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i21 (.D(d7[21]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i22 (.D(d7[22]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i23 (.D(d7[23]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i24 (.D(d7[24]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i25 (.D(d7[25]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i26 (.D(d7[26]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i27 (.D(d7[27]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i28 (.D(d7[28]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i29 (.D(d7[29]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i30 (.D(d7[30]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i31 (.D(d7[31]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i32 (.D(d7[32]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i33 (.D(d7[33]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i34 (.D(d7[34]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i35 (.D(d7[35]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i36 (.D(d7[36]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i37 (.D(d7[37]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i38 (.D(d7[38]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i39 (.D(d7[39]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i40 (.D(d7[40]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i41 (.D(d7[41]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i42 (.D(d7[42]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i43 (.D(d7[43]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i44 (.D(d7[44]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i45 (.D(d7[45]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i46 (.D(d7[46]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i47 (.D(d7[47]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i48 (.D(d7[48]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i49 (.D(d7[49]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i50 (.D(d7[50]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i51 (.D(d7[51]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i52 (.D(d7[52]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i53 (.D(d7[53]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i54 (.D(d7[54]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i55 (.D(d7[55]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i56 (.D(d7[56]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i57 (.D(d7[57]), .SP(clk_80mhz_enable_399), .CK(clk_80mhz), 
            .Q(d_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i58 (.D(d7[58]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i59 (.D(d7[59]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i60 (.D(d7[60]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i61 (.D(d7[61]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i62 (.D(d7[62]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i63 (.D(d7[63]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i64 (.D(d7[64]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i65 (.D(d7[65]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i66 (.D(d7[66]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i67 (.D(d7[67]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i68 (.D(d7[68]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i69 (.D(d7[69]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i70 (.D(d7[70]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d7_i0_i71 (.D(d7[71]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX d8_i0_i1 (.D(d8_71__N_1603[1]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d8_i0_i2 (.D(d8_71__N_1603[2]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d8_i0_i3 (.D(d8_71__N_1603[3]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d8_i0_i4 (.D(d8_71__N_1603[4]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d8_i0_i5 (.D(d8_71__N_1603[5]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d8_i0_i6 (.D(d8_71__N_1603[6]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d8_i0_i7 (.D(d8_71__N_1603[7]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d8_i0_i8 (.D(d8_71__N_1603[8]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d8_i0_i9 (.D(d8_71__N_1603[9]), .SP(clk_80mhz_enable_449), .CK(clk_80mhz), 
            .Q(d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d8_i0_i10 (.D(d8_71__N_1603[10]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d8_i0_i11 (.D(d8_71__N_1603[11]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d8_i0_i12 (.D(d8_71__N_1603[12]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d8_i0_i13 (.D(d8_71__N_1603[13]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d8_i0_i14 (.D(d8_71__N_1603[14]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d8_i0_i15 (.D(d8_71__N_1603[15]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d8_i0_i16 (.D(d8_71__N_1603[16]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d8_i0_i17 (.D(d8_71__N_1603[17]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d8_i0_i18 (.D(d8_71__N_1603[18]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d8_i0_i19 (.D(d8_71__N_1603[19]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d8_i0_i20 (.D(d8_71__N_1603[20]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d8_i0_i21 (.D(d8_71__N_1603[21]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d8_i0_i22 (.D(d8_71__N_1603[22]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d8_i0_i23 (.D(d8_71__N_1603[23]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d8_i0_i24 (.D(d8_71__N_1603[24]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d8_i0_i25 (.D(d8_71__N_1603[25]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d8_i0_i26 (.D(d8_71__N_1603[26]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d8_i0_i27 (.D(d8_71__N_1603[27]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d8_i0_i28 (.D(d8_71__N_1603[28]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d8_i0_i29 (.D(d8_71__N_1603[29]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d8_i0_i30 (.D(d8_71__N_1603[30]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d8_i0_i31 (.D(d8_71__N_1603[31]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d8_i0_i32 (.D(d8_71__N_1603[32]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d8_i0_i33 (.D(d8_71__N_1603[33]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d8_i0_i34 (.D(d8_71__N_1603[34]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d8_i0_i35 (.D(d8_71__N_1603[35]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d8_i0_i36 (.D(d8_71__N_1603[36]), .SP(clk_80mhz_enable_449), 
            .CK(clk_80mhz), .Q(d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d8_i0_i37 (.D(d8_71__N_1603[37]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d8_i0_i38 (.D(d8_71__N_1603[38]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d8_i0_i39 (.D(d8_71__N_1603[39]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d8_i0_i40 (.D(d8_71__N_1603[40]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d8_i0_i41 (.D(d8_71__N_1603[41]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d8_i0_i42 (.D(d8_71__N_1603[42]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d8_i0_i43 (.D(d8_71__N_1603[43]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d8_i0_i44 (.D(d8_71__N_1603[44]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d8_i0_i45 (.D(d8_71__N_1603[45]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d8_i0_i46 (.D(d8_71__N_1603[46]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d8_i0_i47 (.D(d8_71__N_1603[47]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d8_i0_i48 (.D(d8_71__N_1603[48]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d8_i0_i49 (.D(d8_71__N_1603[49]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d8_i0_i50 (.D(d8_71__N_1603[50]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d8_i0_i51 (.D(d8_71__N_1603[51]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d8_i0_i52 (.D(d8_71__N_1603[52]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d8_i0_i53 (.D(d8_71__N_1603[53]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d8_i0_i54 (.D(d8_71__N_1603[54]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d8_i0_i55 (.D(d8_71__N_1603[55]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d8_i0_i56 (.D(d8_71__N_1603[56]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d8_i0_i57 (.D(d8_71__N_1603[57]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d8_i0_i58 (.D(d8_71__N_1603[58]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d8_i0_i59 (.D(d8_71__N_1603[59]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d8_i0_i60 (.D(d8_71__N_1603[60]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d8_i0_i61 (.D(d8_71__N_1603[61]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d8_i0_i62 (.D(d8_71__N_1603[62]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d8_i0_i63 (.D(d8_71__N_1603[63]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d8_i0_i64 (.D(d8_71__N_1603[64]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d8_i0_i65 (.D(d8_71__N_1603[65]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d8_i0_i66 (.D(d8_71__N_1603[66]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d8_i0_i67 (.D(d8_71__N_1603[67]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d8_i0_i68 (.D(d8_71__N_1603[68]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d8_i0_i69 (.D(d8_71__N_1603[69]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d8_i0_i70 (.D(d8_71__N_1603[70]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d8_i0_i71 (.D(d8_71__N_1603[71]), .SP(clk_80mhz_enable_499), 
            .CK(clk_80mhz), .Q(d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i1 (.D(d8[1]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i2 (.D(d8[2]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i3 (.D(d8[3]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i4 (.D(d8[4]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i5 (.D(d8[5]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i6 (.D(d8[6]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i7 (.D(d8[7]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i8 (.D(d8[8]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i9 (.D(d8[9]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i10 (.D(d8[10]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i11 (.D(d8[11]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i12 (.D(d8[12]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i13 (.D(d8[13]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i14 (.D(d8[14]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i15 (.D(d8[15]), .SP(clk_80mhz_enable_499), .CK(clk_80mhz), 
            .Q(d_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i16 (.D(d8[16]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i17 (.D(d8[17]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i18 (.D(d8[18]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i19 (.D(d8[19]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i20 (.D(d8[20]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i21 (.D(d8[21]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i22 (.D(d8[22]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i23 (.D(d8[23]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i24 (.D(d8[24]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i25 (.D(d8[25]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i26 (.D(d8[26]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i27 (.D(d8[27]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i28 (.D(d8[28]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i29 (.D(d8[29]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i30 (.D(d8[30]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i31 (.D(d8[31]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i32 (.D(d8[32]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i33 (.D(d8[33]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i34 (.D(d8[34]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i35 (.D(d8[35]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i36 (.D(d8[36]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i37 (.D(d8[37]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i38 (.D(d8[38]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i39 (.D(d8[39]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i40 (.D(d8[40]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i41 (.D(d8[41]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i42 (.D(d8[42]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i43 (.D(d8[43]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i44 (.D(d8[44]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i45 (.D(d8[45]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i46 (.D(d8[46]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i47 (.D(d8[47]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i48 (.D(d8[48]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i49 (.D(d8[49]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i50 (.D(d8[50]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i51 (.D(d8[51]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i52 (.D(d8[52]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i53 (.D(d8[53]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i54 (.D(d8[54]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i55 (.D(d8[55]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i56 (.D(d8[56]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i57 (.D(d8[57]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i58 (.D(d8[58]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i59 (.D(d8[59]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i60 (.D(d8[60]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i61 (.D(d8[61]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i62 (.D(d8[62]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i63 (.D(d8[63]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i64 (.D(d8[64]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i65 (.D(d8[65]), .SP(clk_80mhz_enable_549), .CK(clk_80mhz), 
            .Q(d_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i66 (.D(d8[66]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i67 (.D(d8[67]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i68 (.D(d8[68]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i69 (.D(d8[69]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i70 (.D(d8[70]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d8_i0_i71 (.D(d8[71]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX d9_i0_i1 (.D(d9_71__N_1675[1]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d9_i0_i2 (.D(d9_71__N_1675[2]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d9_i0_i3 (.D(d9_71__N_1675[3]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d9_i0_i4 (.D(d9_71__N_1675[4]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d9_i0_i5 (.D(d9_71__N_1675[5]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d9_i0_i6 (.D(d9_71__N_1675[6]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d9_i0_i7 (.D(d9_71__N_1675[7]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d9_i0_i8 (.D(d9_71__N_1675[8]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d9_i0_i9 (.D(d9_71__N_1675[9]), .SP(clk_80mhz_enable_599), .CK(clk_80mhz), 
            .Q(d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d9_i0_i10 (.D(d9_71__N_1675[10]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d9_i0_i11 (.D(d9_71__N_1675[11]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d9_i0_i12 (.D(d9_71__N_1675[12]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d9_i0_i13 (.D(d9_71__N_1675[13]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d9_i0_i14 (.D(d9_71__N_1675[14]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d9_i0_i15 (.D(d9_71__N_1675[15]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d9_i0_i16 (.D(d9_71__N_1675[16]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d9_i0_i17 (.D(d9_71__N_1675[17]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d9_i0_i18 (.D(d9_71__N_1675[18]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d9_i0_i19 (.D(d9_71__N_1675[19]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d9_i0_i20 (.D(d9_71__N_1675[20]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d9_i0_i21 (.D(d9_71__N_1675[21]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d9_i0_i22 (.D(d9_71__N_1675[22]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d9_i0_i23 (.D(d9_71__N_1675[23]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d9_i0_i24 (.D(d9_71__N_1675[24]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d9_i0_i25 (.D(d9_71__N_1675[25]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d9_i0_i26 (.D(d9_71__N_1675[26]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d9_i0_i27 (.D(d9_71__N_1675[27]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d9_i0_i28 (.D(d9_71__N_1675[28]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d9_i0_i29 (.D(d9_71__N_1675[29]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d9_i0_i30 (.D(d9_71__N_1675[30]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d9_i0_i31 (.D(d9_71__N_1675[31]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d9_i0_i32 (.D(d9_71__N_1675[32]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d9_i0_i33 (.D(d9_71__N_1675[33]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d9_i0_i34 (.D(d9_71__N_1675[34]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d9_i0_i35 (.D(d9_71__N_1675[35]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d9_i0_i36 (.D(d9_71__N_1675[36]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d9_i0_i37 (.D(d9_71__N_1675[37]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d9_i0_i38 (.D(d9_71__N_1675[38]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d9_i0_i39 (.D(d9_71__N_1675[39]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d9_i0_i40 (.D(d9_71__N_1675[40]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d9_i0_i41 (.D(d9_71__N_1675[41]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d9_i0_i42 (.D(d9_71__N_1675[42]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d9_i0_i43 (.D(d9_71__N_1675[43]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d9_i0_i44 (.D(d9_71__N_1675[44]), .SP(clk_80mhz_enable_599), 
            .CK(clk_80mhz), .Q(d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d9_i0_i45 (.D(d9_71__N_1675[45]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d9_i0_i46 (.D(d9_71__N_1675[46]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d9_i0_i47 (.D(d9_71__N_1675[47]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d9_i0_i48 (.D(d9_71__N_1675[48]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d9_i0_i49 (.D(d9_71__N_1675[49]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d9_i0_i50 (.D(d9_71__N_1675[50]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d9_i0_i51 (.D(d9_71__N_1675[51]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d9_i0_i52 (.D(d9_71__N_1675[52]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d9_i0_i53 (.D(d9_71__N_1675[53]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d9_i0_i54 (.D(d9_71__N_1675[54]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d9_i0_i55 (.D(d9_71__N_1675[55]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d9_i0_i56 (.D(d9_71__N_1675[56]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d9_i0_i57 (.D(d9_71__N_1675[57]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d9_i0_i58 (.D(d9_71__N_1675[58]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d9_i0_i59 (.D(d9_71__N_1675[59]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d9_i0_i60 (.D(d9_71__N_1675[60]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d9_i0_i61 (.D(d9_71__N_1675[61]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d9_i0_i62 (.D(d9_71__N_1675[62]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d9_i0_i63 (.D(d9_71__N_1675[63]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d9_i0_i64 (.D(d9_71__N_1675[64]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d9_i0_i65 (.D(d9_71__N_1675[65]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d9_i0_i66 (.D(d9_71__N_1675[66]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d9_i0_i67 (.D(d9_71__N_1675[67]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d9_i0_i68 (.D(d9_71__N_1675[68]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d9_i0_i69 (.D(d9_71__N_1675[69]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d9_i0_i70 (.D(d9_71__N_1675[70]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d9_i0_i71 (.D(d9_71__N_1675[71]), .SP(clk_80mhz_enable_649), 
            .CK(clk_80mhz), .Q(d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i1 (.D(d9[1]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i2 (.D(d9[2]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i3 (.D(d9[3]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i4 (.D(d9[4]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i5 (.D(d9[5]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i6 (.D(d9[6]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i7 (.D(d9[7]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i8 (.D(d9[8]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i9 (.D(d9[9]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i10 (.D(d9[10]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i11 (.D(d9[11]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i12 (.D(d9[12]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i13 (.D(d9[13]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i14 (.D(d9[14]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i15 (.D(d9[15]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i16 (.D(d9[16]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i17 (.D(d9[17]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i18 (.D(d9[18]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i19 (.D(d9[19]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i20 (.D(d9[20]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i21 (.D(d9[21]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i22 (.D(d9[22]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i23 (.D(d9[23]), .SP(clk_80mhz_enable_649), .CK(clk_80mhz), 
            .Q(d_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i24 (.D(d9[24]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i25 (.D(d9[25]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i26 (.D(d9[26]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i27 (.D(d9[27]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i28 (.D(d9[28]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i29 (.D(d9[29]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i30 (.D(d9[30]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i31 (.D(d9[31]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i32 (.D(d9[32]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i33 (.D(d9[33]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i34 (.D(d9[34]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i35 (.D(d9[35]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i36 (.D(d9[36]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i37 (.D(d9[37]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i38 (.D(d9[38]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i39 (.D(d9[39]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i40 (.D(d9[40]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i41 (.D(d9[41]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i42 (.D(d9[42]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i43 (.D(d9[43]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i44 (.D(d9[44]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i45 (.D(d9[45]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i46 (.D(d9[46]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i47 (.D(d9[47]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i48 (.D(d9[48]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i49 (.D(d9[49]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i50 (.D(d9[50]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i51 (.D(d9[51]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i52 (.D(d9[52]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i53 (.D(d9[53]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i54 (.D(d9[54]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i55 (.D(d9[55]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i56 (.D(d9[56]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i57 (.D(d9[57]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i58 (.D(d9[58]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i59 (.D(d9[59]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i60 (.D(d9[60]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i61 (.D(d9[61]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i62 (.D(d9[62]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i63 (.D(d9[63]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i64 (.D(d9[64]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i65 (.D(d9[65]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i66 (.D(d9[66]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i67 (.D(d9[67]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i68 (.D(d9[68]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i69 (.D(d9[69]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i70 (.D(d9[70]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX d_d9_i0_i71 (.D(d9[71]), .SP(clk_80mhz_enable_699), .CK(clk_80mhz), 
            .Q(d_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX d10__i2 (.D(d10_71__N_1747[57]), .SP(clk_80mhz_enable_699), 
            .CK(clk_80mhz), .Q(d10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i2.GSR = "ENABLED";
    FD1P3AX d10__i3 (.D(d10_71__N_1747[58]), .SP(clk_80mhz_enable_699), 
            .CK(clk_80mhz), .Q(d10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i3.GSR = "ENABLED";
    FD1P3AX d10__i4 (.D(d10_71__N_1747[59]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i4.GSR = "ENABLED";
    FD1P3AX d10__i5 (.D(d10_71__N_1747[60]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i5.GSR = "ENABLED";
    FD1P3AX d10__i6 (.D(d10_71__N_1747[61]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i6.GSR = "ENABLED";
    FD1P3AX d10__i7 (.D(d10_71__N_1747[62]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i7.GSR = "ENABLED";
    FD1P3AX d10__i8 (.D(d10_71__N_1747[63]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i8.GSR = "ENABLED";
    FD1P3AX d10__i9 (.D(d10_71__N_1747[64]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i9.GSR = "ENABLED";
    FD1P3AX d10__i10 (.D(d10_71__N_1747[65]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[65] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i10.GSR = "ENABLED";
    FD1P3AX d10__i11 (.D(d10_71__N_1747[66]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[66] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i11.GSR = "ENABLED";
    FD1P3AX d10__i12 (.D(d10_71__N_1747[67]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[67] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i12.GSR = "ENABLED";
    FD1P3AX d10__i13 (.D(d10_71__N_1747[68]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(\d10[68] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i13.GSR = "ENABLED";
    FD1P3AX d10__i14 (.D(d10_71__N_1747[69]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i14.GSR = "ENABLED";
    FD1P3AX d10__i15 (.D(d10_71__N_1747[70]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i15.GSR = "ENABLED";
    FD1P3AX d10__i16 (.D(d10_71__N_1747[71]), .SP(v_comb), .CK(clk_80mhz), 
            .Q(d10[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d10__i16.GSR = "ENABLED";
    FD1P3AX d_out_i0_i1 (.D(d_out_11__N_1819[1]), .SP(clk_80mhz_enable_700), 
            .CK(clk_80mhz), .Q(MultDataB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i1.GSR = "ENABLED";
    FD1P3AX d_out_i0_i2 (.D(\d_out_11__N_1819[2] ), .SP(clk_80mhz_enable_701), 
            .CK(clk_80mhz), .Q(MultDataB[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i2.GSR = "ENABLED";
    FD1P3AX d_out_i0_i3 (.D(\d_out_11__N_1819[3] ), .SP(clk_80mhz_enable_702), 
            .CK(clk_80mhz), .Q(MultDataB[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i3.GSR = "ENABLED";
    FD1P3AX d_out_i0_i4 (.D(\d_out_11__N_1819[4] ), .SP(clk_80mhz_enable_703), 
            .CK(clk_80mhz), .Q(MultDataB[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i4.GSR = "ENABLED";
    FD1P3AX d_out_i0_i5 (.D(\d_out_11__N_1819[5] ), .SP(clk_80mhz_enable_704), 
            .CK(clk_80mhz), .Q(MultDataB[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i5.GSR = "ENABLED";
    FD1P3AX d_out_i0_i6 (.D(\d_out_11__N_1819[6] ), .SP(clk_80mhz_enable_705), 
            .CK(clk_80mhz), .Q(MultDataB[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i6.GSR = "ENABLED";
    FD1P3AX d_out_i0_i7 (.D(\d_out_11__N_1819[7] ), .SP(clk_80mhz_enable_706), 
            .CK(clk_80mhz), .Q(MultDataB[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i7.GSR = "ENABLED";
    FD1P3AX d_out_i0_i8 (.D(\d_out_11__N_1819[8] ), .SP(clk_80mhz_enable_707), 
            .CK(clk_80mhz), .Q(MultDataB[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i8.GSR = "ENABLED";
    FD1P3AX d_out_i0_i9 (.D(d_out_11__N_1819[9]), .SP(clk_80mhz_enable_708), 
            .CK(clk_80mhz), .Q(MultDataB[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i9.GSR = "ENABLED";
    FD1P3AX d_out_i0_i10 (.D(d_out_11__N_1819[10]), .SP(clk_80mhz_enable_709), 
            .CK(clk_80mhz), .Q(MultDataB[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i10.GSR = "ENABLED";
    FD1P3AX d_out_i0_i11 (.D(d_out_11__N_1819[11]), .SP(clk_80mhz_enable_710), 
            .CK(clk_80mhz), .Q(MultDataB[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(85[12] 104[8])
    defparam d_out_i0_i11.GSR = "ENABLED";
    FD1S3AX d1_i1 (.D(d1_71__N_418[1]), .CK(clk_80mhz), .Q(d1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i1.GSR = "ENABLED";
    FD1S3AX d1_i2 (.D(d1_71__N_418[2]), .CK(clk_80mhz), .Q(d1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i2.GSR = "ENABLED";
    FD1S3AX d1_i3 (.D(d1_71__N_418[3]), .CK(clk_80mhz), .Q(d1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i3.GSR = "ENABLED";
    FD1S3AX d1_i4 (.D(d1_71__N_418[4]), .CK(clk_80mhz), .Q(d1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i4.GSR = "ENABLED";
    FD1S3AX d1_i5 (.D(d1_71__N_418[5]), .CK(clk_80mhz), .Q(d1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i5.GSR = "ENABLED";
    FD1S3AX d1_i6 (.D(d1_71__N_418[6]), .CK(clk_80mhz), .Q(d1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i6.GSR = "ENABLED";
    FD1S3AX d1_i7 (.D(d1_71__N_418[7]), .CK(clk_80mhz), .Q(d1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i7.GSR = "ENABLED";
    FD1S3AX d1_i8 (.D(d1_71__N_418[8]), .CK(clk_80mhz), .Q(d1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i8.GSR = "ENABLED";
    FD1S3AX d1_i9 (.D(d1_71__N_418[9]), .CK(clk_80mhz), .Q(d1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i9.GSR = "ENABLED";
    FD1S3AX d1_i10 (.D(d1_71__N_418[10]), .CK(clk_80mhz), .Q(d1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i10.GSR = "ENABLED";
    FD1S3AX d1_i11 (.D(d1_71__N_418[11]), .CK(clk_80mhz), .Q(d1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i11.GSR = "ENABLED";
    FD1S3AX d1_i12 (.D(d1_71__N_418[12]), .CK(clk_80mhz), .Q(d1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i12.GSR = "ENABLED";
    FD1S3AX d1_i13 (.D(d1_71__N_418[13]), .CK(clk_80mhz), .Q(d1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i13.GSR = "ENABLED";
    FD1S3AX d1_i14 (.D(d1_71__N_418[14]), .CK(clk_80mhz), .Q(d1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i14.GSR = "ENABLED";
    FD1S3AX d1_i15 (.D(d1_71__N_418[15]), .CK(clk_80mhz), .Q(d1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i15.GSR = "ENABLED";
    FD1S3AX d1_i16 (.D(d1_71__N_418[16]), .CK(clk_80mhz), .Q(d1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i16.GSR = "ENABLED";
    FD1S3AX d1_i17 (.D(d1_71__N_418[17]), .CK(clk_80mhz), .Q(d1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i17.GSR = "ENABLED";
    FD1S3AX d1_i18 (.D(d1_71__N_418[18]), .CK(clk_80mhz), .Q(d1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i18.GSR = "ENABLED";
    FD1S3AX d1_i19 (.D(d1_71__N_418[19]), .CK(clk_80mhz), .Q(d1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i19.GSR = "ENABLED";
    FD1S3AX d1_i20 (.D(d1_71__N_418[20]), .CK(clk_80mhz), .Q(d1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i20.GSR = "ENABLED";
    FD1S3AX d1_i21 (.D(d1_71__N_418[21]), .CK(clk_80mhz), .Q(d1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i21.GSR = "ENABLED";
    FD1S3AX d1_i22 (.D(d1_71__N_418[22]), .CK(clk_80mhz), .Q(d1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i22.GSR = "ENABLED";
    FD1S3AX d1_i23 (.D(d1_71__N_418[23]), .CK(clk_80mhz), .Q(d1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i23.GSR = "ENABLED";
    FD1S3AX d1_i24 (.D(d1_71__N_418[24]), .CK(clk_80mhz), .Q(d1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i24.GSR = "ENABLED";
    FD1S3AX d1_i25 (.D(d1_71__N_418[25]), .CK(clk_80mhz), .Q(d1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i25.GSR = "ENABLED";
    FD1S3AX d1_i26 (.D(d1_71__N_418[26]), .CK(clk_80mhz), .Q(d1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i26.GSR = "ENABLED";
    FD1S3AX d1_i27 (.D(d1_71__N_418[27]), .CK(clk_80mhz), .Q(d1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i27.GSR = "ENABLED";
    FD1S3AX d1_i28 (.D(d1_71__N_418[28]), .CK(clk_80mhz), .Q(d1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i28.GSR = "ENABLED";
    FD1S3AX d1_i29 (.D(d1_71__N_418[29]), .CK(clk_80mhz), .Q(d1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i29.GSR = "ENABLED";
    FD1S3AX d1_i30 (.D(d1_71__N_418[30]), .CK(clk_80mhz), .Q(d1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i30.GSR = "ENABLED";
    FD1S3AX d1_i31 (.D(d1_71__N_418[31]), .CK(clk_80mhz), .Q(d1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i31.GSR = "ENABLED";
    FD1S3AX d1_i32 (.D(d1_71__N_418[32]), .CK(clk_80mhz), .Q(d1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i32.GSR = "ENABLED";
    FD1S3AX d1_i33 (.D(d1_71__N_418[33]), .CK(clk_80mhz), .Q(d1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i33.GSR = "ENABLED";
    FD1S3AX d1_i34 (.D(d1_71__N_418[34]), .CK(clk_80mhz), .Q(d1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i34.GSR = "ENABLED";
    FD1S3AX d1_i35 (.D(d1_71__N_418[35]), .CK(clk_80mhz), .Q(d1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i35.GSR = "ENABLED";
    FD1S3AX d1_i36 (.D(d1_71__N_418[36]), .CK(clk_80mhz), .Q(d1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i36.GSR = "ENABLED";
    FD1S3AX d1_i37 (.D(d1_71__N_418[37]), .CK(clk_80mhz), .Q(d1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i37.GSR = "ENABLED";
    FD1S3AX d1_i38 (.D(d1_71__N_418[38]), .CK(clk_80mhz), .Q(d1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i38.GSR = "ENABLED";
    FD1S3AX d1_i39 (.D(d1_71__N_418[39]), .CK(clk_80mhz), .Q(d1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i39.GSR = "ENABLED";
    FD1S3AX d1_i40 (.D(d1_71__N_418[40]), .CK(clk_80mhz), .Q(d1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i40.GSR = "ENABLED";
    FD1S3AX d1_i41 (.D(d1_71__N_418[41]), .CK(clk_80mhz), .Q(d1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i41.GSR = "ENABLED";
    FD1S3AX d1_i42 (.D(d1_71__N_418[42]), .CK(clk_80mhz), .Q(d1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i42.GSR = "ENABLED";
    FD1S3AX d1_i43 (.D(d1_71__N_418[43]), .CK(clk_80mhz), .Q(d1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i43.GSR = "ENABLED";
    FD1S3AX d1_i44 (.D(d1_71__N_418[44]), .CK(clk_80mhz), .Q(d1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i44.GSR = "ENABLED";
    FD1S3AX d1_i45 (.D(d1_71__N_418[45]), .CK(clk_80mhz), .Q(d1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i45.GSR = "ENABLED";
    FD1S3AX d1_i46 (.D(d1_71__N_418[46]), .CK(clk_80mhz), .Q(d1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i46.GSR = "ENABLED";
    FD1S3AX d1_i47 (.D(d1_71__N_418[47]), .CK(clk_80mhz), .Q(d1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i47.GSR = "ENABLED";
    FD1S3AX d1_i48 (.D(d1_71__N_418[48]), .CK(clk_80mhz), .Q(d1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i48.GSR = "ENABLED";
    FD1S3AX d1_i49 (.D(d1_71__N_418[49]), .CK(clk_80mhz), .Q(d1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i49.GSR = "ENABLED";
    FD1S3AX d1_i50 (.D(d1_71__N_418[50]), .CK(clk_80mhz), .Q(d1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i50.GSR = "ENABLED";
    FD1S3AX d1_i51 (.D(d1_71__N_418[51]), .CK(clk_80mhz), .Q(d1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i51.GSR = "ENABLED";
    FD1S3AX d1_i52 (.D(d1_71__N_418[52]), .CK(clk_80mhz), .Q(d1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i52.GSR = "ENABLED";
    FD1S3AX d1_i53 (.D(d1_71__N_418[53]), .CK(clk_80mhz), .Q(d1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i53.GSR = "ENABLED";
    FD1S3AX d1_i54 (.D(d1_71__N_418[54]), .CK(clk_80mhz), .Q(d1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i54.GSR = "ENABLED";
    FD1S3AX d1_i55 (.D(d1_71__N_418[55]), .CK(clk_80mhz), .Q(d1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i55.GSR = "ENABLED";
    FD1S3AX d1_i56 (.D(d1_71__N_418[56]), .CK(clk_80mhz), .Q(d1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i56.GSR = "ENABLED";
    FD1S3AX d1_i57 (.D(d1_71__N_418[57]), .CK(clk_80mhz), .Q(d1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i57.GSR = "ENABLED";
    FD1S3AX d1_i58 (.D(d1_71__N_418[58]), .CK(clk_80mhz), .Q(d1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i58.GSR = "ENABLED";
    FD1S3AX d1_i59 (.D(d1_71__N_418[59]), .CK(clk_80mhz), .Q(d1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i59.GSR = "ENABLED";
    FD1S3AX d1_i60 (.D(d1_71__N_418[60]), .CK(clk_80mhz), .Q(d1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i60.GSR = "ENABLED";
    FD1S3AX d1_i61 (.D(d1_71__N_418[61]), .CK(clk_80mhz), .Q(d1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i61.GSR = "ENABLED";
    FD1S3AX d1_i62 (.D(d1_71__N_418[62]), .CK(clk_80mhz), .Q(d1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i62.GSR = "ENABLED";
    FD1S3AX d1_i63 (.D(d1_71__N_418[63]), .CK(clk_80mhz), .Q(d1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i63.GSR = "ENABLED";
    FD1S3AX d1_i64 (.D(d1_71__N_418[64]), .CK(clk_80mhz), .Q(d1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i64.GSR = "ENABLED";
    FD1S3AX d1_i65 (.D(d1_71__N_418[65]), .CK(clk_80mhz), .Q(d1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i65.GSR = "ENABLED";
    FD1S3AX d1_i66 (.D(d1_71__N_418[66]), .CK(clk_80mhz), .Q(d1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i66.GSR = "ENABLED";
    FD1S3AX d1_i67 (.D(d1_71__N_418[67]), .CK(clk_80mhz), .Q(d1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i67.GSR = "ENABLED";
    FD1S3AX d1_i68 (.D(d1_71__N_418[68]), .CK(clk_80mhz), .Q(d1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i68.GSR = "ENABLED";
    FD1S3AX d1_i69 (.D(d1_71__N_418[69]), .CK(clk_80mhz), .Q(d1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i69.GSR = "ENABLED";
    FD1S3AX d1_i70 (.D(d1_71__N_418[70]), .CK(clk_80mhz), .Q(d1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i70.GSR = "ENABLED";
    FD1S3AX d1_i71 (.D(d1_71__N_418[71]), .CK(clk_80mhz), .Q(d1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam d1_i71.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(n87_adj_126[2]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n87_adj_126[3]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n87_adj_126[4]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n87_adj_126[5]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n87_adj_126[6]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n87_adj_126[7]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n87_adj_126[8]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n87_adj_126[9]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n87_adj_126[10]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_15__N_1442[11]), .CK(clk_80mhz), .CD(d_clk_tmp_N_1831), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i11.GSR = "ENABLED";
    FD1S3IX count__i12 (.D(n87_adj_126[12]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i12.GSR = "ENABLED";
    FD1S3IX count__i13 (.D(n87_adj_126[13]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i13.GSR = "ENABLED";
    FD1S3IX count__i14 (.D(n87_adj_126[14]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i14.GSR = "ENABLED";
    FD1S3IX count__i15 (.D(n87_adj_126[15]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i15.GSR = "ENABLED";
    LUT4 shift_right_31_i62_rep_49_3_lut (.A(d10[61]), .B(d10[62]), .C(\CICGain[0] ), 
         .Z(n17636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i62_rep_49_3_lut.init = 16'hcaca;
    FD1S3IX count__i1 (.D(n87_adj_126[1]), .CK(clk_80mhz), .CD(n12697), 
            .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam count__i1.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i44_1_lut (.A(d_d8[43]), .Z(n30_adj_9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 i6329_4_lut_rep_195 (.A(n17054), .B(n17586), .C(n17562), .D(n17554), 
         .Z(clk_80mhz_enable_129)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i6329_4_lut_rep_195.init = 16'h4000;
    LUT4 shift_right_31_i63_3_lut (.A(d10[62]), .B(d10[63]), .C(\CICGain[0] ), 
         .Z(n63_adj_10)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i135_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65), .D(d10[63]), .Z(n135)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i134_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64), .D(d10[62]), .Z(n134)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i133_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_adj_10), .D(d10[61]), .Z(n133)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_25_inv_0_i66_1_lut (.A(d_d_tmp[65]), .Z(n8_adj_11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i132_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17636), .D(d10[60]), .Z(n132)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i136_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_adj_12), .D(d10[64]), .Z(n136)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i64_3_lut (.A(d10[63]), .B(d10[64]), .C(\CICGain[0] ), 
         .Z(n64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 sub_25_inv_0_i63_1_lut (.A(d_d_tmp[62]), .Z(n11_adj_13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i64_1_lut (.A(d_d_tmp[63]), .Z(n10_adj_14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i136_3_lut_4_lut_adj_26 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n66_adj_15), .D(\d10[64] ), .Z(n136_adj_16)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut_adj_26.init = 16'hf960;
    LUT4 shift_right_31_i135_3_lut_4_lut_adj_27 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n65_adj_17), .D(\d10[63] ), .Z(n135_adj_18)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut_adj_27.init = 16'hf960;
    LUT4 shift_right_31_i133_3_lut_4_lut_adj_28 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n63_adj_19), .D(\d10[61] ), .Z(n133_adj_20)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut_adj_28.init = 16'hf960;
    LUT4 sub_25_inv_0_i61_1_lut (.A(d_d_tmp[60]), .Z(n13_adj_21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i212_3_lut_4_lut_then_3_lut (.A(\CICGain[0] ), .B(\d10[68]_adj_22 ), 
         .C(\d10[69] ), .Z(n17984)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i212_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 shift_right_31_i212_3_lut_4_lut_else_3_lut (.A(\d10[71] ), .B(\CICGain[0] ), 
         .C(\d10[70] ), .Z(n17983)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i212_3_lut_4_lut_else_3_lut.init = 16'he2e2;
    LUT4 shift_right_31_i134_3_lut_4_lut_adj_29 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n64_adj_23), .D(\d10[62] ), .Z(n134_adj_24)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut_adj_29.init = 16'hf960;
    LUT4 sub_28_inv_0_i57_1_lut (.A(d_d8[56]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i58_1_lut (.A(d_d8[57]), .Z(n16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i55_1_lut (.A(d_d8[54]), .Z(n19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i56_1_lut (.A(d_d8[55]), .Z(n18_adj_25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i53_1_lut (.A(d_d8[52]), .Z(n21_adj_26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i54_1_lut (.A(d_d8[53]), .Z(n20_adj_27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i51_1_lut (.A(d_d8[50]), .Z(n23_adj_28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i52_1_lut (.A(d_d8[51]), .Z(n22_adj_29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 i2861_2_lut (.A(n31_c), .B(d_clk_tmp), .Z(n12681)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam i2861_2_lut.init = 16'h8888;
    LUT4 shift_right_31_i132_3_lut_4_lut_adj_30 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17610), .D(\d10[60] ), .Z(n132_adj_30)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut_adj_30.init = 16'hf960;
    LUT4 shift_right_31_i131_3_lut_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17630), .D(\d10[59] ), .Z(n131)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut.init = 16'hf960;
    LUT4 sub_25_inv_0_i62_1_lut (.A(d_d_tmp[61]), .Z(n12_adj_31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i71_1_lut (.A(d_d6[70]), .Z(n3_adj_32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i72_1_lut (.A(d_d6[71]), .Z(n2_adj_33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i64_1_lut (.A(d_d7[63]), .Z(n10_adj_34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i61_1_lut (.A(d_d7[60]), .Z(n13_adj_35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i62_1_lut (.A(d_d7[61]), .Z(n12_adj_36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i59_1_lut (.A(d_d7[58]), .Z(n15_adj_37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i60_1_lut (.A(d_d7[59]), .Z(n14_adj_38)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i57_1_lut (.A(d_d7[56]), .Z(n17_adj_39)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i58_1_lut (.A(d_d7[57]), .Z(n16_adj_40)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i55_1_lut (.A(d_d7[54]), .Z(n19_adj_41)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i131_3_lut_4_lut_adj_31 (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(n17655), .D(d10[59]), .Z(n131_adj_42)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut_adj_31.init = 16'hf960;
    LUT4 i11_3_lut_4_lut_then_3_lut (.A(\CICGain[0] ), .B(\d10[67]_adj_43 ), 
         .C(\d10[68]_adj_22 ), .Z(n17987)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam i11_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 sub_27_inv_0_i56_1_lut (.A(d_d7[55]), .Z(n18_adj_44)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i53_1_lut (.A(d_d7[52]), .Z(n21_adj_45)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i54_1_lut (.A(d_d7[53]), .Z(n20_adj_46)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i51_1_lut (.A(d_d7[50]), .Z(n23_adj_47)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i52_1_lut (.A(d_d7[51]), .Z(n22_adj_48)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i65_3_lut (.A(d10[64]), .B(\d10[65] ), .C(\CICGain[0] ), 
         .Z(n65)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    LUT4 i11_3_lut_4_lut_else_3_lut (.A(\d10[70] ), .B(\CICGain[0] ), .C(\d10[69] ), 
         .Z(n17986)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam i11_3_lut_4_lut_else_3_lut.init = 16'he2e2;
    LUT4 sub_28_inv_0_i49_1_lut (.A(d_d8[48]), .Z(n25_adj_49)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i50_1_lut (.A(d_d8[49]), .Z(n24_adj_50)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i49_1_lut (.A(d_d7[48]), .Z(n25_adj_51)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i50_1_lut (.A(d_d7[49]), .Z(n24_adj_52)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i47_1_lut (.A(d_d7[46]), .Z(n27_adj_53)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i48_1_lut (.A(d_d7[47]), .Z(n26_adj_54)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i45_1_lut (.A(d_d7[44]), .Z(n29_adj_55)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i46_1_lut (.A(d_d7[45]), .Z(n28_adj_56)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i43_1_lut (.A(d_d7[42]), .Z(n31_adj_57)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i44_1_lut (.A(d_d7[43]), .Z(n30_adj_58)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i41_1_lut (.A(d_d7[40]), .Z(n33_adj_59)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i42_1_lut (.A(d_d7[41]), .Z(n32_adj_60)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i47_1_lut (.A(d_d8[46]), .Z(n27_adj_61)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i47_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_182 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_11)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_182.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i39_1_lut (.A(d_d7[38]), .Z(n35_adj_62)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i40_1_lut (.A(d_d7[39]), .Z(n34_adj_63)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i37_1_lut (.A(d_d7[36]), .Z(n37_adj_64)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i38_1_lut (.A(d_d7[37]), .Z(n36_adj_65)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i212_3_lut_4_lut_then_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(\d10[68] ), .D(n17628), .Z(n17990)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((D)+!B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i212_3_lut_4_lut_then_4_lut.init = 16'hf791;
    LUT4 sub_25_inv_0_i59_1_lut (.A(d_d_tmp[58]), .Z(n15_adj_66)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i59_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_185 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_702)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_185.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_187 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_704)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_187.GSR = "ENABLED";
    LUT4 shift_right_31_i212_3_lut_4_lut_else_4_lut (.A(\CICGain[1] ), .B(\CICGain[0] ), 
         .C(\d10[68] ), .D(n17628), .Z(n17989)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (D))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i212_3_lut_4_lut_else_4_lut.init = 16'he680;
    LUT4 shift_right_31_i66_3_lut (.A(\d10[65] ), .B(\d10[66] ), .C(\CICGain[0] ), 
         .Z(n66_adj_12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 i11_3_lut_4_lut_then_3_lut_adj_32 (.A(\CICGain[0] ), .B(\d10[67] ), 
         .C(\d10[68] ), .Z(n17993)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam i11_3_lut_4_lut_then_3_lut_adj_32.init = 16'hd8d8;
    LUT4 i11_3_lut_4_lut_else_3_lut_adj_33 (.A(d10[70]), .B(\CICGain[0] ), 
         .C(d10[69]), .Z(n17992)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam i11_3_lut_4_lut_else_3_lut_adj_33.init = 16'he2e2;
    LUT4 sub_25_inv_0_i60_1_lut (.A(d_d_tmp[59]), .Z(n14_adj_67)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i57_1_lut (.A(d_d_tmp[56]), .Z(n17_adj_68)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i58_1_lut (.A(d_d_tmp[57]), .Z(n16_adj_69)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i58_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_207 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_599)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_207.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i69_1_lut (.A(d_d6[68]), .Z(n5_adj_70)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i70_1_lut (.A(d_d6[69]), .Z(n4_adj_71)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i41_1_lut (.A(d_d8[40]), .Z(n33_adj_72)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i67_1_lut (.A(d_d6[66]), .Z(n7_adj_73)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i42_1_lut (.A(d_d8[41]), .Z(n32_adj_74)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i39_1_lut (.A(d_d8[38]), .Z(n35_adj_75)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i40_1_lut (.A(d_d8[39]), .Z(n34_adj_76)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i68_1_lut (.A(d_d6[67]), .Z(n6_adj_77)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i68_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_206 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_549)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_206.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i65_1_lut (.A(d_d6[64]), .Z(n9_adj_78)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 i1_3_lut (.A(count[8]), .B(count[1]), .C(count[9]), .Z(n17459)) /* synthesis lut_function=(A+(B+(C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_34 (.A(count[10]), .B(count[6]), .C(count[7]), .D(count[5]), 
         .Z(n17463)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i1_4_lut_adj_34.init = 16'hfffe;
    LUT4 i1_4_lut_adj_35 (.A(count[2]), .B(count[4]), .C(count[0]), .D(count[3]), 
         .Z(n17461)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(69[13:41])
    defparam i1_4_lut_adj_35.init = 16'hfffe;
    LUT4 sub_26_inv_0_i66_1_lut (.A(d_d6[65]), .Z(n8_adj_79)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i63_1_lut (.A(d_d6[62]), .Z(n11_adj_80)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i63_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_205 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_499)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_205.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i37_1_lut (.A(d_d8[36]), .Z(n37_adj_81)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i64_1_lut (.A(d_d6[63]), .Z(n10_adj_82)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i38_1_lut (.A(d_d8[37]), .Z(n36_adj_83)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i61_1_lut (.A(d_d6[60]), .Z(n13_adj_84)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i71_1_lut (.A(d_d7[70]), .Z(n3_adj_85)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i72_1_lut (.A(d_d7[71]), .Z(n2_adj_86)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i69_1_lut (.A(d_d7[68]), .Z(n5_adj_87)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i62_1_lut (.A(d_d6[61]), .Z(n12_adj_88)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i62_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_186 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_703)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_186.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i70_1_lut (.A(d_d7[69]), .Z(n4_adj_89)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i67_1_lut (.A(d_d7[66]), .Z(n7_adj_90)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i59_1_lut (.A(d_d6[58]), .Z(n15_adj_91)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i61_rep_68_3_lut (.A(d10[60]), .B(d10[61]), .C(\CICGain[0] ), 
         .Z(n17655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i61_rep_68_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i60_1_lut (.A(d_d6[59]), .Z(n14_adj_92)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i68_1_lut (.A(d_d7[67]), .Z(n6_adj_93)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i70_rep_41_3_lut (.A(d10[69]), .B(d10[70]), .C(\CICGain[0] ), 
         .Z(n17628)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(102[25:52])
    defparam shift_right_31_i70_rep_41_3_lut.init = 16'hcaca;
    LUT4 sub_26_inv_0_i57_1_lut (.A(d_d6[56]), .Z(n17_adj_94)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i55_1_lut (.A(d_d_tmp[54]), .Z(n19_adj_95)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i56_1_lut (.A(d_d_tmp[55]), .Z(n18_adj_96)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i65_1_lut (.A(d_d7[64]), .Z(n9_adj_97)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(95[25:34])
    defparam sub_27_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i58_1_lut (.A(d_d6[57]), .Z(n16_adj_98)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i58_1_lut.init = 16'h5555;
    PFUMX i6441 (.BLUT(n17992), .ALUT(n17993), .C0(\CICGain[1] ), .Z(d_out_11__N_1819[10]));
    PFUMX i6439 (.BLUT(n17989), .ALUT(n17990), .C0(d10[71]), .Z(d_out_11__N_1819[11]));
    PFUMX i6437 (.BLUT(n17986), .ALUT(n17987), .C0(\CICGain[1] ), .Z(\d_out_11__N_1819[10] ));
    LUT4 sub_26_inv_0_i55_1_lut (.A(d_d6[54]), .Z(n19_adj_99)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(93[25:34])
    defparam sub_26_inv_0_i55_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_204 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_449)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_204.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_203 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_399)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_203.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i53_1_lut (.A(d_d_tmp[52]), .Z(n21_adj_100)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i54_1_lut (.A(d_d_tmp[53]), .Z(n20_adj_101)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i54_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_202 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_349)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_202.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_201 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_299)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_201.GSR = "ENABLED";
    PFUMX i6435 (.BLUT(n17983), .ALUT(n17984), .C0(\CICGain[1] ), .Z(\d_out_11__N_1819[11] ));
    FD1S3AX v_comb_66_rep_188 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_705)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_188.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_200 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_249)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_200.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_199 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_199)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_199.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_198 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_149)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_198.GSR = "ENABLED";
    LUT4 i6332_2_lut (.A(n31_c), .B(n18089), .Z(n12697)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam i6332_2_lut.init = 16'hdddd;
    LUT4 sub_25_inv_0_i51_1_lut (.A(d_d_tmp[50]), .Z(n23_adj_102)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i51_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_197 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_65)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_197.GSR = "ENABLED";
    LUT4 i3168_2_lut (.A(n87_adj_126[11]), .B(n31_c), .Z(count_15__N_1442[11])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(78[18] 81[12])
    defparam i3168_2_lut.init = 16'hbbbb;
    LUT4 sub_25_inv_0_i52_1_lut (.A(d_d_tmp[51]), .Z(n22_adj_103)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 i3117_2_lut (.A(n87_adj_126[0]), .B(n31_c), .Z(count_15__N_1442[0])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(78[18] 81[12])
    defparam i3117_2_lut.init = 16'hbbbb;
    PFUMX i6427 (.BLUT(n17971), .ALUT(n17972), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[9]));
    FD1S3AX v_comb_66_rep_193 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_710)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_193.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i49_1_lut (.A(d_d_tmp[48]), .Z(n25_adj_104)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i49_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_192 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_709)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_192.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_191 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_708)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_191.GSR = "ENABLED";
    FD1S3AX v_comb_66_rep_184 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_701)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_184.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i50_1_lut (.A(d_d_tmp[49]), .Z(n24_adj_105)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i50_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_183 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_700)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_183.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i47_1_lut (.A(d_d_tmp[46]), .Z(n27_adj_106)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i48_1_lut (.A(d_d_tmp[47]), .Z(n26_adj_107)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i48_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_190 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_707)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_190.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i45_1_lut (.A(d_d_tmp[44]), .Z(n29_adj_108)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i46_1_lut (.A(d_d_tmp[45]), .Z(n28_adj_109)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i43_1_lut (.A(d_d_tmp[42]), .Z(n31_adj_110)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i44_1_lut (.A(d_d_tmp[43]), .Z(n30_adj_111)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i41_1_lut (.A(d_d_tmp[40]), .Z(n33_adj_112)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i42_1_lut (.A(d_d_tmp[41]), .Z(n32_adj_113)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i39_1_lut (.A(d_d_tmp[38]), .Z(n35_adj_114)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i40_1_lut (.A(d_d_tmp[39]), .Z(n34_adj_115)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i37_1_lut (.A(d_d_tmp[36]), .Z(n37_adj_116)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i38_1_lut (.A(d_d_tmp[37]), .Z(n36_adj_117)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(91[25:40])
    defparam sub_25_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i71_1_lut (.A(d_d8[70]), .Z(n3_adj_118)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i71_1_lut.init = 16'h5555;
    PFUMX i6421 (.BLUT(n17962), .ALUT(n17963), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[1]));
    LUT4 sub_28_inv_0_i72_1_lut (.A(d_d8[71]), .Z(n2_adj_119)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i69_1_lut (.A(d_d8[68]), .Z(n5_adj_120)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i70_1_lut (.A(d_d8[69]), .Z(n4_adj_121)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i67_1_lut (.A(d_d8[66]), .Z(n7_adj_122)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i68_1_lut (.A(d_d8[67]), .Z(n6_adj_123)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i65_1_lut (.A(d_d8[64]), .Z(n9_adj_124)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i65_1_lut.init = 16'h5555;
    FD1S3AX v_comb_66_rep_209 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_699)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_209.GSR = "ENABLED";
    PFUMX i6417 (.BLUT(n17956), .ALUT(n17957), .C0(\CICGain[0] ), .Z(d_out_11__N_1819[0]));
    FD1S3AX v_comb_66_rep_208 (.D(clk_80mhz_enable_129), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_649)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=5, LSE_LLINE=136, LSE_RLINE=142 */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(61[12] 82[8])
    defparam v_comb_66_rep_208.GSR = "ENABLED";
    LUT4 sub_28_inv_0_i66_1_lut (.A(d_d8[65]), .Z(n8_adj_125)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1bitSDRLattice/First_Implementation/source/CIC.v(97[25:34])
    defparam sub_28_inv_0_i66_1_lut.init = 16'h5555;
    
endmodule
