// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.13.0.56.2
// Netlist written on Wed Aug  7 15:42:12 2024
//
// Verilog Description of module top
//

module top (clk_25mhz, rx_serial, rf_in, diff_out, pwm_out, pwm_out_p1, 
            pwm_out_p2, pwm_out_p3, pwm_out_p4, pwm_out_n1, pwm_out_n2, 
            pwm_out_n3, pwm_out_n4, led) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(38[8:11])
    input clk_25mhz;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(39[16:25])
    input rx_serial;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(40[16:25])
    input rf_in;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(41[16:21])
    output diff_out;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(43[23:31])
    output pwm_out;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(44[23:30])
    output pwm_out_p1;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(45[23:33])
    output pwm_out_p2;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(46[23:33])
    output pwm_out_p3;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(47[23:33])
    output pwm_out_p4;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(48[23:33])
    output pwm_out_n1;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(49[23:33])
    output pwm_out_n2;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(50[23:33])
    output pwm_out_n3;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(51[23:33])
    output pwm_out_n4;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(52[23:33])
    output [7:0]led;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(53[23:26])
    
    wire clk_25mhz_c /* synthesis is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(39[16:25])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(64[10:19])
    wire cic_sine_clk /* synthesis SET_AS_NETWORK=cic_sine_clk, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(86[10:22])
    
    wire GND_net, VCC_net, rx_serial_c, rf_in_c, diff_out_c, pwm_out_p4_c, 
        pwm_out_n4_c, led_c_7, led_c_6, led_c_5, led_c_4, led_c_3, 
        led_c_2, led_c_1, led_c_0;
    wire [63:0]phase_inc_gen;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(69[23:36])
    wire [63:0]phase_inc_gen1;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(70[23:37])
    wire [63:0]phase_acc;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(73[17:26])
    wire [12:0]lo_sinewave;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(76[24:35])
    wire [12:0]lo_cosinewave;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(77[24:37])
    wire [11:0]mix_sinewave;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(80[24:36])
    wire [11:0]mix_cosinewave;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(81[24:38])
    
    wire n15536;
    wire [7:0]cic_gain;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(84[15:23])
    wire [11:0]cic_cosine_out;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(87[24:38])
    wire [11:0]amdemod_out;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(91[24:35])
    
    wire n15535, n16, rx_data_valid, rx_data_valid1;
    wire [7:0]rx_byte1;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(97[16:24])
    
    wire n27, n37, n36, n35, n34, n33, n32, n31, n30, n29, 
        n28, n27_adj_2946, n26, n25, n24, n23, n22, n21, n20, 
        n19, n18, n17, n16_adj_2947, n15, n14, n13, n12, n11, 
        n10, n9, n8, n7, n6, n5, n4, n3, n2, n2594, n4_adj_2948, 
        clk_80mhz_enable_1444, n2580, n2579, n15390, n15380, n15389, 
        n15388, clk_80mhz_enable_1507, n2559, n15386, n15385, n15384, 
        n15383, n15382, n15381, n2545, n16348, n15_adj_2949, n14_adj_2950, 
        n13_adj_2951, n12_adj_2952, n11_adj_2953, n10_adj_2954, n9_adj_2955, 
        n8_adj_2956, n7_adj_2957, n6_adj_2958, n5_adj_2959, n4_adj_2960, 
        n12278, n15534, n15533, n3_adj_2961, n2_adj_2962, n15532, 
        n15531;
    wire [63:0]phase_accum;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(26[28:39])
    
    wire n37_adj_2963, n36_adj_2964, n35_adj_2965, n34_adj_2966, n33_adj_2967, 
        n32_adj_2968, n31_adj_2969, n30_adj_2970, n29_adj_2971, n28_adj_2972, 
        n26_adj_2973, n15529, n25_adj_2974, n15742, n15741, n15740, 
        n15739, n15738, n15737, n2102, n15735, n15734, n15733, 
        n15732, n2097, n15731, n15730, n2094, n15729, n15728, 
        n15727, n15726, n15725, n15724, n15723, n15722, n15721, 
        n15720, n15719, n15718, n15714, n15713, n15712, n15711, 
        n15710, n15709, n15708, n15706, n15705, n15704, n15703, 
        n2065, n15702, n15701, n15700, n15699, n71, n68, n65, 
        n62, n59, n56, n53, n2060;
    wire [11:0]sinewave_out_11__N_236;
    wire [11:0]cosinewave_out_11__N_250;
    wire [71:0]integrator_tmp;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(56[41:55])
    wire [71:0]integrator_d_tmp;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(56[57:73])
    wire [71:0]integrator1;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(57[41:52])
    wire [71:0]integrator2;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(57[54:65])
    wire [71:0]integrator3;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(57[67:78])
    wire [71:0]integrator4;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(57[80:91])
    wire [71:0]integrator5;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(57[93:104])
    wire [71:0]comb6;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[41:46])
    wire [71:0]comb_d6;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[48:55])
    wire [71:0]comb7;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[57:62])
    wire [71:0]comb_d7;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[64:71])
    wire [71:0]comb8;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[73:78])
    wire [71:0]comb_d8;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[80:87])
    wire [71:0]comb9;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[89:94])
    wire [71:0]comb_d9;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[96:103])
    
    wire n15528;
    wire [11:0]count;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(60[32:37])
    wire [71:0]integrator1_71__N_418;
    wire [71:0]integrator2_71__N_490;
    wire [71:0]integrator3_71__N_562;
    wire [71:0]integrator4_71__N_634;
    wire [71:0]integrator5_71__N_706;
    
    wire n15379, n15378, n15698, n15697, n15696, n15695, n15694, 
        n15693, n15692, n15691, n15690, n15689;
    wire [71:0]comb6_71__N_1451;
    wire [71:0]comb7_71__N_1523;
    wire [71:0]comb8_71__N_1595;
    wire [71:0]comb9_71__N_1667;
    
    wire n15527, n15526, n15525, n15688;
    wire [71:0]integrator_tmp_adj_6018;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(56[41:55])
    wire [71:0]integrator_d_tmp_adj_6019;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(56[57:73])
    wire [71:0]integrator1_adj_6020;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(57[41:52])
    wire [71:0]integrator2_adj_6021;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(57[54:65])
    wire [71:0]integrator3_adj_6022;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(57[67:78])
    wire [71:0]integrator4_adj_6023;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(57[80:91])
    wire [71:0]integrator5_adj_6024;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(57[93:104])
    wire [71:0]comb6_adj_6025;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[41:46])
    wire [71:0]comb_d6_adj_6026;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[48:55])
    wire [71:0]comb7_adj_6027;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[57:62])
    wire [71:0]comb_d7_adj_6028;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[64:71])
    wire [71:0]comb8_adj_6029;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[73:78])
    wire [71:0]comb_d8_adj_6030;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[80:87])
    wire [71:0]comb9_adj_6031;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[89:94])
    wire [71:0]comb_d9_adj_6032;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[96:103])
    wire [71:0]comb10_adj_6033;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[105:111])
    
    wire n15524;
    wire [11:0]count_adj_6035;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(60[32:37])
    wire [71:0]integrator1_71__N_418_adj_6036;
    wire [71:0]integrator2_71__N_490_adj_6037;
    wire [71:0]integrator3_71__N_562_adj_6038;
    wire [71:0]integrator4_71__N_634_adj_6039;
    wire [71:0]integrator5_71__N_706_adj_6040;
    
    wire n15687, n15686, n15685, n15684, n15683, n15682, n15681, 
        n15680, n15679, n15678;
    wire [71:0]comb6_71__N_1451_adj_6052;
    wire [71:0]comb7_71__N_1523_adj_6053;
    wire [71:0]comb8_71__N_1595_adj_6054;
    wire [71:0]comb9_71__N_1667_adj_6055;
    
    wire n15523, n15377, n15376, n15375, n15374, n15373, n15372, 
        n15371, n15370, n15369, n15367, n15366, n15365, n15364, 
        n15363, n15362, n15677, n15676;
    wire [71:0]data_out_11__N_1811_adj_6058;
    
    wire n15522, n15521, n15520, n16388, n15519, n15518, n15517, 
        n15516, n15515, n15514, n15513, n15512, n15508, n15361, 
        n15360;
    wire [25:0]square_sum;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(31[38:48])
    wire [11:0]mult_i_b;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(34[38:46])
    wire [23:0]mult_result_i;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(35[38:51])
    
    wire n50, n47, n44, n41, n38, n32_adj_4715, n24_adj_4716;
    wire [13:0]amdemod_d_11__N_1830;
    
    wire amdemod_d_11__N_2005, amdemod_d_11__N_2008, amdemod_d_11__N_2011, 
        amdemod_d_11__N_2014, amdemod_d_11__N_2017, amdemod_d_11__N_2020, 
        amdemod_d_11__N_2023, amdemod_d_11__N_2026, n15359;
    wire [13:0]amdemod_d_11__N_1841;
    
    wire n15358;
    wire [13:0]amdemod_d_11__N_1840;
    
    wire amdemod_d_11__N_2065, amdemod_d_11__N_2068, amdemod_d_11__N_2071, 
        amdemod_d_11__N_2074, amdemod_d_11__N_2077, amdemod_d_11__N_2080, 
        amdemod_d_11__N_2083, amdemod_d_11__N_2086, amdemod_d_11__N_2089, 
        amdemod_d_11__N_2092, amdemod_d_11__N_2095, amdemod_d_11__N_2098;
    wire [13:0]amdemod_d_11__N_1851;
    wire [13:0]amdemod_d_11__N_1850;
    
    wire amdemod_d_11__N_2137, amdemod_d_11__N_2140, amdemod_d_11__N_2143, 
        amdemod_d_11__N_2146, amdemod_d_11__N_2149, amdemod_d_11__N_2152, 
        amdemod_d_11__N_2155, amdemod_d_11__N_2158, amdemod_d_11__N_2161, 
        amdemod_d_11__N_2164, amdemod_d_11__N_2167, amdemod_d_11__N_2170;
    wire [13:0]amdemod_d_11__N_1861;
    wire [13:0]amdemod_d_11__N_1860;
    
    wire clk_80mhz_enable_1497, amdemod_d_11__N_2209, amdemod_d_11__N_2212, 
        amdemod_d_11__N_2215, amdemod_d_11__N_2218, amdemod_d_11__N_2221, 
        amdemod_d_11__N_2224, amdemod_d_11__N_2227, amdemod_d_11__N_2230, 
        amdemod_d_11__N_2233, amdemod_d_11__N_2236, amdemod_d_11__N_2239, 
        amdemod_d_11__N_2242;
    wire [13:0]amdemod_d_11__N_1871;
    wire [13:0]amdemod_d_11__N_1870;
    
    wire n17335, amdemod_d_11__N_1874, amdemod_d_11__N_2281, amdemod_d_11__N_2284, 
        amdemod_d_11__N_2287, amdemod_d_11__N_2290, amdemod_d_11__N_2293, 
        amdemod_d_11__N_2296, amdemod_d_11__N_2299, amdemod_d_11__N_2302, 
        amdemod_d_11__N_2305, amdemod_d_11__N_2308, amdemod_d_11__N_2311, 
        amdemod_d_11__N_2314;
    wire [13:0]amdemod_d_11__N_1881;
    wire [13:0]amdemod_d_11__N_1880;
    wire [9:0]count_adj_6105;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(40[27:32])
    wire [11:0]data_in_reg;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(41[27:38])
    
    wire n15507;
    wire [31:0]data_in_reg_11__N_2339;
    
    wire n15357, n15675, n15674, n15673, n23_adj_4727, n15506, n15505, 
        n15504, n15503, n15672, n17134, n15502, n15500, n11789, 
        n15499, n15498, n15497, n15496, n15495, n15494, n15671, 
        n15670, n15669, n2054, n15668, n15667, n15666, n15665, 
        n15664, n15663, n15662, n15661, n15660, n15659, n15658, 
        n15657, n15656, n15655, n15654, n15653, n15652, n15651, 
        n15650, n15649, n15648, n15647, n15646, n15645, n15644, 
        n15643, n15642, n15641, n17152, n17133, n15493, n15640, 
        n15639, n15638, n15637, n15636, n15635, n15634, n15633, 
        n15632, n15356, n15355, n15354, n15492, n15491, n15490, 
        n15489, n15488, n15487, n15486, n15631, n15630, n15629, 
        n15628, n15353, n15352, n15351, n15350, n15349, n15348, 
        n15347, n15346, n15345, n15344, n15343, n15342, n15341, 
        n15340, n15339, n15338, n15337, n15336, n15335, n17132, 
        n17131, n17130, n17150, n17149, n17148, n22_adj_4728, n15485, 
        n15484, n15483, n15482, n11_adj_4729, n71_adj_4730, n15481, 
        n15480, n15479, n68_adj_4731, n65_adj_4732, n62_adj_4733, 
        n59_adj_4734, n56_adj_4735, n53_adj_4736, n50_adj_4737, n47_adj_4738, 
        n44_adj_4739, n41_adj_4740, n38_adj_4741, n32_adj_4742, n15478, 
        n15477, n15476, n21_adj_4743, n17175, n17176, n2040, n2039, 
        n2038, n2037, n2036, n2035, n2034, n2032, n2031, n2030, 
        n2029, n2028, n2027, n2026, n2024, n2021, n2020, n2019, 
        n2018, n2017, n20_adj_4744, n15627, n15626, n15625, n15624, 
        n15623, n2244, n15475, n15622, n2237, n15621, n15619, 
        n2230, n15618, n2226, n11624, n15617, n11622, n15616, 
        n11620, n2214, n15474, n17129, n17128, n62_adj_4745, n63, 
        n64, n65_adj_4746, n66, n17147, n17146, n17144, n17288, 
        n80, n79, n78, n11179, n77, n76, n75, n74, n73, n72, 
        n13_adj_4747, n15473, n15472, n15471, n1827, n19_adj_4748, 
        n15470, n71_adj_4749, n70, n69, n68_adj_4750, n15468, n15467, 
        n15466, n73_adj_4751, n67, n66_adj_4752, n65_adj_4753, n64_adj_4754, 
        n63_adj_4755, n62_adj_4756, n2016, n2015, n2014, n2013, 
        n2012, n2011, n2010, n2009, n2008, n2007, n2006, n2005, 
        n2002, n2001, n2000, n1999, n1998, n1997, n1996, n1995, 
        n1994, n1993, n1991, n1990, n1989, n1988, n1986, n1985, 
        n1984, n6_adj_4757, n61, n60, n59_adj_4758, n58, n57, 
        n70_adj_4759, n15615, n11618, n15614, n15613, n11616, n15612, 
        n2193, n11614, n15611, n11612, n15610, n2187, n15609, 
        n11608, n15608, n15607, n15606, n67_adj_4760, n18_adj_4761, 
        n15605, n15604, n15603, n15465, n15464, n15463, n15462, 
        n15461, n15460, n15459, n15458, n15457, n15456, n15455, 
        n64_adj_4762, n15454, n15453, n15452, n15451, n15450, n15449, 
        n15867, n17_adj_4763, n61_adj_4764, n58_adj_4765, n15602, 
        n2_adj_4766, n3_adj_4767, n4_adj_4768, n5_adj_4769, n6_adj_4770, 
        n7_adj_4771, n8_adj_4772, n9_adj_4773, n10_adj_4774, n11_adj_4775, 
        n12_adj_4776, n13_adj_4777, n14_adj_4778, n15_adj_4779, n16_adj_4780, 
        n17_adj_4781, n18_adj_4782, n19_adj_4783, n20_adj_4784, n21_adj_4785, 
        n22_adj_4786, n23_adj_4787, n24_adj_4788, n25_adj_4789, n26_adj_4790, 
        n27_adj_4791, n28_adj_4792, n29_adj_4793, n30_adj_4794, n31_adj_4795, 
        n32_adj_4796, n33_adj_4797, n34_adj_4798, n35_adj_4799, n36_adj_4800, 
        n37_adj_4801, n2_adj_4802, n3_adj_4803, n4_adj_4804, n5_adj_4805, 
        n6_adj_4806, n7_adj_4807, n8_adj_4808, n9_adj_4809, n10_adj_4810, 
        n11_adj_4811, n12_adj_4812, n13_adj_4813, n14_adj_4814, n15_adj_4815, 
        n16_adj_4816, n17_adj_4817, n18_adj_4818, n19_adj_4819, n20_adj_4820, 
        n21_adj_4821, n22_adj_4822, n23_adj_4823, n24_adj_4824, n25_adj_4825, 
        n26_adj_4826, n27_adj_4827, n28_adj_4828, n29_adj_4829, n30_adj_4830, 
        n31_adj_4831, n32_adj_4832, n33_adj_4833, n34_adj_4834, n35_adj_4835, 
        n36_adj_4836, n37_adj_4837, n2_adj_4838, n3_adj_4839, n4_adj_4840, 
        n5_adj_4841, n6_adj_4842, n7_adj_4843, n8_adj_4844, n9_adj_4845, 
        n10_adj_4846, n11_adj_4847, n12_adj_4848, n13_adj_4849, n14_adj_4850, 
        n15_adj_4851, n16_adj_4852, n17_adj_4853, n18_adj_4854, n19_adj_4855, 
        n20_adj_4856, n21_adj_4857, n22_adj_4858, n23_adj_4859, n24_adj_4860, 
        n25_adj_4861, n26_adj_4862, n27_adj_4863, n28_adj_4864, n29_adj_4865, 
        n30_adj_4866, n31_adj_4867, n32_adj_4868, n33_adj_4869, n34_adj_4870, 
        n35_adj_4871, n36_adj_4872, n37_adj_4873, n2_adj_4874, n3_adj_4875, 
        n4_adj_4876, n5_adj_4877, n6_adj_4878, n7_adj_4879, n8_adj_4880, 
        n9_adj_4881, n10_adj_4882, n11_adj_4883, n12_adj_4884, n13_adj_4885, 
        n14_adj_4886, n15_adj_4887, n16_adj_4888, n17_adj_4889, n18_adj_4890, 
        n19_adj_4891, n20_adj_4892, n21_adj_4893, n22_adj_4894, n23_adj_4895, 
        n24_adj_4896, n25_adj_4897, n26_adj_4898, n27_adj_4899, n28_adj_4900, 
        n29_adj_4901, n30_adj_4902, n31_adj_4903, n32_adj_4904, n33_adj_4905, 
        n34_adj_4906, n35_adj_4907, n36_adj_4908, n37_adj_4909, n2_adj_4910, 
        n3_adj_4911, n4_adj_4912, n5_adj_4913, n6_adj_4914, n7_adj_4915, 
        n8_adj_4916, n9_adj_4917, n10_adj_4918, n11_adj_4919, n12_adj_4920, 
        n13_adj_4921, n14_adj_4922, n15_adj_4923, n16_adj_4924, n17_adj_4925, 
        n18_adj_4926, n19_adj_4927, n20_adj_4928, n21_adj_4929, n22_adj_4930, 
        n23_adj_4931, n24_adj_4932, n25_adj_4933, n26_adj_4934, n27_adj_4935, 
        n28_adj_4936, n29_adj_4937, n30_adj_4938, n31_adj_4939, n32_adj_4940, 
        n33_adj_4941, n34_adj_4942, n35_adj_4943, n36_adj_4944, n37_adj_4945, 
        n15334, n2_adj_4946, n3_adj_4947, n4_adj_4948, n5_adj_4949, 
        n6_adj_4950, n7_adj_4951, n8_adj_4952, n9_adj_4953, n10_adj_4954, 
        n11_adj_4955, n12_adj_4956, n13_adj_4957, n14_adj_4958, n15_adj_4959, 
        n16_adj_4960, n17_adj_4961, n18_adj_4962, n19_adj_4963, n20_adj_4964, 
        n21_adj_4965, n22_adj_4966, n23_adj_4967, n24_adj_4968, n25_adj_4969, 
        n26_adj_4970, n27_adj_4971, n28_adj_4972, n29_adj_4973, n30_adj_4974, 
        n31_adj_4975, n32_adj_4976, n33_adj_4977, n34_adj_4978, n35_adj_4979, 
        n36_adj_4980, n37_adj_4981, n15333, n55, n15332, n15331, 
        n52, n15330, n15329, n49, n15328, n15327, n15326, n46, 
        n15448, n15447, n15446, n15445, n15444, n15443, n15442, 
        n15325, n4_adj_4982, n43, n15324, n15441, n40, n15440, 
        n15439, n15438, n15437, n15323, n15436, n15435, n15434, 
        n15433, n15432, n15431, n15430, n15429, n15428, n15427, 
        n15322, n15426, n15424, n15423, n15422, n34_adj_4983, n78_adj_4984, 
        n81, n84, n87, n90, n93, n96, n99, n102, n105, n108, 
        n111, n114, n117, n120, n123, n126, n129, n132, n135, 
        n138, n141, n144, n147, n150, n153, n156, n159, n162, 
        n165, n168, n171, n174, n177, n180, n183, cout, cout_adj_4985, 
        cout_adj_4986, n78_adj_4987, n81_adj_4988, n84_adj_4989, n87_adj_4990, 
        n90_adj_4991, n93_adj_4992, n96_adj_4993, n99_adj_4994, n102_adj_4995, 
        n105_adj_4996, n108_adj_4997, n111_adj_4998, n114_adj_4999, 
        n117_adj_5000, n120_adj_5001, n123_adj_5002, n126_adj_5003, 
        n129_adj_5004, n132_adj_5005, n135_adj_5006, n138_adj_5007, 
        n141_adj_5008, n144_adj_5009, n147_adj_5010, n150_adj_5011, 
        n153_adj_5012, n156_adj_5013, n159_adj_5014, n162_adj_5015, 
        n165_adj_5016, n168_adj_5017, n171_adj_5018, n174_adj_5019, 
        n177_adj_5020, n180_adj_5021, n183_adj_5022, n78_adj_5023, n81_adj_5024, 
        n84_adj_5025, n87_adj_5026, n90_adj_5027, n93_adj_5028, n96_adj_5029, 
        n99_adj_5030, n102_adj_5031, n105_adj_5032, n108_adj_5033, n111_adj_5034, 
        n114_adj_5035, n117_adj_5036, n120_adj_5037, n123_adj_5038, 
        n126_adj_5039, n129_adj_5040, n132_adj_5041, n135_adj_5042, 
        n138_adj_5043, n141_adj_5044, n144_adj_5045, n147_adj_5046, 
        n150_adj_5047, n153_adj_5048, n156_adj_5049, n159_adj_5050, 
        n162_adj_5051, n165_adj_5052, n168_adj_5053, n171_adj_5054, 
        n174_adj_5055, n177_adj_5056, n180_adj_5057, n183_adj_5058, 
        n32_adj_5059, n38_adj_5060, n41_adj_5061, n44_adj_5062, n47_adj_5063, 
        n50_adj_5064, n53_adj_5065, n56_adj_5066, n59_adj_5067, n62_adj_5068, 
        n65_adj_5069, n68_adj_5070, n71_adj_5071, cout_adj_5072, cout_adj_5073, 
        cout_adj_5074, cout_adj_5075, cout_adj_5076, n28_adj_5077, n31_adj_5078, 
        n34_adj_5079, n37_adj_5080, n40_adj_5081, n43_adj_5082, n46_adj_5083, 
        n49_adj_5084, n52_adj_5085, n55_adj_5086, n58_adj_5087, n61_adj_5088, 
        n78_adj_5089, n81_adj_5090, n84_adj_5091, n87_adj_5092, n90_adj_5093, 
        n93_adj_5094, n96_adj_5095, n99_adj_5096, n102_adj_5097, n105_adj_5098, 
        n108_adj_5099, n111_adj_5100, n114_adj_5101, n117_adj_5102, 
        n120_adj_5103, n123_adj_5104, n126_adj_5105, n129_adj_5106, 
        n132_adj_5107, n135_adj_5108, n138_adj_5109, n141_adj_5110, 
        n144_adj_5111, n147_adj_5112, n150_adj_5113, n153_adj_5114, 
        n156_adj_5115, n159_adj_5116, n162_adj_5117, n165_adj_5118, 
        n168_adj_5119, n171_adj_5120, n174_adj_5121, n177_adj_5122, 
        n180_adj_5123, n183_adj_5124, n15321, n15320, n15318, n15317, 
        n15316, n15315, n15314, n15313, n15311, n15310, n15309, 
        n15308, n15307, n15306, n15305, n15304, n15303, n15302, 
        n15301, n15300, n15299, n15298, n15297, n15296, n15295, 
        n15294, n15290, n15289, n15288, n15287, n15286, n15285, 
        n15284, cout_adj_5125, cout_adj_5126, n78_adj_5127, n81_adj_5128, 
        n84_adj_5129, n87_adj_5130, n90_adj_5131, n93_adj_5132, n96_adj_5133, 
        n99_adj_5134, n102_adj_5135, n105_adj_5136, n108_adj_5137, n111_adj_5138, 
        n114_adj_5139, n117_adj_5140, n120_adj_5141, n123_adj_5142, 
        n126_adj_5143, n129_adj_5144, n132_adj_5145, n135_adj_5146, 
        n138_adj_5147, n141_adj_5148, n144_adj_5149, n147_adj_5150, 
        n150_adj_5151, n153_adj_5152, n156_adj_5153, n159_adj_5154, 
        n162_adj_5155, n165_adj_5156, n168_adj_5157, n171_adj_5158, 
        n174_adj_5159, n177_adj_5160, n180_adj_5161, n183_adj_5162, 
        cout_adj_5163, cout_adj_5164, cout_adj_5165, cout_adj_5166, 
        n28_adj_5167, n31_adj_5168, n34_adj_5169, n37_adj_5170, n40_adj_5171, 
        n43_adj_5172, n46_adj_5173, n49_adj_5174, n52_adj_5175, n55_adj_5176, 
        n58_adj_5177, n61_adj_5178, n22_adj_5179, n25_adj_5180, n28_adj_5181, 
        n31_adj_5182, n34_adj_5183, n37_adj_5184, n40_adj_5185, n43_adj_5186, 
        n46_adj_5187, n78_adj_5188, n81_adj_5189, n84_adj_5190, n87_adj_5191, 
        n90_adj_5192, n93_adj_5193, n96_adj_5194, n99_adj_5195, n102_adj_5196, 
        n105_adj_5197, n108_adj_5198, n111_adj_5199, n114_adj_5200, 
        n117_adj_5201, n120_adj_5202, n123_adj_5203, n126_adj_5204, 
        n129_adj_5205, n132_adj_5206, n135_adj_5207, n138_adj_5208, 
        n141_adj_5209, n144_adj_5210, n147_adj_5211, n150_adj_5212, 
        n153_adj_5213, n156_adj_5214, n159_adj_5215, n162_adj_5216, 
        n165_adj_5217, n168_adj_5218, n171_adj_5219, n174_adj_5220, 
        n177_adj_5221, n180_adj_5222, n183_adj_5223, n22_adj_5224, n25_adj_5225, 
        n28_adj_5226, n31_adj_5227, n34_adj_5228, n37_adj_5229, n40_adj_5230, 
        n43_adj_5231, n46_adj_5232, n78_adj_5233, n81_adj_5234, n84_adj_5235, 
        n87_adj_5236, n90_adj_5237, n93_adj_5238, n96_adj_5239, n99_adj_5240, 
        n102_adj_5241, n105_adj_5242, n108_adj_5243, n111_adj_5244, 
        n114_adj_5245, n117_adj_5246, n120_adj_5247, n123_adj_5248, 
        n126_adj_5249, n129_adj_5250, n132_adj_5251, n135_adj_5252, 
        n138_adj_5253, n141_adj_5254, n144_adj_5255, n147_adj_5256, 
        n150_adj_5257, n153_adj_5258, n156_adj_5259, n159_adj_5260, 
        n162_adj_5261, n165_adj_5262, n168_adj_5263, n171_adj_5264, 
        n174_adj_5265, n177_adj_5266, n180_adj_5267, n183_adj_5268, 
        n78_adj_5269, n81_adj_5270, n84_adj_5271, n87_adj_5272, n90_adj_5273, 
        n93_adj_5274, n96_adj_5275, n99_adj_5276, n102_adj_5277, n105_adj_5278, 
        n108_adj_5279, n111_adj_5280, n114_adj_5281, n117_adj_5282, 
        n120_adj_5283, n123_adj_5284, n126_adj_5285, n129_adj_5286, 
        n132_adj_5287, n135_adj_5288, n138_adj_5289, n141_adj_5290, 
        n144_adj_5291, n147_adj_5292, n150_adj_5293, n153_adj_5294, 
        n156_adj_5295, n159_adj_5296, n162_adj_5297, n165_adj_5298, 
        n168_adj_5299, n171_adj_5300, n174_adj_5301, n177_adj_5302, 
        n180_adj_5303, n183_adj_5304, cout_adj_5305, n15283, n15282, 
        n15281, n15280, n15279, n15278, n15277, n15276, n15275, 
        n15274, n15273, n15272, n15271, n15270, n15269, n15268, 
        n15267, n15266, n15265, n15264, n15263, n15262, n15261, 
        n15260, n15259, n15258, n15257, n15256, n15255, n15254, 
        n15253, n15252, n15251, n15250, n15249, n15248, cout_adj_5306, 
        cout_adj_5307, cout_adj_5308, cout_adj_5309, cout_adj_5310, 
        n78_adj_5311, n81_adj_5312, n84_adj_5313, n87_adj_5314, n90_adj_5315, 
        n93_adj_5316, n96_adj_5317, n99_adj_5318, n102_adj_5319, n105_adj_5320, 
        n108_adj_5321, n111_adj_5322, n114_adj_5323, n117_adj_5324, 
        n120_adj_5325, n123_adj_5326, n126_adj_5327, n129_adj_5328, 
        n132_adj_5329, n135_adj_5330, n138_adj_5331, n141_adj_5332, 
        n144_adj_5333, n147_adj_5334, n150_adj_5335, n153_adj_5336, 
        n156_adj_5337, n159_adj_5338, n162_adj_5339, n165_adj_5340, 
        n168_adj_5341, n171_adj_5342, n174_adj_5343, n177_adj_5344, 
        n180_adj_5345, n183_adj_5346, n134, n137, n140, n143, n146, 
        n149, n152, n155, n158, n161, n164, n167, n170, n173, 
        n176, n179, n182, n185, n188, n191, n194, n197, n200, 
        n203, n206, n209, n212, n215, n218, n221, n224, n227, 
        n230, n233, n236, n239, n242, n245, n248, n251, n254, 
        n257, n260, n263, n266, n269, n272, n275, n278, n281, 
        n284, n287, n290, n293, n296, n299, n302, n305, n308, 
        n311, n314, n317, n320, n323, n15247, n15246, n15245, 
        n15244, n15243, n15242, n15241, n15240, n15239, n15238, 
        cout_adj_5347, n24_adj_5348, n27_adj_5349, n30_adj_5350, n33_adj_5351, 
        n36_adj_5352, n39, n42, n45, n48, n78_adj_5353, n81_adj_5354, 
        n84_adj_5355, n87_adj_5356, n90_adj_5357, n93_adj_5358, n96_adj_5359, 
        n99_adj_5360, n102_adj_5361, n105_adj_5362, n108_adj_5363, n111_adj_5364, 
        n114_adj_5365, n117_adj_5366, n120_adj_5367, n123_adj_5368, 
        n126_adj_5369, n129_adj_5370, n132_adj_5371, n135_adj_5372, 
        n138_adj_5373, n141_adj_5374, n144_adj_5375, n147_adj_5376, 
        n150_adj_5377, n153_adj_5378, n156_adj_5379, n159_adj_5380, 
        n162_adj_5381, n165_adj_5382, n168_adj_5383, n171_adj_5384, 
        n174_adj_5385, n177_adj_5386, n180_adj_5387, n183_adj_5388, 
        n78_adj_5389, n81_adj_5390, n84_adj_5391, n87_adj_5392, n90_adj_5393, 
        n93_adj_5394, n96_adj_5395, n99_adj_5396, n102_adj_5397, n105_adj_5398, 
        n108_adj_5399, n111_adj_5400, n114_adj_5401, n117_adj_5402, 
        n120_adj_5403, n123_adj_5404, n126_adj_5405, n129_adj_5406, 
        n132_adj_5407, n135_adj_5408, n138_adj_5409, n141_adj_5410, 
        n144_adj_5411, n147_adj_5412, n150_adj_5413, n153_adj_5414, 
        n156_adj_5415, n159_adj_5416, n162_adj_5417, n165_adj_5418, 
        n168_adj_5419, n171_adj_5420, n174_adj_5421, n177_adj_5422, 
        n180_adj_5423, n183_adj_5424, n78_adj_5425, n81_adj_5426, n84_adj_5427, 
        n87_adj_5428, n90_adj_5429, n93_adj_5430, n96_adj_5431, n99_adj_5432, 
        n102_adj_5433, n105_adj_5434, n108_adj_5435, n111_adj_5436, 
        n114_adj_5437, n117_adj_5438, n120_adj_5439, n123_adj_5440, 
        n126_adj_5441, n129_adj_5442, n132_adj_5443, n135_adj_5444, 
        n138_adj_5445, n141_adj_5446, n144_adj_5447, n147_adj_5448, 
        n150_adj_5449, n153_adj_5450, n156_adj_5451, n159_adj_5452, 
        n162_adj_5453, n165_adj_5454, n168_adj_5455, n171_adj_5456, 
        n174_adj_5457, n177_adj_5458, n180_adj_5459, n183_adj_5460, 
        n24_adj_5461, n27_adj_5462, n30_adj_5463, n33_adj_5464, n36_adj_5465, 
        n39_adj_5466, n42_adj_5467, n45_adj_5468, n48_adj_5469, n34_adj_5470, 
        n40_adj_5471, n43_adj_5472, n46_adj_5473, n49_adj_5474, n52_adj_5475, 
        n55_adj_5476, n58_adj_5477, n61_adj_5478, n64_adj_5479, n67_adj_5480, 
        n70_adj_5481, n73_adj_5482, n34_adj_5483, n40_adj_5484, n43_adj_5485, 
        n46_adj_5486, n49_adj_5487, n52_adj_5488, n55_adj_5489, n58_adj_5490, 
        n61_adj_5491, n64_adj_5492, n67_adj_5493, n70_adj_5494, n73_adj_5495, 
        n76_adj_5496, n79_adj_5497, n82, n85, n88, n91, n94, n97, 
        n100, n103, n106, n109, n112, n115, n118, n78_adj_5498, 
        n81_adj_5499, n84_adj_5500, n87_adj_5501, n90_adj_5502, n93_adj_5503, 
        n96_adj_5504, n99_adj_5505, n102_adj_5506, n105_adj_5507, n108_adj_5508, 
        n111_adj_5509, n114_adj_5510, n117_adj_5511, n120_adj_5512, 
        n123_adj_5513, n126_adj_5514, n129_adj_5515, n132_adj_5516, 
        n135_adj_5517, n138_adj_5518, n141_adj_5519, n144_adj_5520, 
        n147_adj_5521, n150_adj_5522, n153_adj_5523, n156_adj_5524, 
        n159_adj_5525, n162_adj_5526, n165_adj_5527, n168_adj_5528, 
        n171_adj_5529, n174_adj_5530, n177_adj_5531, n180_adj_5532, 
        n183_adj_5533, n32_adj_5534, n38_adj_5535, n41_adj_5536, n44_adj_5537, 
        n47_adj_5538, n50_adj_5539, n53_adj_5540, n56_adj_5541, n59_adj_5542, 
        n62_adj_5543, n65_adj_5544, n68_adj_5545, n71_adj_5546, n78_adj_5547, 
        n81_adj_5548, n84_adj_5549, n87_adj_5550, n90_adj_5551, n93_adj_5552, 
        n96_adj_5553, n99_adj_5554, n102_adj_5555, n105_adj_5556, n108_adj_5557, 
        n111_adj_5558, n114_adj_5559, n117_adj_5560, n120_adj_5561, 
        n123_adj_5562, n126_adj_5563, n129_adj_5564, n132_adj_5565, 
        n135_adj_5566, n138_adj_5567, n141_adj_5568, n144_adj_5569, 
        n147_adj_5570, n150_adj_5571, n153_adj_5572, n156_adj_5573, 
        n159_adj_5574, n162_adj_5575, n165_adj_5576, n168_adj_5577, 
        n171_adj_5578, n174_adj_5579, n177_adj_5580, n180_adj_5581, 
        n183_adj_5582, n78_adj_5583, n81_adj_5584, n84_adj_5585, n87_adj_5586, 
        n90_adj_5587, n93_adj_5588, n96_adj_5589, n99_adj_5590, n102_adj_5591, 
        n105_adj_5592, n108_adj_5593, n111_adj_5594, n114_adj_5595, 
        n117_adj_5596, n120_adj_5597, n32_adj_5598, n38_adj_5599, n41_adj_5600, 
        n44_adj_5601, n47_adj_5602, n50_adj_5603, n53_adj_5604, n56_adj_5605, 
        n59_adj_5606, n62_adj_5607, n65_adj_5608, n68_adj_5609, n71_adj_5610, 
        n32_adj_5611, n38_adj_5612, n41_adj_5613, n44_adj_5614, n47_adj_5615, 
        n50_adj_5616, n53_adj_5617, n56_adj_5618, n59_adj_5619, n62_adj_5620, 
        n65_adj_5621, n68_adj_5622, n71_adj_5623, n78_adj_5624, n81_adj_5625, 
        n84_adj_5626, n87_adj_5627, n90_adj_5628, n93_adj_5629, n96_adj_5630, 
        n99_adj_5631, n102_adj_5632, n105_adj_5633, n108_adj_5634, n111_adj_5635, 
        n114_adj_5636, n117_adj_5637, n120_adj_5638, n123_adj_5639, 
        n126_adj_5640, n129_adj_5641, n132_adj_5642, n135_adj_5643, 
        n138_adj_5644, n141_adj_5645, n144_adj_5646, n147_adj_5647, 
        n150_adj_5648, n153_adj_5649, n156_adj_5650, n159_adj_5651, 
        n162_adj_5652, n165_adj_5653, n168_adj_5654, n171_adj_5655, 
        n174_adj_5656, n177_adj_5657, n180_adj_5658, n183_adj_5659, 
        n15537, n15421, n15420, n16245, clk_80mhz_enable_1445, n15419, 
        n15418, n15558, n15557, n15417, n15416, n15415, n15556, 
        n15414, n15413, n15555, n15554, n15412, n15411, n15553, 
        n15552, n15410, n15409, n15408, n15407, n15405, n15404, 
        n15403, n15402, n15541, n15401, n15400, n15399, n15849, 
        n15398, n15848, n15397, n15847, n15846, n15540, n15551, 
        n15845, n15550, n15844, n15396, n15842, n15395, n15841, 
        n15549, n15840, n15394, n15839, n15393, n15838, n15837, 
        n15836, n15548, n15835, n15834, n15833, n15832, n15547, 
        n15831, n15830, n15829, n15828, n15392, n15827, n15391, 
        n15826, n15546, n15825, n15824, n15823, n11345, n11351, 
        n11353, n11355, n11357, n11359, n15822, n15821, n15820, 
        n11323, n15819, n132_adj_5660, n11335, n135_adj_5661, n11333, 
        n138_adj_5662, n11331, n141_adj_5663, n144_adj_5664, n147_adj_5665, 
        n150_adj_5666, n153_adj_5667, n156_adj_5668, n159_adj_5669, 
        n162_adj_5670, n165_adj_5671, n168_adj_5672, n171_adj_5673, 
        n174_adj_5674, n177_adj_5675, n15818, n180_adj_5676, n11301, 
        n183_adj_5677, n15598, n186, n11349, n189, n192, n15597, 
        n195, n198, n11395, n201, n204, n11393, n207, n15817, 
        n210, n15816, n213, n11610, n216, n11387, n219, n222, 
        n11385, n225, n15545, n228, n11381, n231, n15815, n234, 
        n15814, n237, n11303, n240, n243, n246, n249, n15813, 
        n252, n255, n15596, n258, n15812, n261, n15595, n264, 
        n11347, n267, n15811, n270, n273, n276, n15594, n279, 
        n282, n285, n288, n291, n294, n15538, n297, n300, n303, 
        n306, n11375, n309, n15807, n312, n15806, n315, n11377, 
        n318, n321, n15237, n15236, n15235, n15234, n15233, n15232, 
        n15231, n15230, n15229, n15228, n15227, n15226, n15225, 
        n15224, n15222, n15221, n14314, n14313, n14312, n2_adj_5678, 
        n4_adj_5679, n6_adj_5680, n8_adj_5681, n10_adj_5682, n12_adj_5683, 
        n14_adj_5684, n16_adj_5685, n18_adj_5686, n20_adj_5687, n22_adj_5688, 
        n24_adj_5689, n26_adj_5690, n28_adj_5691, n30_adj_5692, n32_adj_5693, 
        n34_adj_5694, n36_adj_5695, n38_adj_5696, n40_adj_5697, n42_adj_5698, 
        n44_adj_5699, n46_adj_5700, n48_adj_5701, n52_adj_5702, n55_adj_5703, 
        n58_adj_5704, n61_adj_5705, n64_adj_5706, n67_adj_5707, n70_adj_5708, 
        n73_adj_5709, n76_adj_5710, n79_adj_5711, n15593, n82_adj_5712, 
        n85_adj_5713, n15592, n88_adj_5714, n91_adj_5715, n15805, 
        n94_adj_5716, n15591, n97_adj_5717, n100_adj_5718, n103_adj_5719, 
        n106_adj_5720, n15804, n109_adj_5721, n15803, n112_adj_5722, 
        n14311, n115_adj_5723, n15590, n118_adj_5724, n15802, n121, 
        n15801, n15800, n15589, n15588, n15587, n15586, n15799, 
        n15798, n15797, n15796, n15795, n11_adj_5725, n15585, n15793, 
        n15544, n15792, n15791, n15584, n15790, n15789, n13_adj_5726, 
        n15788, n15787, n15786, n15785, n11259, n15583, n15582, 
        clk_80mhz_enable_1447, n15220, n78_adj_5727, n15219, n81_adj_5728, 
        n15784, n84_adj_5729, n87_adj_5730, n15783, n90_adj_5731, 
        n15782, n93_adj_5732, n96_adj_5733, n99_adj_5734, n15781, 
        n102_adj_5735, n16238, n105_adj_5736, n15780, n108_adj_5737, 
        n15779, n111_adj_5738, n114_adj_5739, n11309, n117_adj_5740, 
        n11311, n120_adj_5741, n15581, n123_adj_5742, n15580, n126_adj_5743, 
        n15778, n129_adj_5744, n132_adj_5745, n15579, n135_adj_5746, 
        n15777, n138_adj_5747, n15578, n141_adj_5748, n15577, n144_adj_5749, 
        n147_adj_5750, n15576, n150_adj_5751, n15575, n153_adj_5752, 
        n156_adj_5753, n15776, n159_adj_5754, n15574, n162_adj_5755, 
        n15573, n165_adj_5756, n15572, n168_adj_5757, n15571, n171_adj_5758, 
        n174_adj_5759, n15570, n177_adj_5760, n15569, n180_adj_5761, 
        n183_adj_5762, n15568, n15772, n15771, n15770, n15769, n15567, 
        n15768, n15767, n15566, n15766, n17127, n15565, n15564, 
        n15563, n15764, n15539, n15543, n15763, n15762, n15562, 
        n15761, n15760, n15759, n15758, n15757, n15561, n15560, 
        n15756, n15755, n11169, n15754, n15753, n11397, n15559, 
        n15752, n15751, n15750, n15749, n15748, n11373, n11339, 
        n11337, n11371, n11369, n11367, n11363, n15542, n17178, 
        n11361, n15747, n11317, n11319, n11327, n11341, n15743, 
        n11307, n15218, n15217, n15216, n15215, n15214, n15213, 
        n15212, n15211, n15210, n15209, n15208, n78_adj_5763, n15207, 
        n81_adj_5764, n15206, n84_adj_5765, n15205, n87_adj_5766, 
        n15204, n90_adj_5767, n15203, n93_adj_5768, n15202, n96_adj_5769, 
        n15201, n99_adj_5770, n15200, n102_adj_5771, n15199, n105_adj_5772, 
        n15198, n108_adj_5773, n15197, n111_adj_5774, n15196, n114_adj_5775, 
        n15195, n117_adj_5776, n15194, n120_adj_5777, n15193, n123_adj_5778, 
        n15192, n126_adj_5779, n15191, n129_adj_5780, n15190, n132_adj_5781, 
        n15189, n135_adj_5782, n15188, n138_adj_5783, n15187, n141_adj_5784, 
        n15185, n144_adj_5785, n15184, n147_adj_5786, n15183, n150_adj_5787, 
        n15182, n153_adj_5788, n15181, n156_adj_5789, n15180, n159_adj_5790, 
        n15179, n162_adj_5791, n15178, n165_adj_5792, n15177, n168_adj_5793, 
        n15176, n171_adj_5794, n15175, n174_adj_5795, n15174, n177_adj_5796, 
        n15173, n180_adj_5797, n15172, n183_adj_5798, n15171, n15170, 
        n15169, n15168, n15167, n15166, n15165, n15164, n15163, 
        n15162, n15161, n15160, n15159, n15158, n15157, n15156, 
        n15155, n15154, n15153, n15152, n15151, n15150, n15149, 
        n15148, n15147, n15146, n15145, n15144, n15143, n15142, 
        n15141, n15140, n15139, n15138, n15137, n15136, n15135, 
        n15134, n15133, n15132, n15131, n15130, n15129, n15128, 
        n15127, n15126, n15125, n15124, n15123, n15122, n15121, 
        n15120, n15119, n15118, n15117, n15116, n15115, n15114, 
        n15113, n15112, n15111, n15110, n15109, n15108, n15107, 
        n15106, n15105, n15104, n15103, n15102, n15101, n15100, 
        n15098, n15097, n15096, n15095, n78_adj_5799, n15094, n81_adj_5800, 
        n15093, n84_adj_5801, n15092, n87_adj_5802, n15091, n90_adj_5803, 
        n15090, n93_adj_5804, n15089, n96_adj_5805, n15088, n99_adj_5806, 
        n15087, n102_adj_5807, n15086, n105_adj_5808, n15085, n108_adj_5809, 
        n15084, n111_adj_5810, n15083, n114_adj_5811, n15082, n117_adj_5812, 
        n15081, n120_adj_5813, n123_adj_5814, n126_adj_5815, n15077, 
        n129_adj_5816, n15076, n132_adj_5817, n15075, n135_adj_5818, 
        n15074, n138_adj_5819, n15073, n141_adj_5820, n15072, n144_adj_5821, 
        n15071, n147_adj_5822, n150_adj_5823, n15069, n153_adj_5824, 
        n15068, n156_adj_5825, n15067, n159_adj_5826, n15066, n162_adj_5827, 
        n15065, n165_adj_5828, n15064, n168_adj_5829, n15063, n171_adj_5830, 
        n15062, n174_adj_5831, n15061, n177_adj_5832, n15060, n180_adj_5833, 
        n15059, n183_adj_5834, n15057, n15056, n15055, n15054, n15053, 
        n15052, n15051, n15050, n15049, n15048, n15047, n15046, 
        n15045, n15044, n15043, n15042, n15041, n15040, n15039, 
        n15038, n15037, n15036, n15035, n15034, n15033, n15032, 
        n15031, n15030, n15029, n15028, n15027, n15026, n15025, 
        n15024, n15023, n15022, n15021, n15020, n15019, n15018, 
        n15017, n15016, n15015, n15014, n15013, n15012, n34_adj_5835, 
        n15011, n15010, n40_adj_5836, n15008, n43_adj_5837, n15007, 
        n46_adj_5838, n15006, n49_adj_5839, n15005, n52_adj_5840, 
        n15004, n55_adj_5841, n15003, n58_adj_5842, n15002, n61_adj_5843, 
        n15001, n64_adj_5844, n15000, n67_adj_5845, n14999, n70_adj_5846, 
        n14998, n73_adj_5847, n14997, n14996, n14995, n14994, n14993, 
        n14992, n14991, n14987, n14986, n14985, n14984, n14983, 
        n14982, n14981, n14979, n14978, n14977, n14976, n14975, 
        n14974, n14973, n14972, n14971, n14970, n14969, n14968, 
        n14967, n14966, n14965, n14964, n14963, n14962, n14958, 
        n14957, n14956, n14955, n14954, n14953, n14952, n14951, 
        n14950, n14949, n14948, n14947, n14946, n14945, n14944, 
        n14943, n14942, n76_adj_5848, n14941, n79_adj_5849, n14940, 
        n82_adj_5850, n14939, n85_adj_5851, n14938, n88_adj_5852, 
        n14937, n91_adj_5853, n14936, n94_adj_5854, n14935, n97_adj_5855, 
        n14934, n100_adj_5856, n14932, n103_adj_5857, n14931, n106_adj_5858, 
        n14930, n109_adj_5859, n14929, n112_adj_5860, n14928, n115_adj_5861, 
        n14927, n118_adj_5862, n14926, n14925, n14924, n14923, n14922, 
        n14921, n14920, n14919, n14918, n14917, n14916, n14915, 
        n14913, n14912, n14911, n14910, n14909, n14908, n14907, 
        n14906, n14905, n14904, n14903, n14902, n14901, n14900, 
        n14899, n14898, n14897, n14896, n14893, n14892, n14891, 
        n14890, n14889, n14888, n14887, n14886, n14885, n14884, 
        n14883, n14882, n14881, n14880, n14879, n14878, n14877, 
        n14876, n14872, n14871, n14870, n14869, n14868, n14867, 
        n14865, n14864, n14863, n14862, n14861, n14860, n14859, 
        n14858, n14857, n14856, n14855, n14854, n14853, n14852, 
        n14851, n14850, n14849, n14848, n14835, n14834, n14833, 
        n14832, n14831, n14830, n14829, n14828, n14827, n14826, 
        n14825, n14819, n14818, n14817, n14816, n14815, n32_adj_5863, 
        n14814, n14813, n14812, n38_adj_5864, n14811, n41_adj_5865, 
        n14810, n44_adj_5866, n14809, n47_adj_5867, n14808, n50_adj_5868, 
        n14807, n53_adj_5869, n14806, n56_adj_5870, n14805, n59_adj_5871, 
        n14804, n62_adj_5872, n14803, n65_adj_5873, n14802, n68_adj_5874, 
        n71_adj_5875, n14800, n14799, n14798, n14797, n14796, n14795, 
        n14794, n14793, n14792, n14791, n14790, n14789, n14788, 
        n14787, n14786, n14785, n14784, n14783, n14782, n14781, 
        n14780, n14779, n14778, n14777, n14776, n14775, n14774, 
        n14773, n14772, n14771, n14770, n14769, n14768, n14767, 
        n14766, n14765, n14764, n14763, n14762, n14761, n14760, 
        n14759, n14758, n14757, n14756, n14755, n14754, n14753, 
        n14752, n14751, n14750, n14749, n14748, n14747, n14746, 
        n14745, n14744, n14743, n14742, n14741, n14740, n14739, 
        n14738, n14737, n14736, n14735, n14734, n14733, n14732, 
        n14731, n14730, n14729, n14728, n14727, n14726, n14725, 
        n14723, n14722, n14721, n14720, n14719, n14718, n14717, 
        n14716, n14715, n14714, n14713, n14712, n14711, n14710, 
        n14709, n14708, n14707, n14706, n14705, n14704, n14703, 
        n14702, n14701, n14700, n14699, n14698, n14697, n14696, 
        n14695, n14694, n14693, n14692, n14691, n14690, n14689, 
        n14688, n14687, n14686, n14685, n14684, n14682, n14681, 
        n14680, n14679, n14678, n14677, n14676, n14675, n14674, 
        n14673, n14672, n14671, n14670, n14669, n14668, n14667, 
        n14666, n34_adj_5876, n14665, n40_adj_5877, n43_adj_5878, 
        n14660, n46_adj_5879, n14659, n49_adj_5880, n14658, n52_adj_5881, 
        n14657, n55_adj_5882, n14656, n58_adj_5883, n14655, n61_adj_5884, 
        n14654, n64_adj_5885, n14653, n67_adj_5886, n14652, n70_adj_5887, 
        n14651, n73_adj_5888, n14650, n14649, n14648, n14647, n14646, 
        n14645, n14644, n14643, n14638, n14637, n14636, n14635, 
        n14634, n14633, n14632, n14631, n14630, n14629, n14628, 
        n14627, n14626, n14625, n14624, n14623, n14622, n14621, 
        n14616, n14615, n14614, n14613, n14612, n14611, n14610, 
        n14609, n14608, n14607, n14606, n14605, n14604, n14603, 
        n14602, n14601, n14600, n14599, n14594, n78_adj_5889, n14593, 
        n81_adj_5890, n14592, n84_adj_5891, n14591, n87_adj_5892, 
        n14590, n90_adj_5893, n14589, n93_adj_5894, n14588, n96_adj_5895, 
        n14587, n99_adj_5896, n14586, n102_adj_5897, n14585, n105_adj_5898, 
        n14584, n108_adj_5899, n14583, n111_adj_5900, n14582, n114_adj_5901, 
        n14581, n117_adj_5902, n14580, n120_adj_5903, n14579, n14578, 
        n14577, n14573, n14572, n14571, n14570, n14569, n14568, 
        n14567, n14566, n14565, n14564, n14563, n14562, n14561, 
        n14560, n14559, n14558, n14557, n14556, n14555, n14554, 
        n14553, n14552, n14551, n14550, n14549, n14548, n14547, 
        n14546, n14545, n14544, n14543, n14542, n14541, n14540, 
        n14539, n14538, n14536, n14535, n14534, n14533, n14532, 
        n14531, n14530, n14529, n14528, n14527, n14526, n14525, 
        n14524, n14523, n14522, n14521, n14520, n14519, n14513, 
        n14512, n14511, n14510, n14509, n14508, n14507, n14506, 
        n14505, n14504, n14503, n14502, n14501, n14500, n14499, 
        n14498, n14497, n14496, n14495, n14494, n14493, n14492, 
        n14491, n14490, n14489, n14488, n14487, n14486, n14485, 
        n14484, n14483, n14482, n14481, n14480, n14479, n14478, 
        n124, n14477, n127, n14476, n130, n14475, n133, n14474, 
        n136, n14473, n139, n14472, n142, n14471, n145, n14470, 
        n148, n14469, n151, n14468, n154, n14467, n157, n14466, 
        n160, n14465, n163, n14464, n166, n14463, n169, n14462, 
        n172, n14461, n175, n14460, n178, n14459, n181, n14458, 
        n184, n14457, n187, n14456, n190, n14455, n193, n14454, 
        n196, n14453, n199, n14452, n202, n14451, n205, n14450, 
        n208, n14449, n211, n14448, n214, n14447, n217, n14446, 
        n220, n14445, n223, n14444, n226, n14443, n229, n14442, 
        n232, n14441, n235, n14440, n238, n14439, n241, n14438, 
        n244, n14437, n247, n14436, n250, n14435, n253, n14434, 
        n256, n14433, n259, n14432, n262, n14431, n265, n14430, 
        n268, n14429, n271, n14428, n274, n14427, n277, n14426, 
        n280, n14425, n283, n14424, n286, n14423, n289, n14422, 
        n292, n14421, n295, n14420, n298, n14419, n301, n14418, 
        n14417, n14416, n14415, n14414, n14413, n14412, n14411, 
        n14410, n14409, n14408, n14407, n14406, n14405, n14404, 
        n14403, n14402, n14401, n14400, n14399, n14398, n14397, 
        n14396, n14395, n14394, n14393, n14392, n14391, n14390, 
        n14389, n14388, n14387, n14386, n14385, n14384, n14383, 
        n14382, n14381, n14380, n14379, n14378, n14377, n14376, 
        n14375, n14374, n14373, n14372, n14371, n14370, n14369, 
        n14368, n14367, n14365, n14364, n14363, n14362, n14360, 
        n14359, n14358, n14357, n130_adj_5904, n14356, n133_adj_5905, 
        n14355, n136_adj_5906, n14354, n139_adj_5907, n14353, n142_adj_5908, 
        n14352, n145_adj_5909, n14351, n148_adj_5910, n14350, n151_adj_5911, 
        n14349, n154_adj_5912, n14348, n157_adj_5913, n14347, n160_adj_5914, 
        n14346, n163_adj_5915, n14345, n166_adj_5916, n14344, n169_adj_5917, 
        n14343, n172_adj_5918, n175_adj_5919, n178_adj_5920, n14339, 
        n181_adj_5921, n14338, n184_adj_5922, n14337, n187_adj_5923, 
        n14336, n190_adj_5924, n14335, n193_adj_5925, n14334, n196_adj_5926, 
        n14333, n199_adj_5927, n14332, n202_adj_5928, n14331, n205_adj_5929, 
        n14330, n208_adj_5930, n14329, n211_adj_5931, n14328, n214_adj_5932, 
        n14327, n217_adj_5933, n14326, n220_adj_5934, n14325, n223_adj_5935, 
        n14324, n226_adj_5936, n14323, n229_adj_5937, n14322, n232_adj_5938, 
        n14321, n235_adj_5939, n14320, n238_adj_5940, n14319, n241_adj_5941, 
        n14318, n244_adj_5942, n14317, n247_adj_5943, n14316, n250_adj_5944, 
        n14315, n253_adj_5945, n256_adj_5946, n259_adj_5947, n262_adj_5948, 
        n265_adj_5949, n268_adj_5950, n271_adj_5951, n274_adj_5952, 
        n277_adj_5953, n280_adj_5954, n283_adj_5955, n286_adj_5956, 
        n289_adj_5957, n292_adj_5958, n295_adj_5959, n298_adj_5960, 
        n301_adj_5961, n304, n307, n310, n313, n316, n32_adj_5962, 
        n38_adj_5963, n41_adj_5964, n44_adj_5965, n47_adj_5966, n50_adj_5967, 
        n53_adj_5968, n56_adj_5969, n59_adj_5970, n62_adj_5971, n65_adj_5972, 
        n68_adj_5973, n71_adj_5974, n34_adj_5975, n40_adj_5976, n43_adj_5977, 
        n46_adj_5978, n49_adj_5979, n52_adj_5980, n55_adj_5981, n58_adj_5982, 
        n61_adj_5983, n64_adj_5984, n67_adj_5985, n70_adj_5986, n73_adj_5987, 
        n16607, n17177, n14310, n14309, n14308, n16957, n14307, 
        n14306, n34_adj_5988, n40_adj_5989, n43_adj_5990, n46_adj_5991, 
        n49_adj_5992, n52_adj_5993, n16451, n55_adj_5994, n58_adj_5995, 
        n61_adj_5996, n64_adj_5997, n67_adj_5998, n70_adj_5999, n73_adj_6000, 
        n14305, n14304, n29_adj_6001, n16220, n17139, n16203, n17137, 
        n14303, n17136, n17049, n16409, n17048, n17163, n17162, 
        n14302, n17043, n17174, n17279, n17158, n14301, n34_adj_6002, 
        n40_adj_6003, n17157, n43_adj_6004, n46_adj_6005, n49_adj_6006, 
        n17173, n52_adj_6007, n55_adj_6008, n58_adj_6009, n17289, 
        n61_adj_6010, n17155, n64_adj_6011, n67_adj_6012, n70_adj_6013, 
        n73_adj_6014, n17278, n17153, n17172;
    
    VHI i2 (.Z(VCC_net));
    \uart_rx(CLKS_PER_BIT=87)  uart_rx_inst (.clk_80mhz(clk_80mhz), .rx_serial_c(rx_serial_c), 
            .rx_byte1({rx_byte1}), .rx_data_valid1(rx_data_valid1), .GND_net(GND_net), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(209[7] 214[6])
    CCU2C _add_1_1250_add_4_3 (.A0(square_sum[11]), .B0(amdemod_d_11__N_1851[13]), 
          .C0(n17132), .D0(amdemod_d_11__N_1850[13]), .A1(n17131), .B1(amdemod_d_11__N_1850[0]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15462), .COUT(n15463), .S0(n68), 
          .S1(n65));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1250_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_1250_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1250_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1250_add_4_3.INJECT1_1 = "NO";
    FD1S3AX rx_byte_i1 (.D(rx_byte1[0]), .CK(clk_80mhz), .Q(led_c_0));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam rx_byte_i1.GSR = "ENABLED";
    AMDemodulator AMDemodulator_inst (.cic_sine_clk(cic_sine_clk), .cic_cosine_out({cic_cosine_out}), 
            .\data_in_reg_11__N_2339[0] (data_in_reg_11__N_2339[0]), .\square_sum[22] (square_sum[22]), 
            .\square_sum[23] (square_sum[23]), .n11179(n11179), .amdemod_d_11__N_1874(amdemod_d_11__N_1874), 
            .amdemod_d_11__N_2023(amdemod_d_11__N_2023), .amdemod_d_11__N_2146(amdemod_d_11__N_2146), 
            .amdemod_d_11__N_2149(amdemod_d_11__N_2149), .amdemod_d_11__N_2020(amdemod_d_11__N_2020), 
            .amdemod_d_11__N_2281(amdemod_d_11__N_2281), .amdemod_d_11__N_2284(amdemod_d_11__N_2284), 
            .amdemod_d_11__N_2026(amdemod_d_11__N_2026), .amdemod_d_11__N_2152(amdemod_d_11__N_2152), 
            .\square_sum[21] (square_sum[21]), .\square_sum[20] (square_sum[20]), 
            .n4(n4_adj_4982), .\amdemod_d_11__N_1870[13] (amdemod_d_11__N_1870[13]), 
            .\amdemod_d_11__N_1871[13] (amdemod_d_11__N_1871[13]), .n17128(n17128), 
            .n80(n80), .n79(n79), .n78(n78), .n77(n77), .n76(n76), 
            .n75(n75), .n74(n74), .n73(n73), .n72(n72), .n71(n71_adj_4749), 
            .n70(n70), .n69(n69), .n68(n68_adj_4750), .n67(n67), .n66(n66_adj_4752), 
            .n65(n65_adj_4753), .n64(n64_adj_4754), .n63(n63_adj_4755), 
            .n62(n62_adj_4756), .n61(n61), .n60(n60), .n59(n59_adj_4758), 
            .n58(n58), .n57(n57), .VCC_net(VCC_net), .GND_net(GND_net), 
            .n17146(n17146), .n17157(n17157), .n34(n34_adj_5988), .n34_adj_225(n34_adj_5835), 
            .n17134(n17134), .n32(n32_adj_5059), .n32_adj_226(n32_adj_4742), 
            .n71_adj_227(n71_adj_5071), .n71_adj_228(n71_adj_4730), .n73_adj_229(n73_adj_6000), 
            .n73_adj_230(n73_adj_5847), .n68_adj_231(n68_adj_5070), .n68_adj_232(n68_adj_4731), 
            .n70_adj_233(n70_adj_5999), .n70_adj_234(n70_adj_5846), .n65_adj_235(n65_adj_5069), 
            .n65_adj_236(n65_adj_4732), .n67_adj_237(n67_adj_5998), .n67_adj_238(n67_adj_5845), 
            .n62_adj_239(n62_adj_5068), .n62_adj_240(n62_adj_4733), .n64_adj_241(n64_adj_5997), 
            .n64_adj_242(n64_adj_5844), .n59_adj_243(n59_adj_5067), .n59_adj_244(n59_adj_4734), 
            .n61_adj_245(n61_adj_5996), .n61_adj_246(n61_adj_5843), .n53(n53_adj_5065), 
            .n53_adj_247(n53_adj_4736), .n55(n55_adj_5994), .n55_adj_248(n55_adj_5841), 
            .n46(n46_adj_5978), .n46_adj_249(n46_adj_6005), .n17132(n17132), 
            .n56(n56_adj_5066), .n56_adj_250(n56_adj_4735), .n58_adj_251(n58_adj_5995), 
            .n58_adj_252(n58_adj_5842), .n41(n41), .n41_adj_253(n41_adj_5964), 
            .n50(n50_adj_5064), .n50_adj_254(n50_adj_4737), .n52(n52_adj_5993), 
            .n52_adj_255(n52_adj_5840), .mult_i_b({mult_i_b}), .mult_result_i({mult_result_i}), 
            .n43(n43_adj_5977), .n43_adj_256(n43_adj_6004), .n47(n47_adj_5063), 
            .n47_adj_257(n47_adj_4738), .n49(n49_adj_5992), .n49_adj_258(n49_adj_5839), 
            .n38(n38), .n38_adj_259(n38_adj_5963), .n40(n40_adj_5976), 
            .n40_adj_260(n40_adj_6003), .n44(n44_adj_5062), .n44_adj_261(n44_adj_4739), 
            .n46_adj_262(n46_adj_5991), .n46_adj_263(n46_adj_5838), .n71_adj_264(n71_adj_5875), 
            .n71_adj_265(n71_adj_5623), .n17130(n17130), .n41_adj_266(n41_adj_5061), 
            .n41_adj_267(n41_adj_4740), .n43_adj_268(n43_adj_5990), .n43_adj_269(n43_adj_5837), 
            .n73_adj_270(n73_adj_5888), .n73_adj_271(n73_adj_5495), .n68_adj_272(n68_adj_5874), 
            .n68_adj_273(n68_adj_5622), .n70_adj_274(n70_adj_5887), .n70_adj_275(n70_adj_5494), 
            .n65_adj_276(n65_adj_5873), .n65_adj_277(n65_adj_5621), .n67_adj_278(n67_adj_5886), 
            .n67_adj_279(n67_adj_5493), .n62_adj_280(n62_adj_5872), .n62_adj_281(n62_adj_5620), 
            .\amdemod_d_11__N_1850[13] (amdemod_d_11__N_1850[13]), .\amdemod_d_11__N_1851[13] (amdemod_d_11__N_1851[13]), 
            .n17131(n17131), .n17129(n17129), .n64_adj_282(n64_adj_5885), 
            .n64_adj_283(n64_adj_5492), .n59_adj_284(n59_adj_5871), .n59_adj_285(n59_adj_5619), 
            .n38_adj_286(n38_adj_5060), .n38_adj_287(n38_adj_4741), .n61_adj_288(n61_adj_5884), 
            .n61_adj_289(n61_adj_5491), .n40_adj_290(n40_adj_5989), .n40_adj_291(n40_adj_5836), 
            .\amdemod_d_11__N_1880[13] (amdemod_d_11__N_1880[13]), .\amdemod_d_11__N_1881[13] (amdemod_d_11__N_1881[13]), 
            .n56_adj_292(n56_adj_5870), .n56_adj_293(n56_adj_5618), .n71_adj_294(n71), 
            .n71_adj_295(n71_adj_5974), .n73_adj_296(n73_adj_5987), .n73_adj_297(n73_adj_6014), 
            .n58_adj_298(n58_adj_5883), .n58_adj_299(n58_adj_5490), .n53_adj_300(n53_adj_5869), 
            .n53_adj_301(n53_adj_5617), .n55_adj_302(n55_adj_5882), .n55_adj_303(n55_adj_5489), 
            .n50_adj_304(n50_adj_5868), .n50_adj_305(n50_adj_5616), .n34_adj_306(n34_adj_5470), 
            .n34_adj_307(n34_adj_4983), .amdemod_d_11__N_2155(amdemod_d_11__N_2155), 
            .\data_in_reg_11__N_2339[1] (data_in_reg_11__N_2339[1]), .\data_in_reg_11__N_2339[2] (data_in_reg_11__N_2339[2]), 
            .\data_in_reg_11__N_2339[3] (data_in_reg_11__N_2339[3]), .\data_in_reg_11__N_2339[4] (data_in_reg_11__N_2339[4]), 
            .\data_in_reg_11__N_2339[5] (data_in_reg_11__N_2339[5]), .\data_in_reg_11__N_2339[6] (data_in_reg_11__N_2339[6]), 
            .\data_in_reg_11__N_2339[7] (data_in_reg_11__N_2339[7]), .\data_in_reg_11__N_2339[8] (data_in_reg_11__N_2339[8]), 
            .\amdemod_out[9] (amdemod_out[9]), .\amdemod_d_11__N_1860[13] (amdemod_d_11__N_1860[13]), 
            .\amdemod_d_11__N_1861[13] (amdemod_d_11__N_1861[13]), .n17127(n17127), 
            .amdemod_d_11__N_2287(amdemod_d_11__N_2287), .\amdemod_d_11__N_1840[11] (amdemod_d_11__N_1840[11]), 
            .\amdemod_d_11__N_1841[11] (amdemod_d_11__N_1841[11]), .n52_adj_308(n52_adj_5881), 
            .n52_adj_309(n52_adj_5488), .n17163(n17163), .n17137(n17137), 
            .n47_adj_310(n47_adj_5867), .n47_adj_311(n47_adj_5615), .n49_adj_312(n49_adj_5880), 
            .n49_adj_313(n49_adj_5487), .n44_adj_314(n44_adj_5866), .n44_adj_315(n44_adj_5614), 
            .n46_adj_316(n46_adj_5879), .n46_adj_317(n46_adj_5486), .n41_adj_318(n41_adj_5865), 
            .n41_adj_319(n41_adj_5613), .n43_adj_320(n43_adj_5878), .n43_adj_321(n43_adj_5485), 
            .n38_adj_322(n38_adj_5864), .n38_adj_323(n38_adj_5612), .n40_adj_324(n40_adj_5877), 
            .n40_adj_325(n40_adj_5484), .n17133(n17133), .n71_adj_326(n71_adj_5610), 
            .n71_adj_327(n71_adj_5546), .n73_adj_328(n73_adj_5482), .n73_adj_329(n73_adj_4751), 
            .n65_adj_330(n65), .n65_adj_331(n65_adj_5972), .n67_adj_332(n67_adj_5985), 
            .n67_adj_333(n67_adj_6012), .n68_adj_334(n68_adj_5609), .n68_adj_335(n68_adj_5545), 
            .n70_adj_336(n70_adj_5481), .n70_adj_337(n70_adj_4759), .n65_adj_338(n65_adj_5608), 
            .n65_adj_339(n65_adj_5544), .n67_adj_340(n67_adj_5480), .n67_adj_341(n67_adj_4760), 
            .n62_adj_342(n62_adj_5607), .n62_adj_343(n62_adj_5543), .n64_adj_344(n64_adj_5479), 
            .n64_adj_345(n64_adj_4762), .n59_adj_346(n59_adj_5606), .n59_adj_347(n59_adj_5542), 
            .n61_adj_348(n61_adj_5478), .n61_adj_349(n61_adj_4764), .amdemod_d_11__N_2290(amdemod_d_11__N_2290), 
            .amdemod_d_11__N_2293(amdemod_d_11__N_2293), .amdemod_d_11__N_2158(amdemod_d_11__N_2158), 
            .amdemod_d_11__N_2296(amdemod_d_11__N_2296), .amdemod_d_11__N_2161(amdemod_d_11__N_2161), 
            .n56_adj_350(n56), .n56_adj_351(n56_adj_5969), .amdemod_d_11__N_2167(amdemod_d_11__N_2167), 
            .amdemod_d_11__N_2299(amdemod_d_11__N_2299), .n34_adj_352(n34_adj_5876), 
            .n34_adj_353(n34_adj_5483), .n68_adj_354(n68), .n68_adj_355(n68_adj_5973), 
            .n17162(n17162), .amdemod_d_11__N_2302(amdemod_d_11__N_2302), 
            .amdemod_d_11__N_2164(amdemod_d_11__N_2164), .n58_adj_356(n58_adj_5982), 
            .n58_adj_357(n58_adj_6009), .n39(n39_adj_5466), .n39_adj_358(n39), 
            .n52_adj_441({n22_adj_5224, n25_adj_5225, n28_adj_5226, n31_adj_5227, 
            n34_adj_5228, n37_adj_5229, n40_adj_5230, n43_adj_5231, 
            n46_adj_5232}), .n52_adj_442({n22_adj_5179, n25_adj_5180, 
            n28_adj_5181, n31_adj_5182, n34_adj_5183, n37_adj_5184, 
            n40_adj_5185, n43_adj_5186, n46_adj_5187}), .n44_adj_372(n44_adj_5601), 
            .n44_adj_373(n44_adj_5537), .n46_adj_374(n46_adj_5473), .n46_adj_375(n46), 
            .n32_adj_376(n32_adj_5863), .n32_adj_377(n32_adj_5611), .amdemod_d_11__N_2305(amdemod_d_11__N_2305), 
            .n70_adj_378(n70_adj_5986), .n70_adj_379(n70_adj_6013), .\amdemod_d_11__N_1830[1] (amdemod_d_11__N_1830[1]), 
            .n34_adj_380(n34_adj_5975), .n34_adj_381(n34_adj_6002), .n32_adj_382(n32_adj_4715), 
            .n32_adj_383(n32_adj_5962), .n48(n48_adj_5469), .n48_adj_384(n48), 
            .n53_adj_385(n53), .n53_adj_386(n53_adj_5968), .amdemod_d_11__N_2308(amdemod_d_11__N_2308), 
            .amdemod_d_11__N_2311(amdemod_d_11__N_2311), .n41_adj_387(n41_adj_5600), 
            .n41_adj_388(n41_adj_5536), .n36(n36_adj_5465), .n36_adj_389(n36_adj_5352), 
            .n42(n42_adj_5467), .n42_adj_390(n42), .amdemod_d_11__N_2314(amdemod_d_11__N_2314), 
            .amdemod_d_11__N_2209(amdemod_d_11__N_2209), .amdemod_d_11__N_2170(amdemod_d_11__N_2170), 
            .n24(n24_adj_5461), .n24_adj_391(n24_adj_5348), .amdemod_d_11__N_2212(amdemod_d_11__N_2212), 
            .n45(n45_adj_5468), .n45_adj_392(n45), .n30(n30_adj_5463), 
            .n30_adj_393(n30_adj_5350), .n33(n33_adj_5464), .n33_adj_394(n33_adj_5351), 
            .amdemod_d_11__N_2215(amdemod_d_11__N_2215), .n27(n27_adj_5462), 
            .n27_adj_395(n27_adj_5349), .amdemod_d_11__N_2218(amdemod_d_11__N_2218), 
            .amdemod_d_11__N_2221(amdemod_d_11__N_2221), .amdemod_d_11__N_2224(amdemod_d_11__N_2224), 
            .n56_adj_396(n56_adj_5605), .n56_adj_397(n56_adj_5541), .amdemod_d_11__N_2227(amdemod_d_11__N_2227), 
            .amdemod_d_11__N_2230(amdemod_d_11__N_2230), .n6(n6_adj_4757), 
            .amdemod_d_11__N_2065(amdemod_d_11__N_2065), .amdemod_d_11__N_2233(amdemod_d_11__N_2233), 
            .n58_adj_398(n58_adj_5477), .n58_adj_399(n58_adj_4765), .amdemod_d_11__N_2236(amdemod_d_11__N_2236), 
            .amdemod_d_11__N_2068(amdemod_d_11__N_2068), .amdemod_d_11__N_2239(amdemod_d_11__N_2239), 
            .n17279(n17279), .amdemod_d_11__N_2242(amdemod_d_11__N_2242), 
            .n53_adj_400(n53_adj_5604), .n53_adj_401(n53_adj_5540), .n4_adj_402(n4_adj_2948), 
            .amdemod_d_11__N_2071(amdemod_d_11__N_2071), .amdemod_d_11__N_2137(amdemod_d_11__N_2137), 
            .amdemod_d_11__N_2074(amdemod_d_11__N_2074), .n62_adj_403(n62), 
            .n62_adj_404(n62_adj_5971), .n64_adj_405(n64_adj_5984), .n64_adj_406(n64_adj_6011), 
            .amdemod_d_11__N_2140(amdemod_d_11__N_2140), .amdemod_d_11__N_2077(amdemod_d_11__N_2077), 
            .n43_adj_407(n43_adj_5472), .n43_adj_408(n43), .n55_adj_409(n55_adj_5981), 
            .n55_adj_410(n55_adj_6008), .n50_adj_411(n50), .n50_adj_412(n50_adj_5967), 
            .amdemod_d_11__N_2143(amdemod_d_11__N_2143), .amdemod_d_11__N_2083(amdemod_d_11__N_2083), 
            .amdemod_d_11__N_2080(amdemod_d_11__N_2080), .n55_adj_413(n55_adj_5476), 
            .n55_adj_414(n55), .amdemod_d_11__N_2086(amdemod_d_11__N_2086), 
            .n38_adj_415(n38_adj_5599), .n38_adj_416(n38_adj_5535), .n59_adj_417(n59), 
            .n59_adj_418(n59_adj_5970), .amdemod_d_11__N_2089(amdemod_d_11__N_2089), 
            .n40_adj_419(n40_adj_5471), .n40_adj_420(n40), .amdemod_d_11__N_2092(amdemod_d_11__N_2092), 
            .n61_adj_421(n61_adj_5983), .n61_adj_422(n61_adj_6010), .amdemod_d_11__N_2095(amdemod_d_11__N_2095), 
            .amdemod_d_11__N_2098(amdemod_d_11__N_2098), .amdemod_d_11__N_2005(amdemod_d_11__N_2005), 
            .n50_adj_423(n50_adj_5603), .n50_adj_424(n50_adj_5539), .n52_adj_425(n52_adj_5475), 
            .n52_adj_426(n52), .n52_adj_427(n52_adj_5980), .n52_adj_428(n52_adj_6007), 
            .n32_adj_429(n32_adj_5598), .n32_adj_430(n32_adj_5534), .amdemod_d_11__N_2011(amdemod_d_11__N_2011), 
            .n47_adj_431(n47), .n47_adj_432(n47_adj_5966), .n47_adj_433(n47_adj_5602), 
            .n47_adj_434(n47_adj_5538), .n49_adj_435(n49_adj_5979), .n49_adj_436(n49_adj_6006), 
            .n49_adj_437(n49_adj_5474), .n49_adj_438(n49), .n44_adj_439(n44), 
            .n44_adj_440(n44_adj_5965), .amdemod_d_11__N_2008(amdemod_d_11__N_2008), 
            .amdemod_d_11__N_2017(amdemod_d_11__N_2017), .amdemod_d_11__N_2014(amdemod_d_11__N_2014)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(184[7] 189[6])
    CCU2C _add_1_1241_add_4_27 (.A0(phase_inc_gen[29]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[30]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15658), .COUT(n15659), .S0(n226), .S1(n223));
    defparam _add_1_1241_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1250_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15462), .S1(n71));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1250_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1250_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1250_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1250_add_4_1.INJECT1_1 = "NO";
    FD1S3AX rx_data_valid_40 (.D(rx_data_valid1), .CK(clk_80mhz), .Q(rx_data_valid));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam rx_data_valid_40.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i0 (.D(phase_inc_gen[0]), .CK(clk_80mhz), .Q(phase_inc_gen1[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i0.GSR = "ENABLED";
    CCU2C _add_1_1112_add_4_38 (.A0(integrator2[71]), .B0(integrator1[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15461), .S0(n78_adj_4984));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1112_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_36 (.A0(integrator2[69]), .B0(integrator1[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[70]), .B1(integrator1[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15460), .COUT(n15461), .S0(n84), 
          .S1(n81));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_34 (.A0(integrator2[67]), .B0(integrator1[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[68]), .B1(integrator1[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15459), .COUT(n15460), .S0(n90), 
          .S1(n87));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_34.INJECT1_1 = "NO";
    PLL PLL_inst (.clk_25mhz_c(clk_25mhz_c), .clk_80mhz(clk_80mhz), .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(102[9] 105[6])
    CCU2C _add_1_1115_add_4_36 (.A0(integrator_d_tmp[33]), .B0(integrator_tmp[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[34]), .B1(integrator_tmp[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15361), .COUT(n15362), .S0(comb6_71__N_1451[33]), 
          .S1(comb6_71__N_1451[34]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_32 (.A0(integrator2[65]), .B0(integrator1[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[66]), .B1(integrator1[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15458), .COUT(n15459), .S0(n96), 
          .S1(n93));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_4 (.A0(integrator1_adj_6020[2]), .B0(mix_cosinewave[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[3]), .B1(mix_cosinewave[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15320), .COUT(n15321), .S0(integrator1_71__N_418_adj_6036[2]), 
          .S1(integrator1_71__N_418_adj_6036[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_2 (.A0(integrator1_adj_6020[0]), .B0(mix_cosinewave[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[1]), .B1(mix_cosinewave[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15320), .S1(integrator1_71__N_418_adj_6036[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_993_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_28 (.A0(integrator_d_tmp[25]), .B0(integrator_tmp[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[26]), .B1(integrator_tmp[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15357), .COUT(n15358), .S0(comb6_71__N_1451[25]), 
          .S1(comb6_71__N_1451[26]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_24 (.A0(integrator4[22]), .B0(integrator3[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[23]), .B1(integrator3[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15398), .COUT(n15399), .S0(integrator4_71__N_634[22]), 
          .S1(integrator4_71__N_634[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_7 (.A0(integrator3_adj_6022[40]), .B0(cout_adj_5165), 
          .C0(n171_adj_5529), .D0(integrator4_adj_6023[40]), .A1(integrator3_adj_6022[41]), 
          .B1(cout_adj_5165), .C1(n168_adj_5528), .D1(integrator4_adj_6023[41]), 
          .CIN(n14993), .COUT(n14994), .S0(integrator4_71__N_634_adj_6039[40]), 
          .S1(integrator4_71__N_634_adj_6039[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_5 (.A0(integrator3_adj_6022[38]), .B0(cout_adj_5165), 
          .C0(n177_adj_5531), .D0(integrator4_adj_6023[38]), .A1(integrator3_adj_6022[39]), 
          .B1(cout_adj_5165), .C1(n174_adj_5530), .D1(integrator4_adj_6023[39]), 
          .CIN(n14992), .COUT(n14993), .S0(integrator4_71__N_634_adj_6039[38]), 
          .S1(integrator4_71__N_634_adj_6039[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_5.INJECT1_1 = "NO";
    FD1S3AX square_sum_e3__i1 (.D(n121), .CK(cic_sine_clk), .Q(square_sum[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i1.GSR = "ENABLED";
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    CCU2C _add_1_1241_add_4_25 (.A0(phase_inc_gen[27]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[28]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15657), .COUT(n15658), .S0(n232), .S1(n229));
    defparam _add_1_1241_add_4_25.INIT0 = 16'haaa0;
    defparam _add_1_1241_add_4_25.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_23 (.A0(phase_inc_gen[25]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[26]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15656), .COUT(n15657), .S0(n238), .S1(n235));
    defparam _add_1_1241_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_21 (.A0(phase_inc_gen[23]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[24]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15655), .COUT(n15656), .S0(n244), .S1(n241));
    defparam _add_1_1241_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_19 (.A0(phase_inc_gen[21]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[22]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15654), .COUT(n15655), .S0(n250), .S1(n247));
    defparam _add_1_1241_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_1241_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_17 (.A0(phase_inc_gen[19]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[20]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15653), .COUT(n15654), .S0(n256), .S1(n253));
    defparam _add_1_1241_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1241_add_4_17.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_15 (.A0(phase_inc_gen[17]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[18]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15652), .COUT(n15653), .S0(n262), .S1(n259));
    defparam _add_1_1241_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_15.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_13 (.A0(phase_inc_gen[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[16]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15651), .COUT(n15652), .S0(n268), .S1(n265));
    defparam _add_1_1241_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1241_add_4_13.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_11 (.A0(phase_inc_gen[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15650), .COUT(n15651), .S0(n274), .S1(n271));
    defparam _add_1_1241_add_4_11.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_9 (.A0(phase_inc_gen[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15649), .COUT(n15650), .S0(n280), .S1(n277));
    defparam _add_1_1241_add_4_9.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_7 (.A0(phase_inc_gen[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15648), .COUT(n15649), .S0(n286), .S1(n283));
    defparam _add_1_1241_add_4_7.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_18 (.A0(integrator2[51]), .B0(integrator1[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[52]), .B1(integrator1[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15451), .COUT(n15452), .S0(n138), 
          .S1(n135));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_5 (.A0(phase_inc_gen[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15647), .COUT(n15648), .S0(n292), .S1(n289));
    defparam _add_1_1241_add_4_5.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_3 (.A0(integrator3_adj_6022[36]), .B0(cout_adj_5165), 
          .C0(n183_adj_5533), .D0(integrator4_adj_6023[36]), .A1(integrator3_adj_6022[37]), 
          .B1(cout_adj_5165), .C1(n180_adj_5532), .D1(integrator4_adj_6023[37]), 
          .CIN(n14991), .COUT(n14992), .S0(integrator4_71__N_634_adj_6039[36]), 
          .S1(integrator4_71__N_634_adj_6039[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1187_add_4_4 (.A0(count_adj_6105[1]), .B0(data_in_reg[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(count_adj_6105[2]), .B1(data_in_reg[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15363), .COUT(n15364));
    defparam _add_1_1187_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1187_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1187_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1187_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_34 (.A0(integrator_d_tmp[31]), .B0(integrator_tmp[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[32]), .B1(integrator_tmp[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15360), .COUT(n15361), .S0(comb6_71__N_1451[31]), 
          .S1(comb6_71__N_1451[32]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_8 (.A0(integrator2[6]), .B0(integrator1[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[7]), .B1(integrator1[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15428), .COUT(n15429), .S0(integrator2_71__N_490[6]), 
          .S1(integrator2_71__N_490[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_2 (.A0(integrator2[0]), .B0(integrator1[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[1]), .B1(integrator1[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15426), .S1(integrator2_71__N_490[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_981_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_34 (.A0(integrator3[32]), .B0(integrator2[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[33]), .B1(integrator2[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15422), .COUT(n15423), .S0(integrator3_71__N_562[32]), 
          .S1(integrator3_71__N_562[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_32 (.A0(integrator3[30]), .B0(integrator2[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[31]), .B1(integrator2[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15421), .COUT(n15422), .S0(integrator3_71__N_562[30]), 
          .S1(integrator3_71__N_562[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_4 (.A0(integrator2[2]), .B0(integrator1[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[3]), .B1(integrator1[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15426), .COUT(n15427), .S0(integrator2_71__N_490[2]), 
          .S1(integrator2_71__N_490[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_6 (.A0(integrator2[4]), .B0(integrator1[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[5]), .B1(integrator1[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15427), .COUT(n15428), .S0(integrator2_71__N_490[4]), 
          .S1(integrator2_71__N_490[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15424), .S0(cout_adj_5073));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_984_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_984_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5165), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14991));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1097_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1097_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_3 (.A0(phase_inc_gen[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15646), .COUT(n15647), .S0(n298), .S1(n295));
    defparam _add_1_1241_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1241_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_28 (.A0(integrator3[26]), .B0(integrator2[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[27]), .B1(integrator2[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15419), .COUT(n15420), .S0(integrator3_71__N_562[26]), 
          .S1(integrator3_71__N_562[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_26 (.A0(integrator3[24]), .B0(integrator2[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[25]), .B1(integrator2[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15418), .COUT(n15419), .S0(integrator3_71__N_562[24]), 
          .S1(integrator3_71__N_562[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_24 (.A0(integrator3[22]), .B0(integrator2[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[23]), .B1(integrator2[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15417), .COUT(n15418), .S0(integrator3_71__N_562[22]), 
          .S1(integrator3_71__N_562[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_22 (.A0(integrator3[20]), .B0(integrator2[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[21]), .B1(integrator2[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15416), .COUT(n15417), .S0(integrator3_71__N_562[20]), 
          .S1(integrator3_71__N_562[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_20 (.A0(integrator3[18]), .B0(integrator2[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[19]), .B1(integrator2[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15415), .COUT(n15416), .S0(integrator3_71__N_562[18]), 
          .S1(integrator3_71__N_562[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_14 (.A0(integrator3[12]), .B0(integrator2[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[13]), .B1(integrator2[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15412), .COUT(n15413), .S0(integrator3_71__N_562[12]), 
          .S1(integrator3_71__N_562[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_6 (.A0(integrator3[4]), .B0(integrator2[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[5]), .B1(integrator2[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15408), .COUT(n15409), .S0(integrator3_71__N_562[4]), 
          .S1(integrator3_71__N_562[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_20 (.A0(integrator1_adj_6020[18]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[19]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15328), .COUT(n15329), .S0(integrator1_71__N_418_adj_6036[18]), 
          .S1(integrator1_71__N_418_adj_6036[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_12 (.A0(integrator3[10]), .B0(integrator2[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[11]), .B1(integrator2[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15411), .COUT(n15412), .S0(integrator3_71__N_562[10]), 
          .S1(integrator3_71__N_562[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_4 (.A0(integrator3[2]), .B0(integrator2[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[3]), .B1(integrator2[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15407), .COUT(n15408), .S0(integrator3_71__N_562[2]), 
          .S1(integrator3_71__N_562[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_18 (.A0(integrator3[16]), .B0(integrator2[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[17]), .B1(integrator2[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15414), .COUT(n15415), .S0(integrator3_71__N_562[16]), 
          .S1(integrator3_71__N_562[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_10 (.A0(integrator3[8]), .B0(integrator2[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[9]), .B1(integrator2[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15410), .COUT(n15411), .S0(integrator3_71__N_562[8]), 
          .S1(integrator3_71__N_562[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_2 (.A0(integrator3[0]), .B0(integrator2[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[1]), .B1(integrator2[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15407), .S1(integrator3_71__N_562[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_984_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_16 (.A0(integrator3[14]), .B0(integrator2[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[15]), .B1(integrator2[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15413), .COUT(n15414), .S0(integrator3_71__N_562[14]), 
          .S1(integrator3_71__N_562[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_8 (.A0(integrator3[6]), .B0(integrator2[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[7]), .B1(integrator2[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15409), .COUT(n15410), .S0(integrator3_71__N_562[6]), 
          .S1(integrator3_71__N_562[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_16 (.A0(integrator_d_tmp[13]), .B0(integrator_tmp[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[14]), .B1(integrator_tmp[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15351), .COUT(n15352), .S0(comb6_71__N_1451[13]), 
          .S1(comb6_71__N_1451[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_16.INJECT1_1 = "NO";
    FD1S3AX rx_byte_i8 (.D(rx_byte1[7]), .CK(clk_80mhz), .Q(led_c_7));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam rx_byte_i8.GSR = "ENABLED";
    CCU2C _add_1_993_add_4_18 (.A0(integrator1_adj_6020[16]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[17]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15327), .COUT(n15328), .S0(integrator1_71__N_418_adj_6036[16]), 
          .S1(integrator1_71__N_418_adj_6036[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_18.INJECT1_1 = "NO";
    FD1S3AX rx_byte_i7 (.D(rx_byte1[6]), .CK(clk_80mhz), .Q(led_c_6));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam rx_byte_i7.GSR = "ENABLED";
    FD1S3AX rx_byte_i6 (.D(rx_byte1[5]), .CK(clk_80mhz), .Q(led_c_5));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam rx_byte_i6.GSR = "ENABLED";
    FD1S3AX rx_byte_i5 (.D(rx_byte1[4]), .CK(clk_80mhz), .Q(led_c_4));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam rx_byte_i5.GSR = "ENABLED";
    FD1S3AX rx_byte_i4 (.D(rx_byte1[3]), .CK(clk_80mhz), .Q(led_c_3));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam rx_byte_i4.GSR = "ENABLED";
    FD1S3AX rx_byte_i3 (.D(rx_byte1[2]), .CK(clk_80mhz), .Q(led_c_2));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam rx_byte_i3.GSR = "ENABLED";
    FD1S3AX rx_byte_i2 (.D(rx_byte1[1]), .CK(clk_80mhz), .Q(led_c_1));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam rx_byte_i2.GSR = "ENABLED";
    CCU2C _add_1_993_add_4_16 (.A0(integrator1_adj_6020[14]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[15]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15326), .COUT(n15327), .S0(integrator1_71__N_418_adj_6036[14]), 
          .S1(integrator1_71__N_418_adj_6036[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_14 (.A0(integrator1_adj_6020[12]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[13]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15325), .COUT(n15326), .S0(integrator1_71__N_418_adj_6036[12]), 
          .S1(integrator1_71__N_418_adj_6036[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_12 (.A0(integrator1_adj_6020[10]), .B0(mix_cosinewave[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[11]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15324), .COUT(n15325), .S0(integrator1_71__N_418_adj_6036[10]), 
          .S1(integrator1_71__N_418_adj_6036[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_10 (.A0(integrator1_adj_6020[8]), .B0(mix_cosinewave[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[9]), .B1(mix_cosinewave[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15323), .COUT(n15324), .S0(integrator1_71__N_418_adj_6036[8]), 
          .S1(integrator1_71__N_418_adj_6036[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_8 (.A0(integrator1_adj_6020[6]), .B0(mix_cosinewave[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[7]), .B1(mix_cosinewave[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15322), .COUT(n15323), .S0(integrator1_71__N_418_adj_6036[6]), 
          .S1(integrator1_71__N_418_adj_6036[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_8.INJECT1_1 = "NO";
    FD1P3AX phase_inc_gen_i0_i1 (.D(n320), .SP(clk_80mhz_enable_1447), .CK(clk_80mhz), 
            .Q(phase_inc_gen[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i1.GSR = "ENABLED";
    CCU2C _add_1_996_add_4_13 (.A0(count[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15318), .S0(n28_adj_5077));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_996_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_996_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_996_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_996_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_996_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15317), .COUT(n15318), .S0(n34_adj_5079), 
          .S1(n31_adj_5078));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_996_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_996_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_996_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_996_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_22 (.A0(integrator2[55]), .B0(integrator1[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[56]), .B1(integrator1[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15453), .COUT(n15454), .S0(n126), 
          .S1(n123));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_22 (.A0(integrator4[20]), .B0(integrator3[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[21]), .B1(integrator3[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15397), .COUT(n15398), .S0(integrator4_71__N_634[20]), 
          .S1(integrator4_71__N_634[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_26 (.A0(integrator2[59]), .B0(integrator1[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[60]), .B1(integrator1[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15455), .COUT(n15456), .S0(n114), 
          .S1(n111));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_36 (.A0(integrator4[34]), .B0(integrator3[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[35]), .B1(integrator3[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15404), .COUT(n15405), .S0(integrator4_71__N_634[34]), 
          .S1(integrator4_71__N_634[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_34 (.A0(integrator4[32]), .B0(integrator3[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[33]), .B1(integrator3[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15403), .COUT(n15404), .S0(integrator4_71__N_634[32]), 
          .S1(integrator4_71__N_634[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_30 (.A0(integrator2[63]), .B0(integrator1[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[64]), .B1(integrator1[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15457), .COUT(n15458), .S0(n102), 
          .S1(n99));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_28 (.A0(integrator2[61]), .B0(integrator1[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[62]), .B1(integrator1[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15456), .COUT(n15457), .S0(n108), 
          .S1(n105));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_24 (.A0(integrator2[57]), .B0(integrator1[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[58]), .B1(integrator1[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15454), .COUT(n15455), .S0(n120), 
          .S1(n117));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_20 (.A0(integrator2[53]), .B0(integrator1[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[54]), .B1(integrator1[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15452), .COUT(n15453), .S0(n132), 
          .S1(n129));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_30 (.A0(integrator4[28]), .B0(integrator3[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[29]), .B1(integrator3[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15401), .COUT(n15402), .S0(integrator4_71__N_634[28]), 
          .S1(integrator4_71__N_634[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_32 (.A0(integrator4[30]), .B0(integrator3[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[31]), .B1(integrator3[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15402), .COUT(n15403), .S0(integrator4_71__N_634[30]), 
          .S1(integrator4_71__N_634[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_32.INJECT1_1 = "NO";
    OB pwm_out_p1_pad (.I(pwm_out_p4_c), .O(pwm_out_p1));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(45[23:33])
    CCU2C _add_1_987_add_4_20 (.A0(integrator4[18]), .B0(integrator3[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[19]), .B1(integrator3[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15396), .COUT(n15397), .S0(integrator4_71__N_634[18]), 
          .S1(integrator4_71__N_634[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_20.INJECT1_1 = "NO";
    OB pwm_out_p2_pad (.I(pwm_out_p4_c), .O(pwm_out_p2));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(46[23:33])
    CCU2C _add_1_987_add_4_28 (.A0(integrator4[26]), .B0(integrator3[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[27]), .B1(integrator3[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15400), .COUT(n15401), .S0(integrator4_71__N_634[26]), 
          .S1(integrator4_71__N_634[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_12 (.A0(integrator_d_tmp[9]), .B0(integrator_tmp[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[10]), .B1(integrator_tmp[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15349), .COUT(n15350), .S0(comb6_71__N_1451[9]), 
          .S1(comb6_71__N_1451[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_12 (.A0(integrator4[10]), .B0(integrator3[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[11]), .B1(integrator3[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15392), .COUT(n15393), .S0(integrator4_71__N_634[10]), 
          .S1(integrator4_71__N_634[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_996_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15316), .COUT(n15317), .S0(n40_adj_5081), .S1(n37_adj_5080));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_996_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_996_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_996_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_996_add_4_9.INJECT1_1 = "NO";
    FD1S3AX square_sum_e1_i0_i0 (.D(n80), .CK(cic_sine_clk), .Q(n48_adj_5701));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i0.GSR = "ENABLED";
    CCU2C _add_1_1241_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_gen[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15646), .S1(n301));
    defparam _add_1_1241_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1241_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_1.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_28 (.A0(phase_inc_gen1[26]), .B0(phase_accum[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[27]), .B1(phase_accum[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15482), .COUT(n15483), .S0(n243), 
          .S1(n240));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_28.INIT0 = 16'h666a;
    defparam phase_accum_add_4_28.INIT1 = 16'h666a;
    defparam phase_accum_add_4_28.INJECT1_0 = "NO";
    defparam phase_accum_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_38 (.A0(comb_d9[71]), .B0(comb9[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15645), .S0(n78_adj_5889));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1154_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_26 (.A0(integrator4[24]), .B0(integrator3[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[25]), .B1(integrator3[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15399), .COUT(n15400), .S0(integrator4_71__N_634[24]), 
          .S1(integrator4_71__N_634[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_16 (.A0(integrator4[14]), .B0(integrator3[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[15]), .B1(integrator3[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15394), .COUT(n15395), .S0(integrator4_71__N_634[14]), 
          .S1(integrator4_71__N_634[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_6 (.A0(integrator4[4]), .B0(integrator3[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[5]), .B1(integrator3[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15389), .COUT(n15390), .S0(integrator4_71__N_634[4]), 
          .S1(integrator4_71__N_634[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_8 (.A0(integrator4[6]), .B0(integrator3[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[7]), .B1(integrator3[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15390), .COUT(n15391), .S0(integrator4_71__N_634[6]), 
          .S1(integrator4_71__N_634[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_18 (.A0(integrator4[16]), .B0(integrator3[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[17]), .B1(integrator3[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15395), .COUT(n15396), .S0(integrator4_71__N_634[16]), 
          .S1(integrator4_71__N_634[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_4 (.A0(integrator4[2]), .B0(integrator3[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[3]), .B1(integrator3[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15388), .COUT(n15389), .S0(integrator4_71__N_634[2]), 
          .S1(integrator4_71__N_634[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_14 (.A0(integrator4[12]), .B0(integrator3[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[13]), .B1(integrator3[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15393), .COUT(n15394), .S0(integrator4_71__N_634[12]), 
          .S1(integrator4_71__N_634[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_2 (.A0(integrator4[0]), .B0(integrator3[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[1]), .B1(integrator3[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15388), .S1(integrator4_71__N_634[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_987_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_16 (.A0(integrator2[49]), .B0(integrator1[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[50]), .B1(integrator1[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15450), .COUT(n15451), .S0(n144), 
          .S1(n141));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_14 (.A0(integrator2[47]), .B0(integrator1[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[48]), .B1(integrator1[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15449), .COUT(n15450), .S0(n150), 
          .S1(n147));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_6 (.A0(integrator2[39]), .B0(integrator1[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[40]), .B1(integrator1[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15445), .COUT(n15446), .S0(n174), 
          .S1(n171));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_4 (.A0(integrator2[37]), .B0(integrator1[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[38]), .B1(integrator1[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15444), .COUT(n15445), .S0(n180), 
          .S1(n177));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator2[36]), .B1(integrator1[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15444), .S1(n183));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1112_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15443), .S0(cout_adj_5072));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_981_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_981_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_12 (.A0(integrator2[45]), .B0(integrator1[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[46]), .B1(integrator1[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15448), .COUT(n15449), .S0(n156), 
          .S1(n153));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_10 (.A0(integrator2[43]), .B0(integrator1[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[44]), .B1(integrator1[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15447), .COUT(n15448), .S0(n162), 
          .S1(n159));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1112_add_4_8 (.A0(integrator2[41]), .B0(integrator1[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[42]), .B1(integrator1[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15446), .COUT(n15447), .S0(n168), 
          .S1(n165));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1112_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1112_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1112_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1112_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_32 (.A0(integrator2[30]), .B0(integrator1[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[31]), .B1(integrator1[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15440), .COUT(n15441), .S0(integrator2_71__N_490[30]), 
          .S1(integrator2_71__N_490[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_30 (.A0(integrator2[28]), .B0(integrator1[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[29]), .B1(integrator1[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15439), .COUT(n15440), .S0(integrator2_71__N_490[28]), 
          .S1(integrator2_71__N_490[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_28 (.A0(integrator2[26]), .B0(integrator1[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[27]), .B1(integrator1[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15438), .COUT(n15439), .S0(integrator2_71__N_490[26]), 
          .S1(integrator2_71__N_490[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_26 (.A0(integrator2[24]), .B0(integrator1[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[25]), .B1(integrator1[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15437), .COUT(n15438), .S0(integrator2_71__N_490[24]), 
          .S1(integrator2_71__N_490[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1196_add_4_16 (.A0(amdemod_d_11__N_2209), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14987), .S0(amdemod_d_11__N_1870[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1196_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1196_add_4_16.INIT1 = 16'h0000;
    defparam _add_1_1196_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1196_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1196_add_4_14 (.A0(amdemod_d_11__N_2215), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2212), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14986), .COUT(n14987), .S0(amdemod_d_11__N_1870[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1196_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_1196_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_1196_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1196_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1196_add_4_12 (.A0(n17137), .B0(amdemod_d_11__N_2221), 
          .C0(GND_net), .D0(VCC_net), .A1(square_sum[23]), .B1(square_sum[22]), 
          .C1(amdemod_d_11__N_2218), .D1(VCC_net), .CIN(n14985), .COUT(n14986), 
          .S0(amdemod_d_11__N_1870[9]), .S1(amdemod_d_11__N_1870[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1196_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1196_add_4_12.INIT1 = 16'he1e1;
    defparam _add_1_1196_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1196_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1196_add_4_10 (.A0(amdemod_d_11__N_2227), .B0(amdemod_d_11__N_1841[11]), 
          .C0(n17134), .D0(amdemod_d_11__N_1840[11]), .A1(n17134), .B1(amdemod_d_11__N_2224), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14984), .COUT(n14985), .S0(amdemod_d_11__N_1870[7]), 
          .S1(amdemod_d_11__N_1870[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1196_add_4_10.INIT0 = 16'h656a;
    defparam _add_1_1196_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1196_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1196_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1196_add_4_8 (.A0(amdemod_d_11__N_2233), .B0(amdemod_d_11__N_1851[13]), 
          .C0(n17132), .D0(amdemod_d_11__N_1850[13]), .A1(n17132), .B1(amdemod_d_11__N_2230), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14983), .COUT(n14984), .S0(amdemod_d_11__N_1870[5]), 
          .S1(amdemod_d_11__N_1870[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1196_add_4_8.INIT0 = 16'h656a;
    defparam _add_1_1196_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1196_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1196_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_30 (.A0(integrator3[28]), .B0(integrator2[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[29]), .B1(integrator2[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15420), .COUT(n15421), .S0(integrator3_71__N_562[28]), 
          .S1(integrator3_71__N_562[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1196_add_4_6 (.A0(amdemod_d_11__N_2239), .B0(amdemod_d_11__N_1861[13]), 
          .C0(n17130), .D0(amdemod_d_11__N_1860[13]), .A1(n17130), .B1(amdemod_d_11__N_2236), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14982), .COUT(n14983), .S0(amdemod_d_11__N_1870[3]), 
          .S1(amdemod_d_11__N_1870[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1196_add_4_6.INIT0 = 16'h656a;
    defparam _add_1_1196_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1196_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1196_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1196_add_4_4 (.A0(n17128), .B0(square_sum[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(n17128), .B1(amdemod_d_11__N_2242), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14981), .COUT(n14982), .S0(amdemod_d_11__N_1870[1]), 
          .S1(amdemod_d_11__N_1870[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1196_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1196_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1196_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1196_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1196_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14981), .S1(amdemod_d_11__N_1870[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1196_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1196_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1196_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1196_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_37 (.A0(comb8_adj_6029[70]), .B0(cout_adj_5310), 
          .C0(n81_adj_5625), .D0(n3_adj_4947), .A1(comb8_adj_6029[71]), 
          .B1(cout_adj_5310), .C1(n78_adj_5624), .D1(n2_adj_4946), .CIN(n14979), 
          .S0(comb9_71__N_1667_adj_6055[70]), .S1(comb9_71__N_1667_adj_6055[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_35 (.A0(comb8_adj_6029[68]), .B0(cout_adj_5310), 
          .C0(n87_adj_5627), .D0(n5_adj_4949), .A1(comb8_adj_6029[69]), 
          .B1(cout_adj_5310), .C1(n84_adj_5626), .D1(n4_adj_4948), .CIN(n14978), 
          .COUT(n14979), .S0(comb9_71__N_1667_adj_6055[68]), .S1(comb9_71__N_1667_adj_6055[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_33 (.A0(comb8_adj_6029[66]), .B0(cout_adj_5310), 
          .C0(n93_adj_5629), .D0(n7_adj_4951), .A1(comb8_adj_6029[67]), 
          .B1(cout_adj_5310), .C1(n90_adj_5628), .D1(n6_adj_4950), .CIN(n14977), 
          .COUT(n14978), .S0(comb9_71__N_1667_adj_6055[66]), .S1(comb9_71__N_1667_adj_6055[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_31 (.A0(comb8_adj_6029[64]), .B0(cout_adj_5310), 
          .C0(n99_adj_5631), .D0(n9_adj_4953), .A1(comb8_adj_6029[65]), 
          .B1(cout_adj_5310), .C1(n96_adj_5630), .D1(n8_adj_4952), .CIN(n14976), 
          .COUT(n14977), .S0(comb9_71__N_1667_adj_6055[64]), .S1(comb9_71__N_1667_adj_6055[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_24 (.A0(integrator2[22]), .B0(integrator1[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[23]), .B1(integrator1[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15436), .COUT(n15437), .S0(integrator2_71__N_490[22]), 
          .S1(integrator2_71__N_490[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_32 (.A0(integrator5[30]), .B0(integrator4[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[31]), .B1(integrator4[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15383), .COUT(n15384), .S0(integrator5_71__N_706[30]), 
          .S1(integrator5_71__N_706[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_26 (.A0(integrator5[24]), .B0(integrator4[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[25]), .B1(integrator4[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15380), .COUT(n15381), .S0(integrator5_71__N_706[24]), 
          .S1(integrator5_71__N_706[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_20 (.A0(integrator5[18]), .B0(integrator4[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[19]), .B1(integrator4[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15377), .COUT(n15378), .S0(integrator5_71__N_706[18]), 
          .S1(integrator5_71__N_706[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_24 (.A0(integrator5[22]), .B0(integrator4[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[23]), .B1(integrator4[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15379), .COUT(n15380), .S0(integrator5_71__N_706[22]), 
          .S1(integrator5_71__N_706[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_30 (.A0(integrator5[28]), .B0(integrator4[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[29]), .B1(integrator4[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15382), .COUT(n15383), .S0(integrator5_71__N_706[28]), 
          .S1(integrator5_71__N_706[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_22 (.A0(integrator5[20]), .B0(integrator4[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[21]), .B1(integrator4[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15378), .COUT(n15379), .S0(integrator5_71__N_706[20]), 
          .S1(integrator5_71__N_706[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_18 (.A0(integrator5[16]), .B0(integrator4[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[17]), .B1(integrator4[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15376), .COUT(n15377), .S0(integrator5_71__N_706[16]), 
          .S1(integrator5_71__N_706[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_28 (.A0(integrator5[26]), .B0(integrator4[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[27]), .B1(integrator4[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15381), .COUT(n15382), .S0(integrator5_71__N_706[26]), 
          .S1(integrator5_71__N_706[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_16 (.A0(integrator5[14]), .B0(integrator4[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[15]), .B1(integrator4[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15375), .COUT(n15376), .S0(integrator5_71__N_706[14]), 
          .S1(integrator5_71__N_706[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_36 (.A0(integrator5[34]), .B0(integrator4[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[35]), .B1(integrator4[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15385), .COUT(n15386), .S0(integrator5_71__N_706[34]), 
          .S1(integrator5_71__N_706[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_14 (.A0(integrator5[12]), .B0(integrator4[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[13]), .B1(integrator4[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15374), .COUT(n15375), .S0(integrator5_71__N_706[12]), 
          .S1(integrator5_71__N_706[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_8 (.A0(integrator5[6]), .B0(integrator4[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[7]), .B1(integrator4[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15371), .COUT(n15372), .S0(integrator5_71__N_706[6]), 
          .S1(integrator5_71__N_706[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_6 (.A0(integrator5[4]), .B0(integrator4[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[5]), .B1(integrator4[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15370), .COUT(n15371), .S0(integrator5_71__N_706[4]), 
          .S1(integrator5_71__N_706[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1187_add_4_12 (.A0(count_adj_6105[9]), .B0(data_in_reg[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15367), .S1(cout_adj_5347));
    defparam _add_1_1187_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1187_add_4_12.INIT1 = 16'h0000;
    defparam _add_1_1187_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1187_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_12 (.A0(integrator5[10]), .B0(integrator4[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[11]), .B1(integrator4[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15373), .COUT(n15374), .S0(integrator5_71__N_706[10]), 
          .S1(integrator5_71__N_706[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_4 (.A0(integrator5[2]), .B0(integrator4[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[3]), .B1(integrator4[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15369), .COUT(n15370), .S0(integrator5_71__N_706[2]), 
          .S1(integrator5_71__N_706[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1187_add_4_10 (.A0(count_adj_6105[7]), .B0(data_in_reg[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(count_adj_6105[8]), .B1(data_in_reg[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15366), .COUT(n15367));
    defparam _add_1_1187_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1187_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1187_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1187_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_10 (.A0(integrator5[8]), .B0(integrator4[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[9]), .B1(integrator4[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15372), .COUT(n15373), .S0(integrator5_71__N_706[8]), 
          .S1(integrator5_71__N_706[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_2 (.A0(integrator5[0]), .B0(integrator4[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[1]), .B1(integrator4[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15369), .S1(integrator5_71__N_706[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_990_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1187_add_4_8 (.A0(count_adj_6105[5]), .B0(data_in_reg[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(count_adj_6105[6]), .B1(data_in_reg[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15365), .COUT(n15366));
    defparam _add_1_1187_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1187_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1187_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1187_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1187_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_6105[0]), .B1(data_in_reg[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15363));
    defparam _add_1_1187_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1187_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1187_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1187_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_32 (.A0(integrator_d_tmp[29]), .B0(integrator_tmp[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[30]), .B1(integrator_tmp[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15359), .COUT(n15360), .S0(comb6_71__N_1451[29]), 
          .S1(comb6_71__N_1451[30]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_38 (.A0(integrator_d_tmp[35]), .B0(integrator_tmp[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15362), .S0(comb6_71__N_1451[35]), .S1(cout));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1115_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_30 (.A0(integrator_d_tmp[27]), .B0(integrator_tmp[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[28]), .B1(integrator_tmp[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15358), .COUT(n15359), .S0(comb6_71__N_1451[27]), 
          .S1(comb6_71__N_1451[28]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1187_add_4_6 (.A0(count_adj_6105[3]), .B0(data_in_reg[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(count_adj_6105[4]), .B1(data_in_reg[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15364), .COUT(n15365));
    defparam _add_1_1187_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1187_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1187_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1187_add_4_6.INJECT1_1 = "NO";
    LUT4 mux_251_i47_4_lut (.A(n11373), .B(n181_adj_5921), .C(n17136), 
         .D(n2244), .Z(n1998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i47_4_lut.init = 16'hcfca;
    CCU2C _add_1_987_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15405), .S0(cout_adj_5074));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_987_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_987_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_cout.INJECT1_1 = "NO";
    LUT4 mux_251_i2_4_lut_then_4_lut (.A(led_c_3), .B(n17150), .C(n16220), 
         .D(led_c_4), .Z(n17173)) /* synthesis lut_function=(!(A+!(B (C (D))+!B ((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i2_4_lut_then_4_lut.init = 16'h5101;
    LUT4 mux_251_i2_4_lut_else_4_lut (.A(led_c_3), .B(n17150), .C(n16220), 
         .Z(n17172)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i2_4_lut_else_4_lut.init = 16'h0101;
    CCU2C _add_1_1115_add_4_26 (.A0(integrator_d_tmp[23]), .B0(integrator_tmp[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[24]), .B1(integrator_tmp[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15356), .COUT(n15357), .S0(comb6_71__N_1451[23]), 
          .S1(comb6_71__N_1451[24]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_24 (.A0(integrator_d_tmp[21]), .B0(integrator_tmp[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[22]), .B1(integrator_tmp[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15355), .COUT(n15356), .S0(comb6_71__N_1451[21]), 
          .S1(comb6_71__N_1451[22]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_24.INJECT1_1 = "NO";
    LUT4 led_c_3_bdd_4_lut (.A(led_c_3), .B(n313), .C(n16220), .D(led_c_4), 
         .Z(n17175)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !(C)))) */ ;
    defparam led_c_3_bdd_4_lut.init = 16'h4505;
    LUT4 mux_251_i4_4_lut_4_lut_4_lut_then_3_lut (.A(led_c_3), .B(n310), 
         .C(led_c_4), .Z(n17177)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam mux_251_i4_4_lut_4_lut_4_lut_then_3_lut.init = 16'h4545;
    LUT4 i2403_2_lut_rep_350 (.A(led_c_4), .B(n1827), .Z(n17147)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i2403_2_lut_rep_350.init = 16'h8888;
    LUT4 mux_251_i48_4_lut (.A(n11375), .B(n178_adj_5920), .C(n17136), 
         .D(n2244), .Z(n1997)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i48_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1115_add_4_22 (.A0(integrator_d_tmp[19]), .B0(integrator_tmp[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[20]), .B1(integrator_tmp[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15354), .COUT(n15355), .S0(comb6_71__N_1451[19]), 
          .S1(comb6_71__N_1451[20]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_22.INJECT1_1 = "NO";
    LUT4 i2567_1_lut_2_lut (.A(led_c_4), .B(n1827), .Z(n2579)) /* synthesis lut_function=(!(A (B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i2567_1_lut_2_lut.init = 16'h7777;
    CCU2C _add_1_1115_add_4_20 (.A0(integrator_d_tmp[17]), .B0(integrator_tmp[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[18]), .B1(integrator_tmp[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15353), .COUT(n15354), .S0(comb6_71__N_1451[17]), 
          .S1(comb6_71__N_1451[18]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_20.INJECT1_1 = "NO";
    LUT4 mux_366_i3_3_lut_rep_351 (.A(led_c_2), .B(led_c_4), .C(n1827), 
         .Z(n17148)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_366_i3_3_lut_rep_351.init = 16'hcaca;
    LUT4 i1456_1_lut_3_lut (.A(led_c_2), .B(led_c_4), .C(n1827), .Z(n11169)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1456_1_lut_3_lut.init = 16'h3535;
    LUT4 mux_251_i4_4_lut_4_lut_4_lut_else_3_lut (.A(led_c_3), .B(n17150), 
         .C(led_c_2), .Z(n17176)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam mux_251_i4_4_lut_4_lut_4_lut_else_3_lut.init = 16'h4040;
    LUT4 mux_251_i45_4_lut (.A(n2065), .B(n187_adj_5923), .C(n17136), 
         .D(n11259), .Z(n2000)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i45_4_lut.init = 16'hc0ca;
    LUT4 mux_251_i46_4_lut (.A(n11371), .B(n184_adj_5922), .C(n17136), 
         .D(n2244), .Z(n1999)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i46_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut_2_lut_rep_367 (.A(n16203), .B(n16409), .Z(n17278)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_4_lut_2_lut_rep_367.init = 16'h8888;
    LUT4 mux_251_i43_4_lut (.A(n11367), .B(n193_adj_5925), .C(n17136), 
         .D(n2244), .Z(n2002)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i43_4_lut.init = 16'hc0ca;
    LUT4 i1_3_lut_4_lut (.A(led_c_4), .B(n17155), .C(led_c_6), .D(n16245), 
         .Z(n11789)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff7f;
    LUT4 mux_251_i44_4_lut (.A(n11369), .B(n190_adj_5924), .C(n17136), 
         .D(n2244), .Z(n2001)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i44_4_lut.init = 16'hc0ca;
    LUT4 i4727_4_lut_rep_418 (.A(n16451), .B(n17153), .C(n17049), .D(n16957), 
         .Z(n17335)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C))) */ ;
    defparam i4727_4_lut_rep_418.init = 16'hc0c8;
    CCU2C _add_1_981_add_4_36 (.A0(integrator2[34]), .B0(integrator1[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[35]), .B1(integrator1[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15442), .COUT(n15443), .S0(integrator2_71__N_490[34]), 
          .S1(integrator2_71__N_490[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_34 (.A0(integrator2[32]), .B0(integrator1[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[33]), .B1(integrator1[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15441), .COUT(n15442), .S0(integrator2_71__N_490[32]), 
          .S1(integrator2_71__N_490[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_34.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_352_3_lut (.A(led_c_6), .B(n17155), .C(led_c_4), 
         .Z(n17149)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i1_2_lut_rep_352_3_lut.init = 16'hf7f7;
    LUT4 i4727_4_lut_rep_419 (.A(n16451), .B(n17153), .C(n17049), .D(n16957), 
         .Z(clk_80mhz_enable_1497)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C))) */ ;
    defparam i4727_4_lut_rep_419.init = 16'hc0c8;
    LUT4 i5754_3_lut_4_lut (.A(led_c_6), .B(n17155), .C(led_c_4), .D(n29_adj_6001), 
         .Z(n16348)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i5754_3_lut_4_lut.init = 16'hf7ff;
    LUT4 i26_4_lut (.A(n2244), .B(n199_adj_5927), .C(n17136), .D(n13_adj_5726), 
         .Z(n11_adj_5725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i26_4_lut.init = 16'hcacf;
    LUT4 i1880_4_lut (.A(n196_adj_5926), .B(n190), .C(led_c_3), .D(n17144), 
         .Z(n11614)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1880_4_lut.init = 16'hcac0;
    LUT4 mux_251_i39_4_lut (.A(n11361), .B(n205_adj_5929), .C(n17136), 
         .D(n2244), .Z(n2006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i39_4_lut.init = 16'hcfca;
    LUT4 i1_3_lut_rep_358 (.A(led_c_5), .B(led_c_7), .C(rx_data_valid), 
         .Z(n17155)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i1_3_lut_rep_358.init = 16'h2020;
    CCU2C _add_1_981_add_4_22 (.A0(integrator2[20]), .B0(integrator1[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[21]), .B1(integrator1[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15435), .COUT(n15436), .S0(integrator2_71__N_490[20]), 
          .S1(integrator2_71__N_490[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_22.INJECT1_1 = "NO";
    FD1S3AX phase_accum_e3_i0_i0 (.D(n321), .CK(clk_80mhz), .Q(phase_accum[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i0.GSR = "ENABLED";
    LUT4 mux_251_i40_4_lut (.A(n11363), .B(n202_adj_5928), .C(n17136), 
         .D(n2244), .Z(n2005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i40_4_lut.init = 16'hcfca;
    LUT4 mux_251_i37_4_lut (.A(n11357), .B(n211_adj_5931), .C(n17136), 
         .D(n2244), .Z(n2008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i37_4_lut.init = 16'hcfca;
    LUT4 i4723_2_lut_rep_355_4_lut (.A(led_c_5), .B(led_c_7), .C(rx_data_valid), 
         .D(led_c_4), .Z(n17152)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i4723_2_lut_rep_355_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_rep_356_4_lut (.A(led_c_5), .B(led_c_7), .C(rx_data_valid), 
         .D(led_c_6), .Z(n17153)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i1_2_lut_rep_356_4_lut.init = 16'h2000;
    LUT4 i5729_3_lut_4_lut (.A(n16203), .B(n16409), .C(n17335), .D(led_c_3), 
         .Z(clk_80mhz_enable_1447)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam i5729_3_lut_4_lut.init = 16'h80f0;
    LUT4 mux_251_i38_4_lut (.A(n11359), .B(n208_adj_5930), .C(n17136), 
         .D(n2244), .Z(n2007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i38_4_lut.init = 16'hcfca;
    LUT4 i45_4_lut_4_lut_4_lut (.A(led_c_3), .B(led_c_0), .C(led_c_1), 
         .D(n17288), .Z(n29_adj_6001)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i45_4_lut_4_lut_4_lut.init = 16'h6014;
    LUT4 i2405_2_lut (.A(led_c_4), .B(n1827), .Z(n2580)) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i2405_2_lut.init = 16'hbbbb;
    LUT4 mux_251_i35_4_lut (.A(n11353), .B(n217_adj_5933), .C(n17136), 
         .D(n2244), .Z(n2010)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i35_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1154_add_4_36 (.A0(comb_d9[69]), .B0(comb9[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[70]), .B1(comb9[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15644), .COUT(n15645), .S0(n84_adj_5891), 
          .S1(n81_adj_5890));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_36.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_361 (.A(led_c_1), .B(led_c_4), .Z(n17158)) /* synthesis lut_function=(!((B)+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i1_2_lut_rep_361.init = 16'h2222;
    LUT4 n17048_bdd_2_lut (.A(n17048), .B(led_c_4), .Z(n17049)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n17048_bdd_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut (.A(led_c_3), .B(led_c_0), .C(led_c_4), 
         .D(led_c_1), .Z(n16238)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(247[13] 258[20])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 led_c_4_bdd_4_lut (.A(n17288), .B(led_c_0), .C(led_c_3), .D(led_c_1), 
         .Z(n17048)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !(B+(C (D)+!C !(D)))) */ ;
    defparam led_c_4_bdd_4_lut.init = 16'hab90;
    LUT4 mux_251_i36_4_lut (.A(n11355), .B(n214_adj_5932), .C(n17136), 
         .D(n2244), .Z(n2009)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i36_4_lut.init = 16'hc0ca;
    LUT4 i1659_3_lut_4_lut (.A(n17288), .B(n17150), .C(led_c_3), .D(n160), 
         .Z(n11381)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1659_3_lut_4_lut.init = 16'hf404;
    OB pwm_out_pad (.I(pwm_out_p4_c), .O(pwm_out));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(44[23:30])
    LUT4 mux_251_i33_4_lut (.A(n11349), .B(n223_adj_5935), .C(n17136), 
         .D(n2244), .Z(n2012)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i33_4_lut.init = 16'hc0ca;
    CCU2C _add_1_981_add_4_20 (.A0(integrator2[18]), .B0(integrator1[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[19]), .B1(integrator1[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15434), .COUT(n15435), .S0(integrator2_71__N_490[18]), 
          .S1(integrator2_71__N_490[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_20.INJECT1_1 = "NO";
    LUT4 mux_251_i34_4_lut (.A(n11351), .B(n220_adj_5934), .C(n17136), 
         .D(n2244), .Z(n2011)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i34_4_lut.init = 16'hcfca;
    LUT4 i1649_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(n17289), .D(n178), 
         .Z(n11371)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1649_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_251_i31_4_lut (.A(n11345), .B(n229_adj_5937), .C(n17136), 
         .D(n2244), .Z(n2014)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i31_4_lut.init = 16'hc0ca;
    LUT4 i1639_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(led_c_3), .D(n199), 
         .Z(n11361)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1639_3_lut_4_lut.init = 16'hf404;
    CCU2C _add_1_996_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15315), .COUT(n15316), .S0(n46_adj_5083), .S1(n43_adj_5082));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_996_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_996_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_996_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_996_add_4_7.INJECT1_1 = "NO";
    LUT4 mux_251_i32_4_lut (.A(n11347), .B(n226_adj_5936), .C(n17136), 
         .D(n2244), .Z(n2013)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i32_4_lut.init = 16'hc0ca;
    LUT4 i1641_3_lut_4_lut (.A(n17288), .B(n17150), .C(n17289), .D(n196), 
         .Z(n11363)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1641_3_lut_4_lut.init = 16'hf404;
    CCU2C _add_1_1088_add_4_29 (.A0(comb8_adj_6029[62]), .B0(cout_adj_5310), 
          .C0(n105_adj_5633), .D0(n11_adj_4955), .A1(comb8_adj_6029[63]), 
          .B1(cout_adj_5310), .C1(n102_adj_5632), .D1(n10_adj_4954), .CIN(n14975), 
          .COUT(n14976), .S0(comb9_71__N_1667_adj_6055[62]), .S1(comb9_71__N_1667_adj_6055[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_29.INJECT1_1 = "NO";
    LUT4 n16254_bdd_4_lut (.A(n17139), .B(led_c_0), .C(led_c_3), .D(n17288), 
         .Z(n17043)) /* synthesis lut_function=(A+(B+!(C (D)+!C !(D)))) */ ;
    defparam n16254_bdd_4_lut.init = 16'heffe;
    LUT4 mux_366_i2_3_lut (.A(led_c_2), .B(led_c_4), .C(n1827), .Z(n2594)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_366_i2_3_lut.init = 16'hc5c5;
    LUT4 mux_251_i29_4_lut (.A(n11341), .B(n235_adj_5939), .C(n17136), 
         .D(n2244), .Z(n2016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i29_4_lut.init = 16'hcfca;
    LUT4 i1635_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(n17289), .D(n205), 
         .Z(n11357)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1635_3_lut_4_lut.init = 16'hf404;
    LUT4 i1633_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(led_c_3), .D(n208), 
         .Z(n11355)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1633_3_lut_4_lut.init = 16'hf404;
    CCU2C _add_1_1088_add_4_27 (.A0(comb8_adj_6029[60]), .B0(cout_adj_5310), 
          .C0(n111_adj_5635), .D0(n13_adj_4957), .A1(comb8_adj_6029[61]), 
          .B1(cout_adj_5310), .C1(n108_adj_5634), .D1(n12_adj_4956), .CIN(n14974), 
          .COUT(n14975), .S0(comb9_71__N_1667_adj_6055[60]), .S1(comb9_71__N_1667_adj_6055[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_25 (.A0(comb8_adj_6029[58]), .B0(cout_adj_5310), 
          .C0(n117_adj_5637), .D0(n15_adj_4959), .A1(comb8_adj_6029[59]), 
          .B1(cout_adj_5310), .C1(n114_adj_5636), .D1(n14_adj_4958), .CIN(n14973), 
          .COUT(n14974), .S0(comb9_71__N_1667_adj_6055[58]), .S1(comb9_71__N_1667_adj_6055[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_25.INJECT1_1 = "NO";
    LUT4 i1625_3_lut_4_lut (.A(n17288), .B(n17150), .C(n17289), .D(n220), 
         .Z(n11347)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1625_3_lut_4_lut.init = 16'hf404;
    LUT4 i1619_3_lut_4_lut (.A(n17288), .B(n17150), .C(n17289), .D(n229), 
         .Z(n11341)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1619_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_251_i30_4_lut (.A(n2214), .B(n232_adj_5938), .C(n17136), 
         .D(n2244), .Z(n2015)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i30_4_lut.init = 16'hc0ca;
    CCU2C _add_1_981_add_4_18 (.A0(integrator2[16]), .B0(integrator1[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[17]), .B1(integrator1[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15433), .COUT(n15434), .S0(integrator2_71__N_490[16]), 
          .S1(integrator2_71__N_490[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_18.INJECT1_1 = "NO";
    LUT4 i1609_3_lut_4_lut (.A(n17288), .B(n17150), .C(n17289), .D(n244), 
         .Z(n11331)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1609_3_lut_4_lut.init = 16'hf404;
    CCU2C add_3221_13 (.A0(square_sum[23]), .B0(square_sum[22]), .C0(amdemod_d_11__N_2284), 
          .D0(VCC_net), .A1(amdemod_d_11__N_2281), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15849), .S1(amdemod_d_11__N_1881[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam add_3221_13.INIT0 = 16'h1e1e;
    defparam add_3221_13.INIT1 = 16'haaa0;
    defparam add_3221_13.INJECT1_0 = "NO";
    defparam add_3221_13.INJECT1_1 = "NO";
    FD1P3AX cic_gain__i1 (.D(led_c_0), .SP(clk_80mhz_enable_1445), .CK(clk_80mhz), 
            .Q(cic_gain[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam cic_gain__i1.GSR = "ENABLED";
    CCU2C add_3221_11 (.A0(n17134), .B0(amdemod_d_11__N_2290), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_d_11__N_2287), .B1(n17162), .C1(n17279), 
          .D1(n17146), .CIN(n15848), .COUT(n15849));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam add_3221_11.INIT0 = 16'h9995;
    defparam add_3221_11.INIT1 = 16'h596a;
    defparam add_3221_11.INJECT1_0 = "NO";
    defparam add_3221_11.INJECT1_1 = "NO";
    CCU2C add_3221_9 (.A0(n17132), .B0(amdemod_d_11__N_2296), .C0(GND_net), 
          .D0(VCC_net), .A1(n17133), .B1(amdemod_d_11__N_2293), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15847), .COUT(n15848));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam add_3221_9.INIT0 = 16'h9995;
    defparam add_3221_9.INIT1 = 16'h9995;
    defparam add_3221_9.INJECT1_0 = "NO";
    defparam add_3221_9.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_16 (.A0(integrator2[14]), .B0(integrator1[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[15]), .B1(integrator1[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15432), .COUT(n15433), .S0(integrator2_71__N_490[14]), 
          .S1(integrator2_71__N_490[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_14 (.A0(integrator2[12]), .B0(integrator1[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[13]), .B1(integrator1[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15431), .COUT(n15432), .S0(integrator2_71__N_490[12]), 
          .S1(integrator2_71__N_490[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_12 (.A0(integrator2[10]), .B0(integrator1[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[11]), .B1(integrator1[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15430), .COUT(n15431), .S0(integrator2_71__N_490[10]), 
          .S1(integrator2_71__N_490[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_12.INJECT1_1 = "NO";
    OB diff_out_pad (.I(diff_out_c), .O(diff_out));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(43[23:31])
    FD1S3AX _add_1_1187_i7 (.D(cout_adj_5347), .CK(clk_80mhz), .Q(pwm_out_p4_c));
    defparam _add_1_1187_i7.GSR = "ENABLED";
    CCU2C add_3221_7 (.A0(n17130), .B0(amdemod_d_11__N_2302), .C0(GND_net), 
          .D0(VCC_net), .A1(n17131), .B1(amdemod_d_11__N_2299), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15846), .COUT(n15847));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam add_3221_7.INIT0 = 16'h9995;
    defparam add_3221_7.INIT1 = 16'h9995;
    defparam add_3221_7.INJECT1_0 = "NO";
    defparam add_3221_7.INJECT1_1 = "NO";
    CCU2C _add_1_984_add_4_36 (.A0(integrator3[34]), .B0(integrator2[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[35]), .B1(integrator2[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15423), .COUT(n15424), .S0(integrator3_71__N_562[34]), 
          .S1(integrator3_71__N_562[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_984_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_984_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_984_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_984_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_996_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15314), .COUT(n15315), .S0(n52_adj_5085), .S1(n49_adj_5084));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_996_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_996_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_996_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_996_add_4_5.INJECT1_1 = "NO";
    LUT4 i1597_3_lut_4_lut (.A(n17288), .B(n17150), .C(led_c_3), .D(n265), 
         .Z(n11319)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1597_3_lut_4_lut.init = 16'hf404;
    CCU2C _add_1_996_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n15313), .COUT(n15314), .S0(n58_adj_5087), .S1(n55_adj_5086));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_996_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_996_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_996_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_996_add_4_3.INJECT1_1 = "NO";
    CCU2C add_3221_5 (.A0(n17128), .B0(amdemod_d_11__N_2308), .C0(GND_net), 
          .D0(VCC_net), .A1(n17129), .B1(amdemod_d_11__N_2305), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15845), .COUT(n15846));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam add_3221_5.INIT0 = 16'h9995;
    defparam add_3221_5.INIT1 = 16'h9995;
    defparam add_3221_5.INJECT1_0 = "NO";
    defparam add_3221_5.INJECT1_1 = "NO";
    LUT4 i1589_3_lut_4_lut (.A(n17288), .B(n17150), .C(led_c_3), .D(n283), 
         .Z(n11311)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1589_3_lut_4_lut.init = 16'hf404;
    LUT4 i1579_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(led_c_3), .D(n301), 
         .Z(n11301)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1579_3_lut_4_lut.init = 16'hf404;
    CCU2C add_3221_3 (.A0(amdemod_d_11__N_1874), .B0(amdemod_d_11__N_2314), 
          .C0(GND_net), .D0(VCC_net), .A1(n17127), .B1(amdemod_d_11__N_2311), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15844), .COUT(n15845));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam add_3221_3.INIT0 = 16'h9995;
    defparam add_3221_3.INIT1 = 16'h9995;
    defparam add_3221_3.INJECT1_0 = "NO";
    defparam add_3221_3.INJECT1_1 = "NO";
    CCU2C _add_1_996_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15313), .S1(n61_adj_5088));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_996_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_996_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_996_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_996_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_37 (.A0(integrator2[70]), .B0(cout_adj_5073), 
          .C0(n81_adj_5312), .D0(integrator3[70]), .A1(integrator2[71]), 
          .B1(cout_adj_5073), .C1(n78_adj_5311), .D1(integrator3[71]), 
          .CIN(n15311), .S0(integrator3_71__N_562[70]), .S1(integrator3_71__N_562[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_35 (.A0(integrator2[68]), .B0(cout_adj_5073), 
          .C0(n87_adj_5314), .D0(integrator3[68]), .A1(integrator2[69]), 
          .B1(cout_adj_5073), .C1(n84_adj_5313), .D1(integrator3[69]), 
          .CIN(n15310), .COUT(n15311), .S0(integrator3_71__N_562[68]), 
          .S1(integrator3_71__N_562[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_35.INJECT1_1 = "NO";
    LUT4 i1663_3_lut_4_lut (.A(n17288), .B(n17150), .C(led_c_3), .D(n154), 
         .Z(n11385)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1663_3_lut_4_lut.init = 16'hf707;
    CCU2C _add_1_1259_add_4_33 (.A0(integrator2[66]), .B0(cout_adj_5073), 
          .C0(n93_adj_5316), .D0(integrator3[66]), .A1(integrator2[67]), 
          .B1(cout_adj_5073), .C1(n90_adj_5315), .D1(integrator3[67]), 
          .CIN(n15309), .COUT(n15310), .S0(integrator3_71__N_562[66]), 
          .S1(integrator3_71__N_562[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_31 (.A0(integrator2[64]), .B0(cout_adj_5073), 
          .C0(n99_adj_5318), .D0(integrator3[64]), .A1(integrator2[65]), 
          .B1(cout_adj_5073), .C1(n96_adj_5317), .D1(integrator3[65]), 
          .CIN(n15308), .COUT(n15309), .S0(integrator3_71__N_562[64]), 
          .S1(integrator3_71__N_562[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_29 (.A0(integrator2[62]), .B0(cout_adj_5073), 
          .C0(n105_adj_5320), .D0(integrator3[62]), .A1(integrator2[63]), 
          .B1(cout_adj_5073), .C1(n102_adj_5319), .D1(integrator3[63]), 
          .CIN(n15307), .COUT(n15308), .S0(integrator3_71__N_562[62]), 
          .S1(integrator3_71__N_562[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_27 (.A0(integrator2[60]), .B0(cout_adj_5073), 
          .C0(n111_adj_5322), .D0(integrator3[60]), .A1(integrator2[61]), 
          .B1(cout_adj_5073), .C1(n108_adj_5321), .D1(integrator3[61]), 
          .CIN(n15306), .COUT(n15307), .S0(integrator3_71__N_562[60]), 
          .S1(integrator3_71__N_562[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_27.INJECT1_1 = "NO";
    LUT4 n16388_bdd_4_lut (.A(n16388), .B(n16238), .C(led_c_2), .D(n17153), 
         .Z(n1827)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n16388_bdd_4_lut.init = 16'hca00;
    CCU2C _add_1_1259_add_4_25 (.A0(integrator2[58]), .B0(cout_adj_5073), 
          .C0(n117_adj_5324), .D0(integrator3[58]), .A1(integrator2[59]), 
          .B1(cout_adj_5073), .C1(n114_adj_5323), .D1(integrator3[59]), 
          .CIN(n15305), .COUT(n15306), .S0(integrator3_71__N_562[58]), 
          .S1(integrator3_71__N_562[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_23 (.A0(integrator2[56]), .B0(cout_adj_5073), 
          .C0(n123_adj_5326), .D0(integrator3[56]), .A1(integrator2[57]), 
          .B1(cout_adj_5073), .C1(n120_adj_5325), .D1(integrator3[57]), 
          .CIN(n15304), .COUT(n15305), .S0(integrator3_71__N_562[56]), 
          .S1(integrator3_71__N_562[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_21 (.A0(integrator2[54]), .B0(cout_adj_5073), 
          .C0(n129_adj_5328), .D0(integrator3[54]), .A1(integrator2[55]), 
          .B1(cout_adj_5073), .C1(n126_adj_5327), .D1(integrator3[55]), 
          .CIN(n15303), .COUT(n15304), .S0(integrator3_71__N_562[54]), 
          .S1(integrator3_71__N_562[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_19 (.A0(integrator2[52]), .B0(cout_adj_5073), 
          .C0(n135_adj_5330), .D0(integrator3[52]), .A1(integrator2[53]), 
          .B1(cout_adj_5073), .C1(n132_adj_5329), .D1(integrator3[53]), 
          .CIN(n15302), .COUT(n15303), .S0(integrator3_71__N_562[52]), 
          .S1(integrator3_71__N_562[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_17 (.A0(integrator2[50]), .B0(cout_adj_5073), 
          .C0(n141_adj_5332), .D0(integrator3[50]), .A1(integrator2[51]), 
          .B1(cout_adj_5073), .C1(n138_adj_5331), .D1(integrator3[51]), 
          .CIN(n15301), .COUT(n15302), .S0(integrator3_71__N_562[50]), 
          .S1(integrator3_71__N_562[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_15 (.A0(integrator2[48]), .B0(cout_adj_5073), 
          .C0(n147_adj_5334), .D0(integrator3[48]), .A1(integrator2[49]), 
          .B1(cout_adj_5073), .C1(n144_adj_5333), .D1(integrator3[49]), 
          .CIN(n15300), .COUT(n15301), .S0(integrator3_71__N_562[48]), 
          .S1(integrator3_71__N_562[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_13 (.A0(integrator2[46]), .B0(cout_adj_5073), 
          .C0(n153_adj_5336), .D0(integrator3[46]), .A1(integrator2[47]), 
          .B1(cout_adj_5073), .C1(n150_adj_5335), .D1(integrator3[47]), 
          .CIN(n15299), .COUT(n15300), .S0(integrator3_71__N_562[46]), 
          .S1(integrator3_71__N_562[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_11 (.A0(integrator2[44]), .B0(cout_adj_5073), 
          .C0(n159_adj_5338), .D0(integrator3[44]), .A1(integrator2[45]), 
          .B1(cout_adj_5073), .C1(n156_adj_5337), .D1(integrator3[45]), 
          .CIN(n15298), .COUT(n15299), .S0(integrator3_71__N_562[44]), 
          .S1(integrator3_71__N_562[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_9 (.A0(integrator2[42]), .B0(cout_adj_5073), 
          .C0(n165_adj_5340), .D0(integrator3[42]), .A1(integrator2[43]), 
          .B1(cout_adj_5073), .C1(n162_adj_5339), .D1(integrator3[43]), 
          .CIN(n15297), .COUT(n15298), .S0(integrator3_71__N_562[42]), 
          .S1(integrator3_71__N_562[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_7 (.A0(integrator2[40]), .B0(cout_adj_5073), 
          .C0(n171_adj_5342), .D0(integrator3[40]), .A1(integrator2[41]), 
          .B1(cout_adj_5073), .C1(n168_adj_5341), .D1(integrator3[41]), 
          .CIN(n15296), .COUT(n15297), .S0(integrator3_71__N_562[40]), 
          .S1(integrator3_71__N_562[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_5 (.A0(integrator2[38]), .B0(cout_adj_5073), 
          .C0(n177_adj_5344), .D0(integrator3[38]), .A1(integrator2[39]), 
          .B1(cout_adj_5073), .C1(n174_adj_5343), .D1(integrator3[39]), 
          .CIN(n15295), .COUT(n15296), .S0(integrator3_71__N_562[38]), 
          .S1(integrator3_71__N_562[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_3 (.A0(integrator2[36]), .B0(cout_adj_5073), 
          .C0(n183_adj_5346), .D0(integrator3[36]), .A1(integrator2[37]), 
          .B1(cout_adj_5073), .C1(n180_adj_5345), .D1(integrator3[37]), 
          .CIN(n15294), .COUT(n15295), .S0(integrator3_71__N_562[36]), 
          .S1(integrator3_71__N_562[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1259_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1259_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1259_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5073), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15294));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1259_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1259_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1259_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1259_add_4_1.INJECT1_1 = "NO";
    LUT4 i4706_2_lut (.A(phase_inc_gen1[0]), .B(phase_accum[0]), .Z(n321)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4706_2_lut.init = 16'h6666;
    CCU2C _add_1_1193_add_4_16 (.A0(amdemod_d_11__N_2137), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15290), .S0(amdemod_d_11__N_1860[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1193_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1193_add_4_16.INIT1 = 16'h0000;
    defparam _add_1_1193_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1193_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1193_add_4_14 (.A0(amdemod_d_11__N_2143), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2140), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15289), .COUT(n15290), .S0(amdemod_d_11__N_1860[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1193_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_1193_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_1193_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1193_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1193_add_4_12 (.A0(amdemod_d_11__N_2149), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2146), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15288), .COUT(n15289), .S0(amdemod_d_11__N_1860[9]), 
          .S1(amdemod_d_11__N_1860[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1193_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_1193_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_1193_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1193_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15386), .S0(cout_adj_5075));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_990_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_990_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_cout.INJECT1_1 = "NO";
    CCU2C add_3221_1 (.A0(square_sum[0]), .B0(GND_net), .C0(GND_net), 
          .D0(square_sum[0]), .A1(amdemod_d_11__N_1874), .B1(square_sum[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15844));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam add_3221_1.INIT0 = 16'h000A;
    defparam add_3221_1.INIT1 = 16'h666a;
    defparam add_3221_1.INJECT1_0 = "NO";
    defparam add_3221_1.INJECT1_1 = "NO";
    CCU2C add_3222_65 (.A0(phase_inc_gen[62]), .B0(n17278), .C0(n11622), 
          .D0(n2545), .A1(phase_inc_gen[63]), .B1(n17278), .C1(n11624), 
          .D1(n2545), .CIN(n15842), .S0(n137), .S1(n134));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_65.INIT0 = 16'h74b8;
    defparam add_3222_65.INIT1 = 16'h74b8;
    defparam add_3222_65.INJECT1_0 = "NO";
    defparam add_3222_65.INJECT1_1 = "NO";
    CCU2C _add_1_987_add_4_10 (.A0(integrator4[8]), .B0(integrator3[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[9]), .B1(integrator3[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15391), .COUT(n15392), .S0(integrator4_71__N_634[8]), 
          .S1(integrator4_71__N_634[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_987_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_987_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_987_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_987_add_4_10.INJECT1_1 = "NO";
    LUT4 i1874_4_lut (.A(n286_adj_5956), .B(n280), .C(led_c_3), .D(n17144), 
         .Z(n11608)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1874_4_lut.init = 16'hcac0;
    LUT4 mux_251_i9_4_lut (.A(n11307), .B(n295_adj_5959), .C(n17136), 
         .D(n2244), .Z(n2036)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i9_4_lut.init = 16'hcfca;
    CCU2C add_3222_63 (.A0(phase_inc_gen[60]), .B0(n17278), .C0(n1984), 
          .D0(n2545), .A1(phase_inc_gen[61]), .B1(n17278), .C1(n11620), 
          .D1(n2545), .CIN(n15841), .COUT(n15842), .S0(n143), .S1(n140));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_63.INIT0 = 16'h74b8;
    defparam add_3222_63.INIT1 = 16'h74b8;
    defparam add_3222_63.INJECT1_0 = "NO";
    defparam add_3222_63.INJECT1_1 = "NO";
    CCU2C add_3222_61 (.A0(phase_inc_gen[58]), .B0(n17278), .C0(n1986), 
          .D0(n2545), .A1(phase_inc_gen[59]), .B1(n17278), .C1(n1985), 
          .D1(n2545), .CIN(n15840), .COUT(n15841), .S0(n149), .S1(n146));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_61.INIT0 = 16'h74b8;
    defparam add_3222_61.INIT1 = 16'h74b8;
    defparam add_3222_61.INJECT1_0 = "NO";
    defparam add_3222_61.INJECT1_1 = "NO";
    FD1S3AX rx_byte_i3_rep_371 (.D(rx_byte1[2]), .CK(clk_80mhz), .Q(n17288));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam rx_byte_i3_rep_371.GSR = "ENABLED";
    CCU2C add_3222_59 (.A0(phase_inc_gen[56]), .B0(n17278), .C0(n1988), 
          .D0(n2545), .A1(phase_inc_gen[57]), .B1(n17278), .C1(n11618), 
          .D1(n2545), .CIN(n15839), .COUT(n15840), .S0(n155), .S1(n152));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_59.INIT0 = 16'h74b8;
    defparam add_3222_59.INIT1 = 16'h74b8;
    defparam add_3222_59.INJECT1_0 = "NO";
    defparam add_3222_59.INJECT1_1 = "NO";
    CCU2C add_3222_57 (.A0(phase_inc_gen[54]), .B0(n17278), .C0(n1990), 
          .D0(n2545), .A1(phase_inc_gen[55]), .B1(n17278), .C1(n1989), 
          .D1(n2545), .CIN(n15838), .COUT(n15839), .S0(n161), .S1(n158));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_57.INIT0 = 16'h74b8;
    defparam add_3222_57.INIT1 = 16'h74b8;
    defparam add_3222_57.INJECT1_0 = "NO";
    defparam add_3222_57.INJECT1_1 = "NO";
    CCU2C add_3222_55 (.A0(phase_inc_gen[52]), .B0(n17278), .C0(n11616), 
          .D0(n2545), .A1(phase_inc_gen[53]), .B1(n17278), .C1(n1991), 
          .D1(n2545), .CIN(n15837), .COUT(n15838), .S0(n167), .S1(n164));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_55.INIT0 = 16'h74b8;
    defparam add_3222_55.INIT1 = 16'h74b8;
    defparam add_3222_55.INJECT1_0 = "NO";
    defparam add_3222_55.INJECT1_1 = "NO";
    CCU2C add_3222_53 (.A0(phase_inc_gen[50]), .B0(n17278), .C0(n1994), 
          .D0(n2559), .A1(phase_inc_gen[51]), .B1(n17278), .C1(n1993), 
          .D1(n2545), .CIN(n15836), .COUT(n15837), .S0(n173), .S1(n170));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_53.INIT0 = 16'h74b8;
    defparam add_3222_53.INIT1 = 16'h74b8;
    defparam add_3222_53.INJECT1_0 = "NO";
    defparam add_3222_53.INJECT1_1 = "NO";
    OB pwm_out_p3_pad (.I(pwm_out_p4_c), .O(pwm_out_p3));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(47[23:33])
    OB pwm_out_p4_pad (.I(pwm_out_p4_c), .O(pwm_out_p4));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(48[23:33])
    OB pwm_out_n1_pad (.I(pwm_out_n4_c), .O(pwm_out_n1));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(49[23:33])
    OB pwm_out_n2_pad (.I(pwm_out_n4_c), .O(pwm_out_n2));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(50[23:33])
    OB pwm_out_n3_pad (.I(pwm_out_n4_c), .O(pwm_out_n3));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(51[23:33])
    OB pwm_out_n4_pad (.I(pwm_out_n4_c), .O(pwm_out_n4));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(52[23:33])
    OB led_pad_7 (.I(led_c_7), .O(led[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(53[23:26])
    OB led_pad_6 (.I(led_c_6), .O(led[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(53[23:26])
    OB led_pad_5 (.I(led_c_5), .O(led[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(53[23:26])
    OB led_pad_4 (.I(led_c_4), .O(led[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(53[23:26])
    OB led_pad_3 (.I(led_c_3), .O(led[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(53[23:26])
    OB led_pad_2 (.I(led_c_2), .O(led[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(53[23:26])
    OB led_pad_1 (.I(led_c_1), .O(led[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(53[23:26])
    OB led_pad_0 (.I(led_c_0), .O(led[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(53[23:26])
    IB clk_25mhz_pad (.I(clk_25mhz), .O(clk_25mhz_c));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(39[16:25])
    IB rx_serial_pad (.I(rx_serial), .O(rx_serial_c));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(40[16:25])
    IB rf_in_pad (.I(rf_in), .O(rf_in_c));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(41[16:21])
    CCU2C add_3222_51 (.A0(phase_inc_gen[48]), .B0(n17278), .C0(n1996), 
          .D0(n2559), .A1(phase_inc_gen[49]), .B1(n17278), .C1(n1995), 
          .D1(n2559), .CIN(n15835), .COUT(n15836), .S0(n179), .S1(n176));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_51.INIT0 = 16'h74b8;
    defparam add_3222_51.INIT1 = 16'h74b8;
    defparam add_3222_51.INJECT1_0 = "NO";
    defparam add_3222_51.INJECT1_1 = "NO";
    FD1S3AX phase_inc_gen1_i1 (.D(phase_inc_gen[1]), .CK(clk_80mhz), .Q(phase_inc_gen1[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i1.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i2 (.D(phase_inc_gen[2]), .CK(clk_80mhz), .Q(phase_inc_gen1[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i2.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i3 (.D(phase_inc_gen[3]), .CK(clk_80mhz), .Q(phase_inc_gen1[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i3.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i4 (.D(phase_inc_gen[4]), .CK(clk_80mhz), .Q(phase_inc_gen1[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i4.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i5 (.D(phase_inc_gen[5]), .CK(clk_80mhz), .Q(phase_inc_gen1[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i5.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i6 (.D(phase_inc_gen[6]), .CK(clk_80mhz), .Q(phase_inc_gen1[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i6.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i7 (.D(phase_inc_gen[7]), .CK(clk_80mhz), .Q(phase_inc_gen1[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i7.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i8 (.D(phase_inc_gen[8]), .CK(clk_80mhz), .Q(phase_inc_gen1[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i8.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i9 (.D(phase_inc_gen[9]), .CK(clk_80mhz), .Q(phase_inc_gen1[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i9.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i10 (.D(phase_inc_gen[10]), .CK(clk_80mhz), .Q(phase_inc_gen1[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i10.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i11 (.D(phase_inc_gen[11]), .CK(clk_80mhz), .Q(phase_inc_gen1[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i11.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i12 (.D(phase_inc_gen[12]), .CK(clk_80mhz), .Q(phase_inc_gen1[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i12.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i13 (.D(phase_inc_gen[13]), .CK(clk_80mhz), .Q(phase_inc_gen1[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i13.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i14 (.D(phase_inc_gen[14]), .CK(clk_80mhz), .Q(phase_inc_gen1[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i14.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i15 (.D(phase_inc_gen[15]), .CK(clk_80mhz), .Q(phase_inc_gen1[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i15.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i16 (.D(phase_inc_gen[16]), .CK(clk_80mhz), .Q(phase_inc_gen1[16]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i16.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i17 (.D(phase_inc_gen[17]), .CK(clk_80mhz), .Q(phase_inc_gen1[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i17.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i18 (.D(phase_inc_gen[18]), .CK(clk_80mhz), .Q(phase_inc_gen1[18]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i18.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i19 (.D(phase_inc_gen[19]), .CK(clk_80mhz), .Q(phase_inc_gen1[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i19.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i20 (.D(phase_inc_gen[20]), .CK(clk_80mhz), .Q(phase_inc_gen1[20]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i20.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i21 (.D(phase_inc_gen[21]), .CK(clk_80mhz), .Q(phase_inc_gen1[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i21.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i22 (.D(phase_inc_gen[22]), .CK(clk_80mhz), .Q(phase_inc_gen1[22]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i22.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i23 (.D(phase_inc_gen[23]), .CK(clk_80mhz), .Q(phase_inc_gen1[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i23.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i24 (.D(phase_inc_gen[24]), .CK(clk_80mhz), .Q(phase_inc_gen1[24]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i24.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i25 (.D(phase_inc_gen[25]), .CK(clk_80mhz), .Q(phase_inc_gen1[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i25.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i26 (.D(phase_inc_gen[26]), .CK(clk_80mhz), .Q(phase_inc_gen1[26]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i26.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i27 (.D(phase_inc_gen[27]), .CK(clk_80mhz), .Q(phase_inc_gen1[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i27.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i28 (.D(phase_inc_gen[28]), .CK(clk_80mhz), .Q(phase_inc_gen1[28]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i28.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i29 (.D(phase_inc_gen[29]), .CK(clk_80mhz), .Q(phase_inc_gen1[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i29.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i30 (.D(phase_inc_gen[30]), .CK(clk_80mhz), .Q(phase_inc_gen1[30]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i30.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i31 (.D(phase_inc_gen[31]), .CK(clk_80mhz), .Q(phase_inc_gen1[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i31.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i32 (.D(phase_inc_gen[32]), .CK(clk_80mhz), .Q(phase_inc_gen1[32]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i32.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i33 (.D(phase_inc_gen[33]), .CK(clk_80mhz), .Q(phase_inc_gen1[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i33.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i34 (.D(phase_inc_gen[34]), .CK(clk_80mhz), .Q(phase_inc_gen1[34]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i34.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i35 (.D(phase_inc_gen[35]), .CK(clk_80mhz), .Q(phase_inc_gen1[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i35.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i36 (.D(phase_inc_gen[36]), .CK(clk_80mhz), .Q(phase_inc_gen1[36]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i36.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i37 (.D(phase_inc_gen[37]), .CK(clk_80mhz), .Q(phase_inc_gen1[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i37.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i38 (.D(phase_inc_gen[38]), .CK(clk_80mhz), .Q(phase_inc_gen1[38]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i38.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i39 (.D(phase_inc_gen[39]), .CK(clk_80mhz), .Q(phase_inc_gen1[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i39.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i40 (.D(phase_inc_gen[40]), .CK(clk_80mhz), .Q(phase_inc_gen1[40]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i40.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i41 (.D(phase_inc_gen[41]), .CK(clk_80mhz), .Q(phase_inc_gen1[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i41.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i42 (.D(phase_inc_gen[42]), .CK(clk_80mhz), .Q(phase_inc_gen1[42]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i42.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i43 (.D(phase_inc_gen[43]), .CK(clk_80mhz), .Q(phase_inc_gen1[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i43.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i44 (.D(phase_inc_gen[44]), .CK(clk_80mhz), .Q(phase_inc_gen1[44]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i44.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i45 (.D(phase_inc_gen[45]), .CK(clk_80mhz), .Q(phase_inc_gen1[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i45.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i46 (.D(phase_inc_gen[46]), .CK(clk_80mhz), .Q(phase_inc_gen1[46]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i46.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i47 (.D(phase_inc_gen[47]), .CK(clk_80mhz), .Q(phase_inc_gen1[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i47.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i48 (.D(phase_inc_gen[48]), .CK(clk_80mhz), .Q(phase_inc_gen1[48]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i48.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i49 (.D(phase_inc_gen[49]), .CK(clk_80mhz), .Q(phase_inc_gen1[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i49.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i50 (.D(phase_inc_gen[50]), .CK(clk_80mhz), .Q(phase_inc_gen1[50]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i50.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i51 (.D(phase_inc_gen[51]), .CK(clk_80mhz), .Q(phase_inc_gen1[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i51.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i52 (.D(phase_inc_gen[52]), .CK(clk_80mhz), .Q(phase_inc_gen1[52]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i52.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i53 (.D(phase_inc_gen[53]), .CK(clk_80mhz), .Q(phase_inc_gen1[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i53.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i54 (.D(phase_inc_gen[54]), .CK(clk_80mhz), .Q(phase_inc_gen1[54]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i54.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i55 (.D(phase_inc_gen[55]), .CK(clk_80mhz), .Q(phase_inc_gen1[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i55.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i56 (.D(phase_inc_gen[56]), .CK(clk_80mhz), .Q(phase_inc_gen1[56]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i56.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i57 (.D(phase_inc_gen[57]), .CK(clk_80mhz), .Q(phase_inc_gen1[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i57.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i58 (.D(phase_inc_gen[58]), .CK(clk_80mhz), .Q(phase_inc_gen1[58]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i58.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i59 (.D(phase_inc_gen[59]), .CK(clk_80mhz), .Q(phase_inc_gen1[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i59.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i60 (.D(phase_inc_gen[60]), .CK(clk_80mhz), .Q(phase_inc_gen1[60]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i60.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i61 (.D(phase_inc_gen[61]), .CK(clk_80mhz), .Q(phase_inc_gen1[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i61.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i62 (.D(phase_inc_gen[62]), .CK(clk_80mhz), .Q(phase_inc_gen1[62]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i62.GSR = "ENABLED";
    FD1S3AX phase_inc_gen1_i63 (.D(phase_inc_gen[63]), .CK(clk_80mhz), .Q(phase_inc_gen1[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen1_i63.GSR = "ENABLED";
    LUT4 i1655_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(n17289), .D(n169), 
         .Z(n11377)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1655_3_lut_4_lut.init = 16'hf808;
    LUT4 i5717_4_lut (.A(led_c_2), .B(n17152), .C(led_c_3), .D(led_c_6), 
         .Z(clk_80mhz_enable_1445)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i5717_4_lut.init = 16'h0004;
    CCU2C add_3222_49 (.A0(phase_inc_gen[46]), .B0(n17278), .C0(n1998), 
          .D0(n11169), .A1(phase_inc_gen[47]), .B1(n17278), .C1(n1997), 
          .D1(n11169), .CIN(n15834), .COUT(n15835), .S0(n185), .S1(n182));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_49.INIT0 = 16'h74b8;
    defparam add_3222_49.INIT1 = 16'h74b8;
    defparam add_3222_49.INJECT1_0 = "NO";
    defparam add_3222_49.INJECT1_1 = "NO";
    CCU2C add_3222_47 (.A0(phase_inc_gen[44]), .B0(n17278), .C0(n2000), 
          .D0(n17148), .A1(phase_inc_gen[45]), .B1(n17278), .C1(n1999), 
          .D1(n2545), .CIN(n15833), .COUT(n15834), .S0(n191), .S1(n188));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_47.INIT0 = 16'h74b8;
    defparam add_3222_47.INIT1 = 16'h74b8;
    defparam add_3222_47.INJECT1_0 = "NO";
    defparam add_3222_47.INJECT1_1 = "NO";
    CCU2C add_3222_45 (.A0(phase_inc_gen[42]), .B0(n17278), .C0(n2002), 
          .D0(n17147), .A1(phase_inc_gen[43]), .B1(n17278), .C1(n2001), 
          .D1(n2579), .CIN(n15832), .COUT(n15833), .S0(n197), .S1(n194));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_45.INIT0 = 16'h74b8;
    defparam add_3222_45.INIT1 = 16'h74b8;
    defparam add_3222_45.INJECT1_0 = "NO";
    defparam add_3222_45.INJECT1_1 = "NO";
    CCU2C _add_1_990_add_4_34 (.A0(integrator5[32]), .B0(integrator4[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5[33]), .B1(integrator4[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15384), .COUT(n15385), .S0(integrator5_71__N_706[32]), 
          .S1(integrator5_71__N_706[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_990_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_990_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_990_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_990_add_4_34.INJECT1_1 = "NO";
    CCU2C add_3222_43 (.A0(phase_inc_gen[40]), .B0(n17278), .C0(n11_adj_5725), 
          .D0(n2559), .A1(phase_inc_gen[41]), .B1(n17278), .C1(n11614), 
          .D1(n2579), .CIN(n15831), .COUT(n15832), .S0(n203), .S1(n200));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_43.INIT0 = 16'h74b8;
    defparam add_3222_43.INIT1 = 16'h74b8;
    defparam add_3222_43.INJECT1_0 = "NO";
    defparam add_3222_43.INJECT1_1 = "NO";
    CCU2C add_3222_41 (.A0(phase_inc_gen[38]), .B0(n17278), .C0(n2006), 
          .D0(n2545), .A1(phase_inc_gen[39]), .B1(n17278), .C1(n2005), 
          .D1(n2545), .CIN(n15830), .COUT(n15831), .S0(n209), .S1(n206));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_41.INIT0 = 16'h74b8;
    defparam add_3222_41.INIT1 = 16'h74b8;
    defparam add_3222_41.INJECT1_0 = "NO";
    defparam add_3222_41.INJECT1_1 = "NO";
    CCU2C add_3222_39 (.A0(phase_inc_gen[36]), .B0(n17278), .C0(n2008), 
          .D0(n17148), .A1(phase_inc_gen[37]), .B1(n17278), .C1(n2007), 
          .D1(n2580), .CIN(n15829), .COUT(n15830), .S0(n215), .S1(n212));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_39.INIT0 = 16'h74b8;
    defparam add_3222_39.INIT1 = 16'h74b8;
    defparam add_3222_39.INJECT1_0 = "NO";
    defparam add_3222_39.INJECT1_1 = "NO";
    CCU2C _add_1_1193_add_4_10 (.A0(n17137), .B0(amdemod_d_11__N_2155), 
          .C0(GND_net), .D0(VCC_net), .A1(square_sum[23]), .B1(square_sum[22]), 
          .C1(amdemod_d_11__N_2152), .D1(VCC_net), .CIN(n15287), .COUT(n15288), 
          .S0(amdemod_d_11__N_1860[7]), .S1(amdemod_d_11__N_1860[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1193_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1193_add_4_10.INIT1 = 16'he1e1;
    defparam _add_1_1193_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1193_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_34 (.A0(comb_d9[67]), .B0(comb9[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[68]), .B1(comb9[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15643), .COUT(n15644), .S0(n90_adj_5893), 
          .S1(n87_adj_5892));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_32 (.A0(comb_d9[65]), .B0(comb9[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[66]), .B1(comb9[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15642), .COUT(n15643), .S0(n96_adj_5895), 
          .S1(n93_adj_5894));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_30 (.A0(comb_d9[63]), .B0(comb9[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[64]), .B1(comb9[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15641), .COUT(n15642), .S0(n102_adj_5897), 
          .S1(n99_adj_5896));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_28 (.A0(comb_d9[61]), .B0(comb9[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[62]), .B1(comb9[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15640), .COUT(n15641), .S0(n108_adj_5899), 
          .S1(n105_adj_5898));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_26 (.A0(comb_d9[59]), .B0(comb9[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[60]), .B1(comb9[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15639), .COUT(n15640), .S0(n114_adj_5901), 
          .S1(n111_adj_5900));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_24 (.A0(comb_d9[57]), .B0(comb9[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[58]), .B1(comb9[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15638), .COUT(n15639), .S0(n120_adj_5903), 
          .S1(n117_adj_5902));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_22 (.A0(comb_d9[55]), .B0(comb9[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[56]), .B1(comb9[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15637), .COUT(n15638));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_20 (.A0(comb_d9[53]), .B0(comb9[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[54]), .B1(comb9[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15636), .COUT(n15637));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_18 (.A0(comb_d9[51]), .B0(comb9[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[52]), .B1(comb9[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15635), .COUT(n15636));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_16 (.A0(comb_d9[49]), .B0(comb9[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[50]), .B1(comb9[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15634), .COUT(n15635));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_16.INJECT1_1 = "NO";
    CCU2C add_3222_37 (.A0(phase_inc_gen[34]), .B0(n17278), .C0(n2010), 
          .D0(n17148), .A1(phase_inc_gen[35]), .B1(n17278), .C1(n2009), 
          .D1(n2545), .CIN(n15828), .COUT(n15829), .S0(n221), .S1(n218));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_37.INIT0 = 16'h74b8;
    defparam add_3222_37.INIT1 = 16'h74b8;
    defparam add_3222_37.INJECT1_0 = "NO";
    defparam add_3222_37.INJECT1_1 = "NO";
    CCU2C add_3222_35 (.A0(phase_inc_gen[32]), .B0(n17278), .C0(n2012), 
          .D0(n2559), .A1(phase_inc_gen[33]), .B1(n17278), .C1(n2011), 
          .D1(n2580), .CIN(n15827), .COUT(n15828), .S0(n227), .S1(n224));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_35.INIT0 = 16'h74b8;
    defparam add_3222_35.INIT1 = 16'h74b8;
    defparam add_3222_35.INJECT1_0 = "NO";
    defparam add_3222_35.INJECT1_1 = "NO";
    CCU2C add_3222_33 (.A0(phase_inc_gen[30]), .B0(n17278), .C0(n2014), 
          .D0(n2559), .A1(phase_inc_gen[31]), .B1(n17278), .C1(n2013), 
          .D1(n2594), .CIN(n15826), .COUT(n15827), .S0(n233), .S1(n230));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_33.INIT0 = 16'h74b8;
    defparam add_3222_33.INIT1 = 16'h74b8;
    defparam add_3222_33.INJECT1_0 = "NO";
    defparam add_3222_33.INJECT1_1 = "NO";
    CCU2C add_3222_31 (.A0(phase_inc_gen[28]), .B0(n17278), .C0(n2016), 
          .D0(n2579), .A1(phase_inc_gen[29]), .B1(n17278), .C1(n2015), 
          .D1(n17147), .CIN(n15825), .COUT(n15826), .S0(n239), .S1(n236));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_31.INIT0 = 16'h74b8;
    defparam add_3222_31.INIT1 = 16'h74b8;
    defparam add_3222_31.INJECT1_0 = "NO";
    defparam add_3222_31.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_14 (.A0(comb_d9[47]), .B0(comb9[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[48]), .B1(comb9[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15633), .COUT(n15634));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_12 (.A0(comb_d9[45]), .B0(comb9[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[46]), .B1(comb9[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15632), .COUT(n15633));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_10 (.A0(comb_d9[43]), .B0(comb9[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[44]), .B1(comb9[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15631), .COUT(n15632));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_8 (.A0(comb_d9[41]), .B0(comb9[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[42]), .B1(comb9[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15630), .COUT(n15631));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_6 (.A0(comb_d9[39]), .B0(comb9[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[40]), .B1(comb9[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15629), .COUT(n15630));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_4 (.A0(comb_d9[37]), .B0(comb9[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[38]), .B1(comb9[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15628), .COUT(n15629));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1154_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1154_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[36]), .B1(comb9[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15628));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1154_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1154_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1154_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1154_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1223_add_4_16 (.A0(amdemod_d_11__N_1860[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15627), .S0(n34_adj_5876));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1223_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1223_add_4_16.INIT1 = 16'h0000;
    defparam _add_1_1223_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1223_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1223_add_4_14 (.A0(amdemod_d_11__N_1860[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1860[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15626), .COUT(n15627), .S0(n40_adj_5877));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1223_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_1223_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_1223_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1223_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1223_add_4_12 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1860[7]), .D0(VCC_net), .A1(amdemod_d_11__N_1860[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n15625), .COUT(n15626), 
          .S0(n46_adj_5879), .S1(n43_adj_5878));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1223_add_4_12.INIT0 = 16'he1e1;
    defparam _add_1_1223_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_1223_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1223_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_23 (.A0(comb8_adj_6029[56]), .B0(cout_adj_5310), 
          .C0(n123_adj_5639), .D0(n17_adj_4961), .A1(comb8_adj_6029[57]), 
          .B1(cout_adj_5310), .C1(n120_adj_5638), .D1(n16_adj_4960), .CIN(n14972), 
          .COUT(n14973), .S0(comb9_71__N_1667_adj_6055[56]), .S1(comb9_71__N_1667_adj_6055[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_21 (.A0(comb8_adj_6029[54]), .B0(cout_adj_5310), 
          .C0(n129_adj_5641), .D0(n19_adj_4963), .A1(comb8_adj_6029[55]), 
          .B1(cout_adj_5310), .C1(n126_adj_5640), .D1(n18_adj_4962), .CIN(n14971), 
          .COUT(n14972), .S0(comb9_71__N_1667_adj_6055[54]), .S1(comb9_71__N_1667_adj_6055[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_19 (.A0(comb8_adj_6029[52]), .B0(cout_adj_5310), 
          .C0(n135_adj_5643), .D0(n21_adj_4965), .A1(comb8_adj_6029[53]), 
          .B1(cout_adj_5310), .C1(n132_adj_5642), .D1(n20_adj_4964), .CIN(n14970), 
          .COUT(n14971), .S0(comb9_71__N_1667_adj_6055[52]), .S1(comb9_71__N_1667_adj_6055[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_17 (.A0(comb8_adj_6029[50]), .B0(cout_adj_5310), 
          .C0(n141_adj_5645), .D0(n23_adj_4967), .A1(comb8_adj_6029[51]), 
          .B1(cout_adj_5310), .C1(n138_adj_5644), .D1(n22_adj_4966), .CIN(n14969), 
          .COUT(n14970), .S0(comb9_71__N_1667_adj_6055[50]), .S1(comb9_71__N_1667_adj_6055[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_15 (.A0(comb8_adj_6029[48]), .B0(cout_adj_5310), 
          .C0(n147_adj_5647), .D0(n25_adj_4969), .A1(comb8_adj_6029[49]), 
          .B1(cout_adj_5310), .C1(n144_adj_5646), .D1(n24_adj_4968), .CIN(n14968), 
          .COUT(n14969), .S0(comb9_71__N_1667_adj_6055[48]), .S1(comb9_71__N_1667_adj_6055[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_13 (.A0(comb8_adj_6029[46]), .B0(cout_adj_5310), 
          .C0(n153_adj_5649), .D0(n27_adj_4971), .A1(comb8_adj_6029[47]), 
          .B1(cout_adj_5310), .C1(n150_adj_5648), .D1(n26_adj_4970), .CIN(n14967), 
          .COUT(n14968), .S0(comb9_71__N_1667_adj_6055[46]), .S1(comb9_71__N_1667_adj_6055[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_11 (.A0(comb8_adj_6029[44]), .B0(cout_adj_5310), 
          .C0(n159_adj_5651), .D0(n29_adj_4973), .A1(comb8_adj_6029[45]), 
          .B1(cout_adj_5310), .C1(n156_adj_5650), .D1(n28_adj_4972), .CIN(n14966), 
          .COUT(n14967), .S0(comb9_71__N_1667_adj_6055[44]), .S1(comb9_71__N_1667_adj_6055[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_9 (.A0(comb8_adj_6029[42]), .B0(cout_adj_5310), 
          .C0(n165_adj_5653), .D0(n31_adj_4975), .A1(comb8_adj_6029[43]), 
          .B1(cout_adj_5310), .C1(n162_adj_5652), .D1(n30_adj_4974), .CIN(n14965), 
          .COUT(n14966), .S0(comb9_71__N_1667_adj_6055[42]), .S1(comb9_71__N_1667_adj_6055[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_7 (.A0(comb8_adj_6029[40]), .B0(cout_adj_5310), 
          .C0(n171_adj_5655), .D0(n33_adj_4977), .A1(comb8_adj_6029[41]), 
          .B1(cout_adj_5310), .C1(n168_adj_5654), .D1(n32_adj_4976), .CIN(n14964), 
          .COUT(n14965), .S0(comb9_71__N_1667_adj_6055[40]), .S1(comb9_71__N_1667_adj_6055[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_5 (.A0(comb8_adj_6029[38]), .B0(cout_adj_5310), 
          .C0(n177_adj_5657), .D0(n35_adj_4979), .A1(comb8_adj_6029[39]), 
          .B1(cout_adj_5310), .C1(n174_adj_5656), .D1(n34_adj_4978), .CIN(n14963), 
          .COUT(n14964), .S0(comb9_71__N_1667_adj_6055[38]), .S1(comb9_71__N_1667_adj_6055[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_3 (.A0(comb8_adj_6029[36]), .B0(cout_adj_5310), 
          .C0(n183_adj_5659), .D0(n37_adj_4981), .A1(comb8_adj_6029[37]), 
          .B1(cout_adj_5310), .C1(n180_adj_5658), .D1(n36_adj_4980), .CIN(n14962), 
          .COUT(n14963), .S0(comb9_71__N_1667_adj_6055[36]), .S1(comb9_71__N_1667_adj_6055[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1088_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1088_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1088_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5310), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14962));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1088_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1088_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1088_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1088_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1061_add_4_15 (.A0(amdemod_d_11__N_1861[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14958), .S0(n32_adj_5611));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1061_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1061_add_4_15.INIT1 = 16'h0000;
    defparam _add_1_1061_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1061_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1061_add_4_13 (.A0(amdemod_d_11__N_1861[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1861[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14957), .COUT(n14958), .S0(n38_adj_5612));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1061_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1061_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1061_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1061_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1061_add_4_11 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1861[7]), .D0(VCC_net), .A1(amdemod_d_11__N_1861[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n14956), .COUT(n14957), 
          .S0(n44_adj_5614), .S1(n41_adj_5613));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1061_add_4_11.INIT0 = 16'h1e1e;
    defparam _add_1_1061_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1061_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1061_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1061_add_4_9 (.A0(n17134), .B0(amdemod_d_11__N_1861[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1861[6]), .B1(n17162), 
          .C1(n17279), .D1(n17146), .CIN(n14955), .COUT(n14956), .S0(n50_adj_5616), 
          .S1(n47_adj_5615));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1061_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1061_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_1061_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1061_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1061_add_4_7 (.A0(n17132), .B0(amdemod_d_11__N_1861[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17133), .B1(amdemod_d_11__N_1861[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14954), .COUT(n14955), .S0(n56_adj_5618), 
          .S1(n53_adj_5617));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1061_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1061_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1061_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1061_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1061_add_4_5 (.A0(n17130), .B0(amdemod_d_11__N_1861[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17131), .B1(amdemod_d_11__N_1861[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14953), .COUT(n14954), .S0(n62_adj_5620), 
          .S1(n59_adj_5619));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1061_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1061_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1061_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1061_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1061_add_4_3 (.A0(square_sum[7]), .B0(amdemod_d_11__N_1861[13]), 
          .C0(n17130), .D0(amdemod_d_11__N_1860[13]), .A1(n17129), .B1(amdemod_d_11__N_1861[0]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14952), .COUT(n14953), .S0(n68_adj_5622), 
          .S1(n65_adj_5621));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1061_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_1061_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1061_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1061_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1061_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14952), .S1(n71_adj_5623));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1061_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1061_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1061_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1061_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14951), .S0(cout_adj_5164));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1002_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1002_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_36 (.A0(integrator3_adj_6022[34]), .B0(integrator2_adj_6021[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[35]), .B1(integrator2_adj_6021[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14950), .COUT(n14951), .S0(integrator3_71__N_562_adj_6038[34]), 
          .S1(integrator3_71__N_562_adj_6038[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_34 (.A0(integrator3_adj_6022[32]), .B0(integrator2_adj_6021[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[33]), .B1(integrator2_adj_6021[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14949), .COUT(n14950), .S0(integrator3_71__N_562_adj_6038[32]), 
          .S1(integrator3_71__N_562_adj_6038[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_32 (.A0(integrator3_adj_6022[30]), .B0(integrator2_adj_6021[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[31]), .B1(integrator2_adj_6021[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14948), .COUT(n14949), .S0(integrator3_71__N_562_adj_6038[30]), 
          .S1(integrator3_71__N_562_adj_6038[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_30 (.A0(integrator3_adj_6022[28]), .B0(integrator2_adj_6021[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[29]), .B1(integrator2_adj_6021[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14947), .COUT(n14948), .S0(integrator3_71__N_562_adj_6038[28]), 
          .S1(integrator3_71__N_562_adj_6038[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_28 (.A0(integrator3_adj_6022[26]), .B0(integrator2_adj_6021[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[27]), .B1(integrator2_adj_6021[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14946), .COUT(n14947), .S0(integrator3_71__N_562_adj_6038[26]), 
          .S1(integrator3_71__N_562_adj_6038[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_26 (.A0(integrator3_adj_6022[24]), .B0(integrator2_adj_6021[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[25]), .B1(integrator2_adj_6021[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14945), .COUT(n14946), .S0(integrator3_71__N_562_adj_6038[24]), 
          .S1(integrator3_71__N_562_adj_6038[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_24 (.A0(integrator3_adj_6022[22]), .B0(integrator2_adj_6021[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[23]), .B1(integrator2_adj_6021[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14944), .COUT(n14945), .S0(integrator3_71__N_562_adj_6038[22]), 
          .S1(integrator3_71__N_562_adj_6038[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_22 (.A0(integrator3_adj_6022[20]), .B0(integrator2_adj_6021[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[21]), .B1(integrator2_adj_6021[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14943), .COUT(n14944), .S0(integrator3_71__N_562_adj_6038[20]), 
          .S1(integrator3_71__N_562_adj_6038[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_20 (.A0(integrator3_adj_6022[18]), .B0(integrator2_adj_6021[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[19]), .B1(integrator2_adj_6021[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14942), .COUT(n14943), .S0(integrator3_71__N_562_adj_6038[18]), 
          .S1(integrator3_71__N_562_adj_6038[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_18 (.A0(integrator3_adj_6022[16]), .B0(integrator2_adj_6021[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[17]), .B1(integrator2_adj_6021[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14941), .COUT(n14942), .S0(integrator3_71__N_562_adj_6038[16]), 
          .S1(integrator3_71__N_562_adj_6038[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_16 (.A0(integrator3_adj_6022[14]), .B0(integrator2_adj_6021[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[15]), .B1(integrator2_adj_6021[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14940), .COUT(n14941), .S0(integrator3_71__N_562_adj_6038[14]), 
          .S1(integrator3_71__N_562_adj_6038[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_14 (.A0(integrator3_adj_6022[12]), .B0(integrator2_adj_6021[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[13]), .B1(integrator2_adj_6021[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14939), .COUT(n14940), .S0(integrator3_71__N_562_adj_6038[12]), 
          .S1(integrator3_71__N_562_adj_6038[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_12 (.A0(integrator3_adj_6022[10]), .B0(integrator2_adj_6021[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[11]), .B1(integrator2_adj_6021[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14938), .COUT(n14939), .S0(integrator3_71__N_562_adj_6038[10]), 
          .S1(integrator3_71__N_562_adj_6038[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_12.INJECT1_1 = "NO";
    FD1S3AX square_sum_e3__i2 (.D(n118_adj_5724), .CK(cic_sine_clk), .Q(square_sum[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i2.GSR = "ENABLED";
    CCU2C add_3222_29 (.A0(phase_inc_gen[26]), .B0(n17278), .C0(n2018), 
          .D0(n2545), .A1(phase_inc_gen[27]), .B1(n17278), .C1(n2017), 
          .D1(n2580), .CIN(n15824), .COUT(n15825), .S0(n245), .S1(n242));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_29.INIT0 = 16'h74b8;
    defparam add_3222_29.INIT1 = 16'h74b8;
    defparam add_3222_29.INJECT1_0 = "NO";
    defparam add_3222_29.INJECT1_1 = "NO";
    CCU2C add_3222_27 (.A0(phase_inc_gen[24]), .B0(n17278), .C0(n2020), 
          .D0(n2545), .A1(phase_inc_gen[25]), .B1(n17278), .C1(n2019), 
          .D1(n2545), .CIN(n15823), .COUT(n15824), .S0(n251), .S1(n248));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_27.INIT0 = 16'h74b8;
    defparam add_3222_27.INIT1 = 16'h74b8;
    defparam add_3222_27.INJECT1_0 = "NO";
    defparam add_3222_27.INJECT1_1 = "NO";
    CCU2C add_3222_25 (.A0(phase_inc_gen[22]), .B0(n17278), .C0(n11_adj_4729), 
          .D0(n17148), .A1(phase_inc_gen[23]), .B1(n17278), .C1(n2021), 
          .D1(n17147), .CIN(n15822), .COUT(n15823), .S0(n257), .S1(n254));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_25.INIT0 = 16'h74b8;
    defparam add_3222_25.INIT1 = 16'h74b8;
    defparam add_3222_25.INJECT1_0 = "NO";
    defparam add_3222_25.INJECT1_1 = "NO";
    CCU2C add_3222_23 (.A0(phase_inc_gen[20]), .B0(n17278), .C0(n2024), 
          .D0(n2545), .A1(phase_inc_gen[21]), .B1(n17278), .C1(n11612), 
          .D1(n2559), .CIN(n15821), .COUT(n15822), .S0(n263), .S1(n260));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_23.INIT0 = 16'h74b8;
    defparam add_3222_23.INIT1 = 16'h74b8;
    defparam add_3222_23.INJECT1_0 = "NO";
    defparam add_3222_23.INJECT1_1 = "NO";
    CCU2C add_3222_21 (.A0(phase_inc_gen[18]), .B0(n17278), .C0(n2026), 
          .D0(n17147), .A1(phase_inc_gen[19]), .B1(n17278), .C1(n11610), 
          .D1(n2580), .CIN(n15820), .COUT(n15821), .S0(n269), .S1(n266));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_21.INIT0 = 16'h74b8;
    defparam add_3222_21.INIT1 = 16'h74b8;
    defparam add_3222_21.INJECT1_0 = "NO";
    defparam add_3222_21.INJECT1_1 = "NO";
    CCU2C add_3222_19 (.A0(phase_inc_gen[16]), .B0(n17278), .C0(n2028), 
          .D0(n2594), .A1(phase_inc_gen[17]), .B1(n17278), .C1(n2027), 
          .D1(n11169), .CIN(n15819), .COUT(n15820), .S0(n275), .S1(n272));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_19.INIT0 = 16'h74b8;
    defparam add_3222_19.INIT1 = 16'h74b8;
    defparam add_3222_19.INJECT1_0 = "NO";
    defparam add_3222_19.INJECT1_1 = "NO";
    CCU2C add_3222_17 (.A0(phase_inc_gen[14]), .B0(n17278), .C0(n2030), 
          .D0(n17148), .A1(phase_inc_gen[15]), .B1(n17278), .C1(n2029), 
          .D1(n2580), .CIN(n15818), .COUT(n15819), .S0(n281), .S1(n278));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_17.INIT0 = 16'h74b8;
    defparam add_3222_17.INIT1 = 16'h74b8;
    defparam add_3222_17.INJECT1_0 = "NO";
    defparam add_3222_17.INJECT1_1 = "NO";
    CCU2C add_3222_15 (.A0(phase_inc_gen[12]), .B0(n17278), .C0(n2032), 
          .D0(n17148), .A1(phase_inc_gen[13]), .B1(n17278), .C1(n2031), 
          .D1(n2594), .CIN(n15817), .COUT(n15818), .S0(n287), .S1(n284));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_15.INIT0 = 16'h74b8;
    defparam add_3222_15.INIT1 = 16'h74b8;
    defparam add_3222_15.INJECT1_0 = "NO";
    defparam add_3222_15.INJECT1_1 = "NO";
    CCU2C add_3222_13 (.A0(phase_inc_gen[10]), .B0(n17278), .C0(n2034), 
          .D0(n2594), .A1(phase_inc_gen[11]), .B1(n17278), .C1(n11608), 
          .D1(n2545), .CIN(n15816), .COUT(n15817), .S0(n293), .S1(n290));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_13.INIT0 = 16'h74b8;
    defparam add_3222_13.INIT1 = 16'h74b8;
    defparam add_3222_13.INJECT1_0 = "NO";
    defparam add_3222_13.INJECT1_1 = "NO";
    CCU2C add_3222_11 (.A0(phase_inc_gen[8]), .B0(n17278), .C0(n2036), 
          .D0(n2579), .A1(phase_inc_gen[9]), .B1(n17278), .C1(n2035), 
          .D1(n17147), .CIN(n15815), .COUT(n15816), .S0(n299), .S1(n296));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_11.INIT0 = 16'h74b8;
    defparam add_3222_11.INIT1 = 16'h74b8;
    defparam add_3222_11.INJECT1_0 = "NO";
    defparam add_3222_11.INJECT1_1 = "NO";
    CCU2C _add_1_1193_add_4_8 (.A0(amdemod_d_11__N_2161), .B0(amdemod_d_11__N_1841[11]), 
          .C0(n17134), .D0(amdemod_d_11__N_1840[11]), .A1(n17134), .B1(amdemod_d_11__N_2158), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15286), .COUT(n15287), .S0(amdemod_d_11__N_1860[5]), 
          .S1(amdemod_d_11__N_1860[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1193_add_4_8.INIT0 = 16'h656a;
    defparam _add_1_1193_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1193_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1193_add_4_8.INJECT1_1 = "NO";
    FD1S3AX square_sum_e3__i3 (.D(n115_adj_5723), .CK(cic_sine_clk), .Q(square_sum[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i3.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i4 (.D(n112_adj_5722), .CK(cic_sine_clk), .Q(square_sum[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i4.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i5 (.D(n109_adj_5721), .CK(cic_sine_clk), .Q(square_sum[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i5.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i6 (.D(n106_adj_5720), .CK(cic_sine_clk), .Q(square_sum[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i6.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i7 (.D(n103_adj_5719), .CK(cic_sine_clk), .Q(square_sum[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i7.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i8 (.D(n100_adj_5718), .CK(cic_sine_clk), .Q(square_sum[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i8.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i9 (.D(n97_adj_5717), .CK(cic_sine_clk), .Q(square_sum[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i9.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i10 (.D(n94_adj_5716), .CK(cic_sine_clk), .Q(square_sum[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i10.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i11 (.D(n91_adj_5715), .CK(cic_sine_clk), .Q(square_sum[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i11.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i12 (.D(n88_adj_5714), .CK(cic_sine_clk), .Q(square_sum[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i12.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i13 (.D(n85_adj_5713), .CK(cic_sine_clk), .Q(square_sum[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i13.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i14 (.D(n82_adj_5712), .CK(cic_sine_clk), .Q(square_sum[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i14.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i15 (.D(n79_adj_5711), .CK(cic_sine_clk), .Q(square_sum[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i15.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i16 (.D(n76_adj_5710), .CK(cic_sine_clk), .Q(square_sum[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i16.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i17 (.D(n73_adj_5709), .CK(cic_sine_clk), .Q(square_sum[16]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i17.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i18 (.D(n70_adj_5708), .CK(cic_sine_clk), .Q(square_sum[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i18.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i19 (.D(n67_adj_5707), .CK(cic_sine_clk), .Q(square_sum[18]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i19.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i20 (.D(n64_adj_5706), .CK(cic_sine_clk), .Q(square_sum[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i20.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i21 (.D(n61_adj_5705), .CK(cic_sine_clk), .Q(square_sum[20]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i21.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i22 (.D(n58_adj_5704), .CK(cic_sine_clk), .Q(square_sum[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i22.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i23 (.D(n55_adj_5703), .CK(cic_sine_clk), .Q(square_sum[22]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i23.GSR = "ENABLED";
    FD1S3AX square_sum_e3__i24 (.D(n52_adj_5702), .CK(cic_sine_clk), .Q(square_sum[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e3__i24.GSR = "ENABLED";
    CCU2C _add_1_1223_add_4_10 (.A0(n17134), .B0(amdemod_d_11__N_1860[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17137), .B1(amdemod_d_11__N_1860[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15624), .COUT(n15625), .S0(n52_adj_5881), 
          .S1(n49_adj_5880));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1223_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1223_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1223_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1223_add_4_10.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_26 (.A0(phase_inc_gen1[24]), .B0(phase_accum[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[25]), .B1(phase_accum[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15481), .COUT(n15482), .S0(n249), 
          .S1(n246));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_26.INIT0 = 16'h666a;
    defparam phase_accum_add_4_26.INIT1 = 16'h666a;
    defparam phase_accum_add_4_26.INJECT1_0 = "NO";
    defparam phase_accum_add_4_26.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_353_4_lut_4_lut (.A(led_c_0), .B(n17158), .C(n17155), 
         .D(led_c_6), .Z(n17150)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_3_lut_rep_353_4_lut_4_lut.init = 16'h4000;
    CCU2C _add_1_1193_add_4_6 (.A0(amdemod_d_11__N_2167), .B0(amdemod_d_11__N_1851[13]), 
          .C0(n17132), .D0(amdemod_d_11__N_1850[13]), .A1(n17132), .B1(amdemod_d_11__N_2164), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15285), .COUT(n15286), .S0(amdemod_d_11__N_1860[3]), 
          .S1(amdemod_d_11__N_1860[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1193_add_4_6.INIT0 = 16'h656a;
    defparam _add_1_1193_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1193_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1193_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1223_add_4_8 (.A0(n17132), .B0(amdemod_d_11__N_1860[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1860[4]), .B1(amdemod_d_11__N_1841[11]), 
          .C1(n17134), .D1(amdemod_d_11__N_1840[11]), .CIN(n15623), .COUT(n15624), 
          .S0(n58_adj_5883), .S1(n55_adj_5882));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1223_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1223_add_4_8.INIT1 = 16'h656a;
    defparam _add_1_1223_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1223_add_4_8.INJECT1_1 = "NO";
    CCU2C add_3222_9 (.A0(phase_inc_gen[6]), .B0(n17278), .C0(n2038), 
          .D0(n2580), .A1(phase_inc_gen[7]), .B1(n17278), .C1(n2037), 
          .D1(n17147), .CIN(n15814), .COUT(n15815), .S0(n305), .S1(n302));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_9.INIT0 = 16'h74b8;
    defparam add_3222_9.INIT1 = 16'h74b8;
    defparam add_3222_9.INJECT1_0 = "NO";
    defparam add_3222_9.INJECT1_1 = "NO";
    CCU2C add_3222_7 (.A0(phase_inc_gen[4]), .B0(n17278), .C0(n2040), 
          .D0(n2580), .A1(phase_inc_gen[5]), .B1(n17278), .C1(n2039), 
          .D1(n2580), .CIN(n15813), .COUT(n15814), .S0(n311), .S1(n308));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_7.INIT0 = 16'h74b8;
    defparam add_3222_7.INIT1 = 16'h74b8;
    defparam add_3222_7.INJECT1_0 = "NO";
    defparam add_3222_7.INJECT1_1 = "NO";
    CCU2C add_3222_5 (.A0(phase_inc_gen[2]), .B0(n17278), .C0(n17175), 
          .D0(n11169), .A1(phase_inc_gen[3]), .B1(n17278), .C1(n17178), 
          .D1(n11169), .CIN(n15812), .COUT(n15813), .S0(n317), .S1(n314));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_5.INIT0 = 16'h74b8;
    defparam add_3222_5.INIT1 = 16'h74b8;
    defparam add_3222_5.INJECT1_0 = "NO";
    defparam add_3222_5.INJECT1_1 = "NO";
    CCU2C add_3222_3 (.A0(phase_inc_gen[0]), .B0(n17278), .C0(n15867), 
          .D0(n17147), .A1(phase_inc_gen[1]), .B1(n17278), .C1(n17174), 
          .D1(n2594), .CIN(n15811), .COUT(n15812), .S0(n323), .S1(n320));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_3.INIT0 = 16'h74b8;
    defparam add_3222_3.INIT1 = 16'h74b8;
    defparam add_3222_3.INJECT1_0 = "NO";
    defparam add_3222_3.INJECT1_1 = "NO";
    CCU2C add_3222_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n16348), .B1(n12278), .C1(led_c_4), .D1(n1827), .COUT(n15811));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam add_3222_1.INIT0 = 16'h0000;
    defparam add_3222_1.INIT1 = 16'hf7ff;
    defparam add_3222_1.INJECT1_0 = "NO";
    defparam add_3222_1.INJECT1_1 = "NO";
    CCU2C _add_1_1223_add_4_6 (.A0(n17130), .B0(amdemod_d_11__N_1860[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1860[2]), .B1(amdemod_d_11__N_1851[13]), 
          .C1(n17132), .D1(amdemod_d_11__N_1850[13]), .CIN(n15622), .COUT(n15623), 
          .S0(n64_adj_5885), .S1(n61_adj_5884));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1223_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1223_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_1223_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1223_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1226_add_4_16 (.A0(amdemod_d_11__N_1851[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15807), .S0(n34_adj_6002));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1226_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1226_add_4_16.INIT1 = 16'h0000;
    defparam _add_1_1226_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1226_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1226_add_4_14 (.A0(amdemod_d_11__N_1851[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1851[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15806), .COUT(n15807), .S0(n40_adj_6003));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1226_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_1226_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_1226_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1226_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1226_add_4_12 (.A0(amdemod_d_11__N_1851[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1851[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15805), .COUT(n15806), .S0(n46_adj_6005), 
          .S1(n43_adj_6004));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1226_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_1226_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_1226_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1226_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1223_add_4_4 (.A0(n17129), .B0(square_sum[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_d_11__N_1860[0]), .B1(amdemod_d_11__N_1861[13]), 
          .C1(n17130), .D1(amdemod_d_11__N_1860[13]), .CIN(n15621), .COUT(n15622), 
          .S0(n70_adj_5887), .S1(n67_adj_5886));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1223_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1223_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_1223_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1223_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1226_add_4_10 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1851[5]), .D0(VCC_net), .A1(amdemod_d_11__N_1851[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n15804), .COUT(n15805), 
          .S0(n52_adj_6007), .S1(n49_adj_6006));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1226_add_4_10.INIT0 = 16'he1e1;
    defparam _add_1_1226_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_1226_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1226_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1226_add_4_8 (.A0(n17134), .B0(amdemod_d_11__N_1851[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17137), .B1(amdemod_d_11__N_1851[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15803), .COUT(n15804), .S0(n58_adj_6009), 
          .S1(n55_adj_6008));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1226_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1226_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1226_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1226_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1223_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15621), .S1(n73_adj_5888));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1223_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1223_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1223_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1223_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1226_add_4_6 (.A0(n17132), .B0(amdemod_d_11__N_1851[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1851[2]), .B1(amdemod_d_11__N_1841[11]), 
          .C1(n17134), .D1(amdemod_d_11__N_1840[11]), .CIN(n15802), .COUT(n15803), 
          .S0(n64_adj_6011), .S1(n61_adj_6010));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1226_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1226_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_1226_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1226_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1226_add_4_4 (.A0(n17131), .B0(square_sum[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_d_11__N_1851[0]), .B1(amdemod_d_11__N_1851[13]), 
          .C1(n17132), .D1(amdemod_d_11__N_1850[13]), .CIN(n15801), .COUT(n15802), 
          .S0(n70_adj_6013), .S1(n67_adj_6012));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1226_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1226_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_1226_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1226_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1226_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15801), .S1(n73_adj_6014));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1226_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1226_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1226_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1226_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1238_add_4_13 (.A0(n17134), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15800), .S0(amdemod_d_11__N_1841[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1238_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1238_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_1238_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1238_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1238_add_4_11 (.A0(amdemod_d_11__N_2005), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(n17134), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15799), .COUT(n15800), .S0(amdemod_d_11__N_1841[9]), 
          .S1(amdemod_d_11__N_1841[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1238_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1238_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1238_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1238_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1238_add_4_9 (.A0(amdemod_d_11__N_2011), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2008), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15798), .COUT(n15799), .S0(amdemod_d_11__N_1841[7]), 
          .S1(amdemod_d_11__N_1841[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1238_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1238_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1238_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1238_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1238_add_4_7 (.A0(amdemod_d_11__N_2017), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2014), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15797), .COUT(n15798), .S0(amdemod_d_11__N_1841[5]), 
          .S1(amdemod_d_11__N_1841[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1238_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1238_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1238_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1238_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1238_add_4_5 (.A0(amdemod_d_11__N_2023), .B0(n17162), .C0(n17279), 
          .D0(n17146), .A1(square_sum[23]), .B1(square_sum[22]), .C1(amdemod_d_11__N_2020), 
          .D1(VCC_net), .CIN(n15796), .COUT(n15797), .S0(amdemod_d_11__N_1841[3]), 
          .S1(amdemod_d_11__N_1841[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1238_add_4_5.INIT0 = 16'h596a;
    defparam _add_1_1238_add_4_5.INIT1 = 16'h1e1e;
    defparam _add_1_1238_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1238_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1238_add_4_3 (.A0(n17134), .B0(square_sum[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(n17134), .B1(amdemod_d_11__N_2026), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15795), .COUT(n15796), .S0(amdemod_d_11__N_1841[1]), 
          .S1(amdemod_d_11__N_1841[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1238_add_4_3.INIT0 = 16'h666a;
    defparam _add_1_1238_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1238_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1238_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1238_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[16]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15795), .S1(amdemod_d_11__N_1841[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1238_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1238_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1238_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1238_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_37 (.A0(integrator4_adj_6023[70]), .B0(cout_adj_5166), 
          .C0(n81_adj_5548), .D0(integrator5_adj_6024[70]), .A1(integrator4_adj_6023[71]), 
          .B1(cout_adj_5166), .C1(n78_adj_5547), .D1(integrator5_adj_6024[71]), 
          .CIN(n15793), .S0(integrator5_71__N_706_adj_6040[70]), .S1(integrator5_71__N_706_adj_6040[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_35 (.A0(integrator4_adj_6023[68]), .B0(cout_adj_5166), 
          .C0(n87_adj_5550), .D0(integrator5_adj_6024[68]), .A1(integrator4_adj_6023[69]), 
          .B1(cout_adj_5166), .C1(n84_adj_5549), .D1(integrator5_adj_6024[69]), 
          .CIN(n15792), .COUT(n15793), .S0(integrator5_71__N_706_adj_6040[68]), 
          .S1(integrator5_71__N_706_adj_6040[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_33 (.A0(integrator4_adj_6023[66]), .B0(cout_adj_5166), 
          .C0(n93_adj_5552), .D0(integrator5_adj_6024[66]), .A1(integrator4_adj_6023[67]), 
          .B1(cout_adj_5166), .C1(n90_adj_5551), .D1(integrator5_adj_6024[67]), 
          .CIN(n15791), .COUT(n15792), .S0(integrator5_71__N_706_adj_6040[66]), 
          .S1(integrator5_71__N_706_adj_6040[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_31 (.A0(integrator4_adj_6023[64]), .B0(cout_adj_5166), 
          .C0(n99_adj_5554), .D0(integrator5_adj_6024[64]), .A1(integrator4_adj_6023[65]), 
          .B1(cout_adj_5166), .C1(n96_adj_5553), .D1(integrator5_adj_6024[65]), 
          .CIN(n15790), .COUT(n15791), .S0(integrator5_71__N_706_adj_6040[64]), 
          .S1(integrator5_71__N_706_adj_6040[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_29 (.A0(integrator4_adj_6023[62]), .B0(cout_adj_5166), 
          .C0(n105_adj_5556), .D0(integrator5_adj_6024[62]), .A1(integrator4_adj_6023[63]), 
          .B1(cout_adj_5166), .C1(n102_adj_5555), .D1(integrator5_adj_6024[63]), 
          .CIN(n15789), .COUT(n15790), .S0(integrator5_71__N_706_adj_6040[62]), 
          .S1(integrator5_71__N_706_adj_6040[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_27 (.A0(integrator4_adj_6023[60]), .B0(cout_adj_5166), 
          .C0(n111_adj_5558), .D0(integrator5_adj_6024[60]), .A1(integrator4_adj_6023[61]), 
          .B1(cout_adj_5166), .C1(n108_adj_5557), .D1(integrator5_adj_6024[61]), 
          .CIN(n15788), .COUT(n15789), .S0(integrator5_71__N_706_adj_6040[60]), 
          .S1(integrator5_71__N_706_adj_6040[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_25 (.A0(integrator4_adj_6023[58]), .B0(cout_adj_5166), 
          .C0(n117_adj_5560), .D0(integrator5_adj_6024[58]), .A1(integrator4_adj_6023[59]), 
          .B1(cout_adj_5166), .C1(n114_adj_5559), .D1(integrator5_adj_6024[59]), 
          .CIN(n15787), .COUT(n15788), .S0(integrator5_71__N_706_adj_6040[58]), 
          .S1(integrator5_71__N_706_adj_6040[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_23 (.A0(integrator4_adj_6023[56]), .B0(cout_adj_5166), 
          .C0(n123_adj_5562), .D0(integrator5_adj_6024[56]), .A1(integrator4_adj_6023[57]), 
          .B1(cout_adj_5166), .C1(n120_adj_5561), .D1(integrator5_adj_6024[57]), 
          .CIN(n15786), .COUT(n15787), .S0(integrator5_71__N_706_adj_6040[56]), 
          .S1(integrator5_71__N_706_adj_6040[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_21 (.A0(integrator4_adj_6023[54]), .B0(cout_adj_5166), 
          .C0(n129_adj_5564), .D0(integrator5_adj_6024[54]), .A1(integrator4_adj_6023[55]), 
          .B1(cout_adj_5166), .C1(n126_adj_5563), .D1(integrator5_adj_6024[55]), 
          .CIN(n15785), .COUT(n15786), .S0(integrator5_71__N_706_adj_6040[54]), 
          .S1(integrator5_71__N_706_adj_6040[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_19 (.A0(integrator4_adj_6023[52]), .B0(cout_adj_5166), 
          .C0(n135_adj_5566), .D0(integrator5_adj_6024[52]), .A1(integrator4_adj_6023[53]), 
          .B1(cout_adj_5166), .C1(n132_adj_5565), .D1(integrator5_adj_6024[53]), 
          .CIN(n15784), .COUT(n15785), .S0(integrator5_71__N_706_adj_6040[52]), 
          .S1(integrator5_71__N_706_adj_6040[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_17 (.A0(integrator4_adj_6023[50]), .B0(cout_adj_5166), 
          .C0(n141_adj_5568), .D0(integrator5_adj_6024[50]), .A1(integrator4_adj_6023[51]), 
          .B1(cout_adj_5166), .C1(n138_adj_5567), .D1(integrator5_adj_6024[51]), 
          .CIN(n15783), .COUT(n15784), .S0(integrator5_71__N_706_adj_6040[50]), 
          .S1(integrator5_71__N_706_adj_6040[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_15 (.A0(integrator4_adj_6023[48]), .B0(cout_adj_5166), 
          .C0(n147_adj_5570), .D0(integrator5_adj_6024[48]), .A1(integrator4_adj_6023[49]), 
          .B1(cout_adj_5166), .C1(n144_adj_5569), .D1(integrator5_adj_6024[49]), 
          .CIN(n15782), .COUT(n15783), .S0(integrator5_71__N_706_adj_6040[48]), 
          .S1(integrator5_71__N_706_adj_6040[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_13 (.A0(integrator4_adj_6023[46]), .B0(cout_adj_5166), 
          .C0(n153_adj_5572), .D0(integrator5_adj_6024[46]), .A1(integrator4_adj_6023[47]), 
          .B1(cout_adj_5166), .C1(n150_adj_5571), .D1(integrator5_adj_6024[47]), 
          .CIN(n15781), .COUT(n15782), .S0(integrator5_71__N_706_adj_6040[46]), 
          .S1(integrator5_71__N_706_adj_6040[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_11 (.A0(integrator4_adj_6023[44]), .B0(cout_adj_5166), 
          .C0(n159_adj_5574), .D0(integrator5_adj_6024[44]), .A1(integrator4_adj_6023[45]), 
          .B1(cout_adj_5166), .C1(n156_adj_5573), .D1(integrator5_adj_6024[45]), 
          .CIN(n15780), .COUT(n15781), .S0(integrator5_71__N_706_adj_6040[44]), 
          .S1(integrator5_71__N_706_adj_6040[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_9 (.A0(integrator4_adj_6023[42]), .B0(cout_adj_5166), 
          .C0(n165_adj_5576), .D0(integrator5_adj_6024[42]), .A1(integrator4_adj_6023[43]), 
          .B1(cout_adj_5166), .C1(n162_adj_5575), .D1(integrator5_adj_6024[43]), 
          .CIN(n15779), .COUT(n15780), .S0(integrator5_71__N_706_adj_6040[42]), 
          .S1(integrator5_71__N_706_adj_6040[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_7 (.A0(integrator4_adj_6023[40]), .B0(cout_adj_5166), 
          .C0(n171_adj_5578), .D0(integrator5_adj_6024[40]), .A1(integrator4_adj_6023[41]), 
          .B1(cout_adj_5166), .C1(n168_adj_5577), .D1(integrator5_adj_6024[41]), 
          .CIN(n15778), .COUT(n15779), .S0(integrator5_71__N_706_adj_6040[40]), 
          .S1(integrator5_71__N_706_adj_6040[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_5 (.A0(integrator4_adj_6023[38]), .B0(cout_adj_5166), 
          .C0(n177_adj_5580), .D0(integrator5_adj_6024[38]), .A1(integrator4_adj_6023[39]), 
          .B1(cout_adj_5166), .C1(n174_adj_5579), .D1(integrator5_adj_6024[39]), 
          .CIN(n15777), .COUT(n15778), .S0(integrator5_71__N_706_adj_6040[38]), 
          .S1(integrator5_71__N_706_adj_6040[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_3 (.A0(integrator4_adj_6023[36]), .B0(cout_adj_5166), 
          .C0(n183_adj_5582), .D0(integrator5_adj_6024[36]), .A1(integrator4_adj_6023[37]), 
          .B1(cout_adj_5166), .C1(n180_adj_5581), .D1(integrator5_adj_6024[37]), 
          .CIN(n15776), .COUT(n15777), .S0(integrator5_71__N_706_adj_6040[36]), 
          .S1(integrator5_71__N_706_adj_6040[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1094_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1094_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1094_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5166), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15776));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1094_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1094_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1094_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1094_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_37 (.A0(comb6[70]), .B0(cout_adj_4985), .C0(n81_adj_5390), 
          .D0(n3), .A1(comb6[71]), .B1(cout_adj_4985), .C1(n78_adj_5389), 
          .D1(n2), .CIN(n15619), .S0(comb7_71__N_1523[70]), .S1(comb7_71__N_1523[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1235_add_4_16 (.A0(amdemod_d_11__N_1840[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15772), .S0(n34_adj_5988));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1235_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1235_add_4_16.INIT1 = 16'h0000;
    defparam _add_1_1235_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1235_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1235_add_4_14 (.A0(amdemod_d_11__N_1840[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1840[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15771), .COUT(n15772), .S0(n40_adj_5989));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1235_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_1235_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_1235_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1235_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1235_add_4_12 (.A0(amdemod_d_11__N_1840[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1840[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15770), .COUT(n15771), .S0(n46_adj_5991), 
          .S1(n43_adj_5990));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1235_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_1235_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_1235_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1235_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1235_add_4_10 (.A0(amdemod_d_11__N_1840[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1840[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15769), .COUT(n15770), .S0(n52_adj_5993), 
          .S1(n49_adj_5992));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1235_add_4_10.INIT0 = 16'h555f;
    defparam _add_1_1235_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_1235_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1235_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_35 (.A0(comb6[68]), .B0(cout_adj_4985), .C0(n87_adj_5392), 
          .D0(n5), .A1(comb6[69]), .B1(cout_adj_4985), .C1(n84_adj_5391), 
          .D1(n4), .CIN(n15618), .COUT(n15619), .S0(comb7_71__N_1523[68]), 
          .S1(comb7_71__N_1523[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1235_add_4_8 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1840[3]), .D0(VCC_net), .A1(amdemod_d_11__N_1840[4]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n15768), .COUT(n15769), 
          .S0(n58_adj_5995), .S1(n55_adj_5994));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1235_add_4_8.INIT0 = 16'he1e1;
    defparam _add_1_1235_add_4_8.INIT1 = 16'h555f;
    defparam _add_1_1235_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1235_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1235_add_4_6 (.A0(n17134), .B0(amdemod_d_11__N_1840[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17137), .B1(amdemod_d_11__N_1840[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15767), .COUT(n15768), .S0(n64_adj_5997), 
          .S1(n61_adj_5996));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1235_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1235_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1235_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1235_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1235_add_4_4 (.A0(n17133), .B0(square_sum[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_d_11__N_1840[0]), .B1(amdemod_d_11__N_1841[11]), 
          .C1(n17134), .D1(amdemod_d_11__N_1840[11]), .CIN(n15766), .COUT(n15767), 
          .S0(n70_adj_5999), .S1(n67_adj_5998));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1235_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1235_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_1235_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1235_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1235_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15766), .S1(n73_adj_6000));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1235_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1235_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1235_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1235_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_37 (.A0(comb8[70]), .B0(cout_adj_5305), .C0(n81_adj_5234), 
          .D0(n3_adj_4803), .A1(comb8[71]), .B1(cout_adj_5305), .C1(n78_adj_5233), 
          .D1(n2_adj_4802), .CIN(n15764), .S0(comb9_71__N_1667[70]), .S1(comb9_71__N_1667[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_35 (.A0(comb8[68]), .B0(cout_adj_5305), .C0(n87_adj_5236), 
          .D0(n5_adj_4805), .A1(comb8[69]), .B1(cout_adj_5305), .C1(n84_adj_5235), 
          .D1(n4_adj_4804), .CIN(n15763), .COUT(n15764), .S0(comb9_71__N_1667[68]), 
          .S1(comb9_71__N_1667[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_33 (.A0(comb8[66]), .B0(cout_adj_5305), .C0(n93_adj_5238), 
          .D0(n7_adj_4807), .A1(comb8[67]), .B1(cout_adj_5305), .C1(n90_adj_5237), 
          .D1(n6_adj_4806), .CIN(n15762), .COUT(n15763), .S0(comb9_71__N_1667[66]), 
          .S1(comb9_71__N_1667[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_33.INJECT1_1 = "NO";
    FD1P3AX phase_inc_gen_i0_i0 (.D(n323), .SP(clk_80mhz_enable_1444), .CK(clk_80mhz), 
            .Q(phase_inc_gen[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i0.GSR = "ENABLED";
    CCU2C _add_1_1073_add_4_31 (.A0(comb8[64]), .B0(cout_adj_5305), .C0(n99_adj_5240), 
          .D0(n9_adj_4809), .A1(comb8[65]), .B1(cout_adj_5305), .C1(n96_adj_5239), 
          .D1(n8_adj_4808), .CIN(n15761), .COUT(n15762), .S0(comb9_71__N_1667[64]), 
          .S1(comb9_71__N_1667[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_29 (.A0(comb8[62]), .B0(cout_adj_5305), .C0(n105_adj_5242), 
          .D0(n11_adj_4811), .A1(comb8[63]), .B1(cout_adj_5305), .C1(n102_adj_5241), 
          .D1(n10_adj_4810), .CIN(n15760), .COUT(n15761), .S0(comb9_71__N_1667[62]), 
          .S1(comb9_71__N_1667[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_27 (.A0(comb8[60]), .B0(cout_adj_5305), .C0(n111_adj_5244), 
          .D0(n13_adj_4813), .A1(comb8[61]), .B1(cout_adj_5305), .C1(n108_adj_5243), 
          .D1(n12_adj_4812), .CIN(n15759), .COUT(n15760), .S0(comb9_71__N_1667[60]), 
          .S1(comb9_71__N_1667[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_25 (.A0(comb8[58]), .B0(cout_adj_5305), .C0(n117_adj_5246), 
          .D0(n15_adj_4815), .A1(comb8[59]), .B1(cout_adj_5305), .C1(n114_adj_5245), 
          .D1(n14_adj_4814), .CIN(n15758), .COUT(n15759), .S0(comb9_71__N_1667[58]), 
          .S1(comb9_71__N_1667[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_23 (.A0(comb8[56]), .B0(cout_adj_5305), .C0(n123_adj_5248), 
          .D0(n17_adj_4817), .A1(comb8[57]), .B1(cout_adj_5305), .C1(n120_adj_5247), 
          .D1(n16_adj_4816), .CIN(n15757), .COUT(n15758), .S0(comb9_71__N_1667[56]), 
          .S1(comb9_71__N_1667[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_21 (.A0(comb8[54]), .B0(cout_adj_5305), .C0(n129_adj_5250), 
          .D0(n19_adj_4819), .A1(comb8[55]), .B1(cout_adj_5305), .C1(n126_adj_5249), 
          .D1(n18_adj_4818), .CIN(n15756), .COUT(n15757), .S0(comb9_71__N_1667[54]), 
          .S1(comb9_71__N_1667[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_19 (.A0(comb8[52]), .B0(cout_adj_5305), .C0(n135_adj_5252), 
          .D0(n21_adj_4821), .A1(comb8[53]), .B1(cout_adj_5305), .C1(n132_adj_5251), 
          .D1(n20_adj_4820), .CIN(n15755), .COUT(n15756), .S0(comb9_71__N_1667[52]), 
          .S1(comb9_71__N_1667[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_33 (.A0(comb6[66]), .B0(cout_adj_4985), .C0(n93_adj_5394), 
          .D0(n7), .A1(comb6[67]), .B1(cout_adj_4985), .C1(n90_adj_5393), 
          .D1(n6), .CIN(n15617), .COUT(n15618), .S0(comb7_71__N_1523[66]), 
          .S1(comb7_71__N_1523[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_31 (.A0(comb6[64]), .B0(cout_adj_4985), .C0(n99_adj_5396), 
          .D0(n9), .A1(comb6[65]), .B1(cout_adj_4985), .C1(n96_adj_5395), 
          .D1(n8), .CIN(n15616), .COUT(n15617), .S0(comb7_71__N_1523[64]), 
          .S1(comb7_71__N_1523[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_29 (.A0(comb6[62]), .B0(cout_adj_4985), .C0(n105_adj_5398), 
          .D0(n11), .A1(comb6[63]), .B1(cout_adj_4985), .C1(n102_adj_5397), 
          .D1(n10), .CIN(n15615), .COUT(n15616), .S0(comb7_71__N_1523[62]), 
          .S1(comb7_71__N_1523[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_27 (.A0(comb6[60]), .B0(cout_adj_4985), .C0(n111_adj_5400), 
          .D0(n13), .A1(comb6[61]), .B1(cout_adj_4985), .C1(n108_adj_5399), 
          .D1(n12), .CIN(n15614), .COUT(n15615), .S0(comb7_71__N_1523[60]), 
          .S1(comb7_71__N_1523[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_25 (.A0(comb6[58]), .B0(cout_adj_4985), .C0(n117_adj_5402), 
          .D0(n15), .A1(comb6[59]), .B1(cout_adj_4985), .C1(n114_adj_5401), 
          .D1(n14), .CIN(n15613), .COUT(n15614), .S0(comb7_71__N_1523[58]), 
          .S1(comb7_71__N_1523[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_23 (.A0(comb6[56]), .B0(cout_adj_4985), .C0(n123_adj_5404), 
          .D0(n17), .A1(comb6[57]), .B1(cout_adj_4985), .C1(n120_adj_5403), 
          .D1(n16_adj_2947), .CIN(n15612), .COUT(n15613), .S0(comb7_71__N_1523[56]), 
          .S1(comb7_71__N_1523[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_21 (.A0(comb6[54]), .B0(cout_adj_4985), .C0(n129_adj_5406), 
          .D0(n19), .A1(comb6[55]), .B1(cout_adj_4985), .C1(n126_adj_5405), 
          .D1(n18), .CIN(n15611), .COUT(n15612), .S0(comb7_71__N_1523[54]), 
          .S1(comb7_71__N_1523[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_19 (.A0(comb6[52]), .B0(cout_adj_4985), .C0(n135_adj_5408), 
          .D0(n21), .A1(comb6[53]), .B1(cout_adj_4985), .C1(n132_adj_5407), 
          .D1(n20), .CIN(n15610), .COUT(n15611), .S0(comb7_71__N_1523[52]), 
          .S1(comb7_71__N_1523[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_17 (.A0(comb6[50]), .B0(cout_adj_4985), .C0(n141_adj_5410), 
          .D0(n23), .A1(comb6[51]), .B1(cout_adj_4985), .C1(n138_adj_5409), 
          .D1(n22), .CIN(n15609), .COUT(n15610), .S0(comb7_71__N_1523[50]), 
          .S1(comb7_71__N_1523[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_17 (.A0(comb8[50]), .B0(cout_adj_5305), .C0(n141_adj_5254), 
          .D0(n23_adj_4823), .A1(comb8[51]), .B1(cout_adj_5305), .C1(n138_adj_5253), 
          .D1(n22_adj_4822), .CIN(n15754), .COUT(n15755), .S0(comb9_71__N_1667[50]), 
          .S1(comb9_71__N_1667[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_15 (.A0(comb8[48]), .B0(cout_adj_5305), .C0(n147_adj_5256), 
          .D0(n25_adj_4825), .A1(comb8[49]), .B1(cout_adj_5305), .C1(n144_adj_5255), 
          .D1(n24_adj_4824), .CIN(n15753), .COUT(n15754), .S0(comb9_71__N_1667[48]), 
          .S1(comb9_71__N_1667[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_13 (.A0(comb8[46]), .B0(cout_adj_5305), .C0(n153_adj_5258), 
          .D0(n27_adj_4827), .A1(comb8[47]), .B1(cout_adj_5305), .C1(n150_adj_5257), 
          .D1(n26_adj_4826), .CIN(n15752), .COUT(n15753), .S0(comb9_71__N_1667[46]), 
          .S1(comb9_71__N_1667[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_11 (.A0(comb8[44]), .B0(cout_adj_5305), .C0(n159_adj_5260), 
          .D0(n29_adj_4829), .A1(comb8[45]), .B1(cout_adj_5305), .C1(n156_adj_5259), 
          .D1(n28_adj_4828), .CIN(n15751), .COUT(n15752), .S0(comb9_71__N_1667[44]), 
          .S1(comb9_71__N_1667[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_9 (.A0(comb8[42]), .B0(cout_adj_5305), .C0(n165_adj_5262), 
          .D0(n31_adj_4831), .A1(comb8[43]), .B1(cout_adj_5305), .C1(n162_adj_5261), 
          .D1(n30_adj_4830), .CIN(n15750), .COUT(n15751), .S0(comb9_71__N_1667[42]), 
          .S1(comb9_71__N_1667[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_15 (.A0(comb6[48]), .B0(cout_adj_4985), .C0(n147_adj_5412), 
          .D0(n25), .A1(comb6[49]), .B1(cout_adj_4985), .C1(n144_adj_5411), 
          .D1(n24), .CIN(n15608), .COUT(n15609), .S0(comb7_71__N_1523[48]), 
          .S1(comb7_71__N_1523[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_15.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_24 (.A0(phase_inc_gen1[22]), .B0(phase_accum[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[23]), .B1(phase_accum[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15480), .COUT(n15481), .S0(n255), 
          .S1(n252));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_24.INIT0 = 16'h666a;
    defparam phase_accum_add_4_24.INIT1 = 16'h666a;
    defparam phase_accum_add_4_24.INJECT1_0 = "NO";
    defparam phase_accum_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_7 (.A0(comb8[40]), .B0(cout_adj_5305), .C0(n171_adj_5264), 
          .D0(n33_adj_4833), .A1(comb8[41]), .B1(cout_adj_5305), .C1(n168_adj_5263), 
          .D1(n32_adj_4832), .CIN(n15749), .COUT(n15750), .S0(comb9_71__N_1667[40]), 
          .S1(comb9_71__N_1667[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_5 (.A0(comb8[38]), .B0(cout_adj_5305), .C0(n177_adj_5266), 
          .D0(n35_adj_4835), .A1(comb8[39]), .B1(cout_adj_5305), .C1(n174_adj_5265), 
          .D1(n34_adj_4834), .CIN(n15748), .COUT(n15749), .S0(comb9_71__N_1667[38]), 
          .S1(comb9_71__N_1667[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_3 (.A0(comb8[36]), .B0(cout_adj_5305), .C0(n183_adj_5268), 
          .D0(n37_adj_4837), .A1(comb8[37]), .B1(cout_adj_5305), .C1(n180_adj_5267), 
          .D1(n36_adj_4836), .CIN(n15747), .COUT(n15748), .S0(comb9_71__N_1667[36]), 
          .S1(comb9_71__N_1667[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1073_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1073_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1073_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5305), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15747));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1073_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1073_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1073_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1073_add_4_1.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_22 (.A0(phase_inc_gen1[20]), .B0(phase_accum[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[21]), .B1(phase_accum[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15479), .COUT(n15480), .S0(n261), 
          .S1(n258));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_22.INIT0 = 16'h666a;
    defparam phase_accum_add_4_22.INIT1 = 16'h666a;
    defparam phase_accum_add_4_22.INJECT1_0 = "NO";
    defparam phase_accum_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1229_add_4_16 (.A0(amdemod_d_11__N_1850[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15743), .S0(n34_adj_5975));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1229_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1229_add_4_16.INIT1 = 16'h0000;
    defparam _add_1_1229_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1229_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1229_add_4_14 (.A0(amdemod_d_11__N_1850[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1850[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15742), .COUT(n15743), .S0(n40_adj_5976));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1229_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_1229_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_1229_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1229_add_4_14.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_20 (.A0(phase_inc_gen1[18]), .B0(phase_accum[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[19]), .B1(phase_accum[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15478), .COUT(n15479), .S0(n267), 
          .S1(n264));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_20.INIT0 = 16'h666a;
    defparam phase_accum_add_4_20.INIT1 = 16'h666a;
    defparam phase_accum_add_4_20.INJECT1_0 = "NO";
    defparam phase_accum_add_4_20.INJECT1_1 = "NO";
    LUT4 i4704_2_lut (.A(integrator3[0]), .B(integrator2[0]), .Z(integrator3_71__N_562[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4704_2_lut.init = 16'h6666;
    CCU2C _add_1_1193_add_4_4 (.A0(n17130), .B0(square_sum[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(n17130), .B1(amdemod_d_11__N_2170), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15284), .COUT(n15285), .S0(amdemod_d_11__N_1860[1]), 
          .S1(amdemod_d_11__N_1860[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1193_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1193_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1193_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1193_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1193_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15284), .S1(amdemod_d_11__N_1860[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1193_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1193_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1193_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1193_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1262_add_4_14 (.A0(n17134), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15283), .S0(amdemod_d_11__N_1840[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1262_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_1262_add_4_14.INIT1 = 16'h0000;
    defparam _add_1_1262_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1262_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_10 (.A0(integrator3_adj_6022[8]), .B0(integrator2_adj_6021[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[9]), .B1(integrator2_adj_6021[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14937), .COUT(n14938), .S0(integrator3_71__N_562_adj_6038[8]), 
          .S1(integrator3_71__N_562_adj_6038[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_8 (.A0(integrator3_adj_6022[6]), .B0(integrator2_adj_6021[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[7]), .B1(integrator2_adj_6021[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14936), .COUT(n14937), .S0(integrator3_71__N_562_adj_6038[6]), 
          .S1(integrator3_71__N_562_adj_6038[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_6 (.A0(integrator3_adj_6022[4]), .B0(integrator2_adj_6021[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[5]), .B1(integrator2_adj_6021[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14935), .COUT(n14936), .S0(integrator3_71__N_562_adj_6038[4]), 
          .S1(integrator3_71__N_562_adj_6038[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_4 (.A0(integrator3_adj_6022[2]), .B0(integrator2_adj_6021[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[3]), .B1(integrator2_adj_6021[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14934), .COUT(n14935), .S0(integrator3_71__N_562_adj_6038[2]), 
          .S1(integrator3_71__N_562_adj_6038[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1002_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1002_add_4_2 (.A0(integrator3_adj_6022[0]), .B0(integrator2_adj_6021[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[1]), .B1(integrator2_adj_6021[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14934), .S1(integrator3_71__N_562_adj_6038[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1002_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1002_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1002_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1002_add_4_2.INJECT1_1 = "NO";
    LUT4 i1651_3_lut_4_lut (.A(n17288), .B(n17150), .C(n17289), .D(n175), 
         .Z(n11373)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1651_3_lut_4_lut.init = 16'hf707;
    CCU2C _add_1_1005_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14932), .S0(cout_adj_5165));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1005_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1005_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_36 (.A0(integrator4_adj_6023[34]), .B0(integrator3_adj_6022[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[35]), .B1(integrator3_adj_6022[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14931), .COUT(n14932), .S0(integrator4_71__N_634_adj_6039[34]), 
          .S1(integrator4_71__N_634_adj_6039[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_34 (.A0(integrator4_adj_6023[32]), .B0(integrator3_adj_6022[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[33]), .B1(integrator3_adj_6022[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14930), .COUT(n14931), .S0(integrator4_71__N_634_adj_6039[32]), 
          .S1(integrator4_71__N_634_adj_6039[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_32 (.A0(integrator4_adj_6023[30]), .B0(integrator3_adj_6022[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[31]), .B1(integrator3_adj_6022[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14929), .COUT(n14930), .S0(integrator4_71__N_634_adj_6039[30]), 
          .S1(integrator4_71__N_634_adj_6039[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_30 (.A0(integrator4_adj_6023[28]), .B0(integrator3_adj_6022[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[29]), .B1(integrator3_adj_6022[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14928), .COUT(n14929), .S0(integrator4_71__N_634_adj_6039[28]), 
          .S1(integrator4_71__N_634_adj_6039[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_28 (.A0(integrator4_adj_6023[26]), .B0(integrator3_adj_6022[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[27]), .B1(integrator3_adj_6022[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14927), .COUT(n14928), .S0(integrator4_71__N_634_adj_6039[26]), 
          .S1(integrator4_71__N_634_adj_6039[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_26 (.A0(integrator4_adj_6023[24]), .B0(integrator3_adj_6022[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[25]), .B1(integrator3_adj_6022[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14926), .COUT(n14927), .S0(integrator4_71__N_634_adj_6039[24]), 
          .S1(integrator4_71__N_634_adj_6039[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_24 (.A0(integrator4_adj_6023[22]), .B0(integrator3_adj_6022[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[23]), .B1(integrator3_adj_6022[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14925), .COUT(n14926), .S0(integrator4_71__N_634_adj_6039[22]), 
          .S1(integrator4_71__N_634_adj_6039[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_22 (.A0(integrator4_adj_6023[20]), .B0(integrator3_adj_6022[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[21]), .B1(integrator3_adj_6022[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14924), .COUT(n14925), .S0(integrator4_71__N_634_adj_6039[20]), 
          .S1(integrator4_71__N_634_adj_6039[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_20 (.A0(integrator4_adj_6023[18]), .B0(integrator3_adj_6022[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[19]), .B1(integrator3_adj_6022[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14923), .COUT(n14924), .S0(integrator4_71__N_634_adj_6039[18]), 
          .S1(integrator4_71__N_634_adj_6039[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_18 (.A0(integrator4_adj_6023[16]), .B0(integrator3_adj_6022[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[17]), .B1(integrator3_adj_6022[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14922), .COUT(n14923), .S0(integrator4_71__N_634_adj_6039[16]), 
          .S1(integrator4_71__N_634_adj_6039[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_16 (.A0(integrator4_adj_6023[14]), .B0(integrator3_adj_6022[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[15]), .B1(integrator3_adj_6022[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14921), .COUT(n14922), .S0(integrator4_71__N_634_adj_6039[14]), 
          .S1(integrator4_71__N_634_adj_6039[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_14 (.A0(integrator4_adj_6023[12]), .B0(integrator3_adj_6022[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[13]), .B1(integrator3_adj_6022[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14920), .COUT(n14921), .S0(integrator4_71__N_634_adj_6039[12]), 
          .S1(integrator4_71__N_634_adj_6039[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_12 (.A0(integrator4_adj_6023[10]), .B0(integrator3_adj_6022[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[11]), .B1(integrator3_adj_6022[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14919), .COUT(n14920), .S0(integrator4_71__N_634_adj_6039[10]), 
          .S1(integrator4_71__N_634_adj_6039[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_10 (.A0(integrator4_adj_6023[8]), .B0(integrator3_adj_6022[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[9]), .B1(integrator3_adj_6022[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14918), .COUT(n14919), .S0(integrator4_71__N_634_adj_6039[8]), 
          .S1(integrator4_71__N_634_adj_6039[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_8 (.A0(integrator4_adj_6023[6]), .B0(integrator3_adj_6022[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[7]), .B1(integrator3_adj_6022[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14917), .COUT(n14918), .S0(integrator4_71__N_634_adj_6039[6]), 
          .S1(integrator4_71__N_634_adj_6039[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_6 (.A0(integrator4_adj_6023[4]), .B0(integrator3_adj_6022[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[5]), .B1(integrator3_adj_6022[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14916), .COUT(n14917), .S0(integrator4_71__N_634_adj_6039[4]), 
          .S1(integrator4_71__N_634_adj_6039[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_4 (.A0(integrator4_adj_6023[2]), .B0(integrator3_adj_6022[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[3]), .B1(integrator3_adj_6022[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14915), .COUT(n14916), .S0(integrator4_71__N_634_adj_6039[2]), 
          .S1(integrator4_71__N_634_adj_6039[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1005_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1005_add_4_2 (.A0(integrator4_adj_6023[0]), .B0(integrator3_adj_6022[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[1]), .B1(integrator3_adj_6022[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14915), .S1(integrator4_71__N_634_adj_6039[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1005_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1005_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1005_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1005_add_4_2.INJECT1_1 = "NO";
    LUT4 i4703_2_lut (.A(integrator4[0]), .B(integrator3[0]), .Z(integrator4_71__N_634[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4703_2_lut.init = 16'h6666;
    CCU2C _add_1_1008_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14913), .S0(cout_adj_5166));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1008_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1008_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_36 (.A0(integrator5_adj_6024[34]), .B0(integrator4_adj_6023[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[35]), .B1(integrator4_adj_6023[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14912), .COUT(n14913), .S0(integrator5_71__N_706_adj_6040[34]), 
          .S1(integrator5_71__N_706_adj_6040[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_34 (.A0(integrator5_adj_6024[32]), .B0(integrator4_adj_6023[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[33]), .B1(integrator4_adj_6023[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14911), .COUT(n14912), .S0(integrator5_71__N_706_adj_6040[32]), 
          .S1(integrator5_71__N_706_adj_6040[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_32 (.A0(integrator5_adj_6024[30]), .B0(integrator4_adj_6023[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[31]), .B1(integrator4_adj_6023[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14910), .COUT(n14911), .S0(integrator5_71__N_706_adj_6040[30]), 
          .S1(integrator5_71__N_706_adj_6040[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_30 (.A0(integrator5_adj_6024[28]), .B0(integrator4_adj_6023[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[29]), .B1(integrator4_adj_6023[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14909), .COUT(n14910), .S0(integrator5_71__N_706_adj_6040[28]), 
          .S1(integrator5_71__N_706_adj_6040[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_28 (.A0(integrator5_adj_6024[26]), .B0(integrator4_adj_6023[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[27]), .B1(integrator4_adj_6023[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14908), .COUT(n14909), .S0(integrator5_71__N_706_adj_6040[26]), 
          .S1(integrator5_71__N_706_adj_6040[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_26 (.A0(integrator5_adj_6024[24]), .B0(integrator4_adj_6023[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[25]), .B1(integrator4_adj_6023[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14907), .COUT(n14908), .S0(integrator5_71__N_706_adj_6040[24]), 
          .S1(integrator5_71__N_706_adj_6040[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_24 (.A0(integrator5_adj_6024[22]), .B0(integrator4_adj_6023[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[23]), .B1(integrator4_adj_6023[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14906), .COUT(n14907), .S0(integrator5_71__N_706_adj_6040[22]), 
          .S1(integrator5_71__N_706_adj_6040[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_22 (.A0(integrator5_adj_6024[20]), .B0(integrator4_adj_6023[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[21]), .B1(integrator4_adj_6023[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14905), .COUT(n14906), .S0(integrator5_71__N_706_adj_6040[20]), 
          .S1(integrator5_71__N_706_adj_6040[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_20 (.A0(integrator5_adj_6024[18]), .B0(integrator4_adj_6023[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[19]), .B1(integrator4_adj_6023[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14904), .COUT(n14905), .S0(integrator5_71__N_706_adj_6040[18]), 
          .S1(integrator5_71__N_706_adj_6040[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_18 (.A0(integrator5_adj_6024[16]), .B0(integrator4_adj_6023[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[17]), .B1(integrator4_adj_6023[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14903), .COUT(n14904), .S0(integrator5_71__N_706_adj_6040[16]), 
          .S1(integrator5_71__N_706_adj_6040[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_16 (.A0(integrator5_adj_6024[14]), .B0(integrator4_adj_6023[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[15]), .B1(integrator4_adj_6023[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14902), .COUT(n14903), .S0(integrator5_71__N_706_adj_6040[14]), 
          .S1(integrator5_71__N_706_adj_6040[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_14 (.A0(integrator5_adj_6024[12]), .B0(integrator4_adj_6023[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[13]), .B1(integrator4_adj_6023[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14901), .COUT(n14902), .S0(integrator5_71__N_706_adj_6040[12]), 
          .S1(integrator5_71__N_706_adj_6040[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_12 (.A0(integrator5_adj_6024[10]), .B0(integrator4_adj_6023[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[11]), .B1(integrator4_adj_6023[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14900), .COUT(n14901), .S0(integrator5_71__N_706_adj_6040[10]), 
          .S1(integrator5_71__N_706_adj_6040[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_10 (.A0(integrator5_adj_6024[8]), .B0(integrator4_adj_6023[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[9]), .B1(integrator4_adj_6023[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14899), .COUT(n14900), .S0(integrator5_71__N_706_adj_6040[8]), 
          .S1(integrator5_71__N_706_adj_6040[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_8 (.A0(integrator5_adj_6024[6]), .B0(integrator4_adj_6023[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[7]), .B1(integrator4_adj_6023[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14898), .COUT(n14899), .S0(integrator5_71__N_706_adj_6040[6]), 
          .S1(integrator5_71__N_706_adj_6040[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_6 (.A0(integrator5_adj_6024[4]), .B0(integrator4_adj_6023[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[5]), .B1(integrator4_adj_6023[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14897), .COUT(n14898), .S0(integrator5_71__N_706_adj_6040[4]), 
          .S1(integrator5_71__N_706_adj_6040[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_4 (.A0(integrator5_adj_6024[2]), .B0(integrator4_adj_6023[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[3]), .B1(integrator4_adj_6023[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14896), .COUT(n14897), .S0(integrator5_71__N_706_adj_6040[2]), 
          .S1(integrator5_71__N_706_adj_6040[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1008_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1008_add_4_2 (.A0(integrator5_adj_6024[0]), .B0(integrator4_adj_6023[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[1]), .B1(integrator4_adj_6023[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14896), .S1(integrator5_71__N_706_adj_6040[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1008_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1008_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1008_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1008_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_37 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n81_adj_5354), .D0(integrator1[70]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n78_adj_5353), .D1(integrator1[71]), 
          .CIN(n14893), .S0(integrator1_71__N_418[70]), .S1(integrator1_71__N_418[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_35 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n87_adj_5356), .D0(integrator1[68]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n84_adj_5355), .D1(integrator1[69]), 
          .CIN(n14892), .COUT(n14893), .S0(integrator1_71__N_418[68]), 
          .S1(integrator1_71__N_418[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_33 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n93_adj_5358), .D0(integrator1[66]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n90_adj_5357), .D1(integrator1[67]), 
          .CIN(n14891), .COUT(n14892), .S0(integrator1_71__N_418[66]), 
          .S1(integrator1_71__N_418[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_31 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n99_adj_5360), .D0(integrator1[64]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n96_adj_5359), .D1(integrator1[65]), 
          .CIN(n14890), .COUT(n14891), .S0(integrator1_71__N_418[64]), 
          .S1(integrator1_71__N_418[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_29 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n105_adj_5362), .D0(integrator1[62]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n102_adj_5361), .D1(integrator1[63]), 
          .CIN(n14889), .COUT(n14890), .S0(integrator1_71__N_418[62]), 
          .S1(integrator1_71__N_418[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_27 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n111_adj_5364), .D0(integrator1[60]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n108_adj_5363), .D1(integrator1[61]), 
          .CIN(n14888), .COUT(n14889), .S0(integrator1_71__N_418[60]), 
          .S1(integrator1_71__N_418[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_25 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n117_adj_5366), .D0(integrator1[58]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n114_adj_5365), .D1(integrator1[59]), 
          .CIN(n14887), .COUT(n14888), .S0(integrator1_71__N_418[58]), 
          .S1(integrator1_71__N_418[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_23 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n123_adj_5368), .D0(integrator1[56]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n120_adj_5367), .D1(integrator1[57]), 
          .CIN(n14886), .COUT(n14887), .S0(integrator1_71__N_418[56]), 
          .S1(integrator1_71__N_418[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_21 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n129_adj_5370), .D0(integrator1[54]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n126_adj_5369), .D1(integrator1[55]), 
          .CIN(n14885), .COUT(n14886), .S0(integrator1_71__N_418[54]), 
          .S1(integrator1_71__N_418[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_19 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n135_adj_5372), .D0(integrator1[52]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n132_adj_5371), .D1(integrator1[53]), 
          .CIN(n14884), .COUT(n14885), .S0(integrator1_71__N_418[52]), 
          .S1(integrator1_71__N_418[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_17 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n141_adj_5374), .D0(integrator1[50]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n138_adj_5373), .D1(integrator1[51]), 
          .CIN(n14883), .COUT(n14884), .S0(integrator1_71__N_418[50]), 
          .S1(integrator1_71__N_418[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_15 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n147_adj_5376), .D0(integrator1[48]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n144_adj_5375), .D1(integrator1[49]), 
          .CIN(n14882), .COUT(n14883), .S0(integrator1_71__N_418[48]), 
          .S1(integrator1_71__N_418[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_13 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n153_adj_5378), .D0(integrator1[46]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n150_adj_5377), .D1(integrator1[47]), 
          .CIN(n14881), .COUT(n14882), .S0(integrator1_71__N_418[46]), 
          .S1(integrator1_71__N_418[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_11 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n159_adj_5380), .D0(integrator1[44]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n156_adj_5379), .D1(integrator1[45]), 
          .CIN(n14880), .COUT(n14881), .S0(integrator1_71__N_418[44]), 
          .S1(integrator1_71__N_418[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_9 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n165_adj_5382), .D0(integrator1[42]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n162_adj_5381), .D1(integrator1[43]), 
          .CIN(n14879), .COUT(n14880), .S0(integrator1_71__N_418[42]), 
          .S1(integrator1_71__N_418[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_7 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n171_adj_5384), .D0(integrator1[40]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n168_adj_5383), .D1(integrator1[41]), 
          .CIN(n14878), .COUT(n14879), .S0(integrator1_71__N_418[40]), 
          .S1(integrator1_71__N_418[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_5 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n177_adj_5386), .D0(integrator1[38]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n174_adj_5385), .D1(integrator1[39]), 
          .CIN(n14877), .COUT(n14878), .S0(integrator1_71__N_418[38]), 
          .S1(integrator1_71__N_418[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_3 (.A0(mix_sinewave[11]), .B0(cout_adj_5126), 
          .C0(n183_adj_5388), .D0(integrator1[36]), .A1(mix_sinewave[11]), 
          .B1(cout_adj_5126), .C1(n180_adj_5387), .D1(integrator1[37]), 
          .CIN(n14876), .COUT(n14877), .S0(integrator1_71__N_418[36]), 
          .S1(integrator1_71__N_418[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1011_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1011_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1011_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5126), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14876));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1011_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1011_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1011_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1011_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1014_add_4_13 (.A0(count_adj_6035[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14872), .S0(n28_adj_5167));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_1014_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1014_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_1014_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1014_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1014_add_4_11 (.A0(count_adj_6035[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_6035[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14871), .COUT(n14872), .S0(n34_adj_5169), 
          .S1(n31_adj_5168));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_1014_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1014_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1014_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1014_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1014_add_4_9 (.A0(count_adj_6035[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_6035[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14870), .COUT(n14871), .S0(n40_adj_5171), 
          .S1(n37_adj_5170));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_1014_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1014_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1014_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1014_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_13 (.A0(comb6[46]), .B0(cout_adj_4985), .C0(n153_adj_5414), 
          .D0(n27_adj_2946), .A1(comb6[47]), .B1(cout_adj_4985), .C1(n150_adj_5413), 
          .D1(n26), .CIN(n15607), .COUT(n15608), .S0(comb7_71__N_1523[46]), 
          .S1(comb7_71__N_1523[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_11 (.A0(comb6[44]), .B0(cout_adj_4985), .C0(n159_adj_5416), 
          .D0(n29), .A1(comb6[45]), .B1(cout_adj_4985), .C1(n156_adj_5415), 
          .D1(n28), .CIN(n15606), .COUT(n15607), .S0(comb7_71__N_1523[44]), 
          .S1(comb7_71__N_1523[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_9 (.A0(comb6[42]), .B0(cout_adj_4985), .C0(n165_adj_5418), 
          .D0(n31), .A1(comb6[43]), .B1(cout_adj_4985), .C1(n162_adj_5417), 
          .D1(n30), .CIN(n15605), .COUT(n15606), .S0(comb7_71__N_1523[42]), 
          .S1(comb7_71__N_1523[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_7 (.A0(comb6[40]), .B0(cout_adj_4985), .C0(n171_adj_5420), 
          .D0(n33), .A1(comb6[41]), .B1(cout_adj_4985), .C1(n168_adj_5419), 
          .D1(n32), .CIN(n15604), .COUT(n15605), .S0(comb7_71__N_1523[40]), 
          .S1(comb7_71__N_1523[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_5 (.A0(comb6[38]), .B0(cout_adj_4985), .C0(n177_adj_5422), 
          .D0(n35), .A1(comb6[39]), .B1(cout_adj_4985), .C1(n174_adj_5421), 
          .D1(n34), .CIN(n15603), .COUT(n15604), .S0(comb7_71__N_1523[38]), 
          .S1(comb7_71__N_1523[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_5.INJECT1_1 = "NO";
    LUT4 i4702_2_lut (.A(integrator5[0]), .B(integrator4[0]), .Z(integrator5_71__N_706[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4702_2_lut.init = 16'h6666;
    CCU2C _add_1_1067_add_4_3 (.A0(comb6[36]), .B0(cout_adj_4985), .C0(n183_adj_5424), 
          .D0(n37), .A1(comb6[37]), .B1(cout_adj_4985), .C1(n180_adj_5423), 
          .D1(n36), .CIN(n15602), .COUT(n15603), .S0(comb7_71__N_1523[36]), 
          .S1(comb7_71__N_1523[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1067_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1067_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1067_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_4985), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15602));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1067_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1067_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1067_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1067_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_15 (.A0(amdemod_d_11__N_1860[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15598), .S0(n32_adj_5863));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1064_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1064_add_4_15.INIT1 = 16'h0000;
    defparam _add_1_1064_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_13 (.A0(amdemod_d_11__N_1860[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1860[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15597), .COUT(n15598), .S0(n38_adj_5864));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1064_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1064_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1064_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_11 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1860[7]), .D0(VCC_net), .A1(amdemod_d_11__N_1860[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n15596), .COUT(n15597), 
          .S0(n44_adj_5866), .S1(n41_adj_5865));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1064_add_4_11.INIT0 = 16'h1e1e;
    defparam _add_1_1064_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1064_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_9 (.A0(n17134), .B0(amdemod_d_11__N_1860[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1860[6]), .B1(n17162), 
          .C1(n17279), .D1(n17146), .CIN(n15595), .COUT(n15596), .S0(n50_adj_5868), 
          .S1(n47_adj_5867));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1064_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1064_add_4_9.INIT1 = 16'h596a;
    defparam _add_1_1064_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_7 (.A0(n17132), .B0(amdemod_d_11__N_1860[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17133), .B1(amdemod_d_11__N_1860[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15594), .COUT(n15595), .S0(n56_adj_5870), 
          .S1(n53_adj_5869));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1064_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1064_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1064_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_5 (.A0(n17130), .B0(amdemod_d_11__N_1860[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17131), .B1(amdemod_d_11__N_1860[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15593), .COUT(n15594), .S0(n62_adj_5872), 
          .S1(n59_adj_5871));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1064_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1064_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1064_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_3 (.A0(square_sum[7]), .B0(amdemod_d_11__N_1861[13]), 
          .C0(n17130), .D0(amdemod_d_11__N_1860[13]), .A1(n17129), .B1(amdemod_d_11__N_1860[0]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15592), .COUT(n15593), .S0(n68_adj_5874), 
          .S1(n65_adj_5873));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1064_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_1064_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1064_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1064_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15592), .S1(n71_adj_5875));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1064_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1064_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1064_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1064_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_37 (.A0(comb_d9[71]), .B0(comb9[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15591), .S0(n76_adj_5848));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_37.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_37.INIT1 = 16'h0000;
    defparam _add_1_1076_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_35 (.A0(comb_d9[69]), .B0(comb9[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[70]), .B1(comb9[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15590), .COUT(n15591), .S0(n82_adj_5850), 
          .S1(n79_adj_5849));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_35.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_35.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_33 (.A0(comb_d9[67]), .B0(comb9[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[68]), .B1(comb9[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15589), .COUT(n15590), .S0(n88_adj_5852), 
          .S1(n85_adj_5851));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_33.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_33.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_31 (.A0(comb_d9[65]), .B0(comb9[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[66]), .B1(comb9[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15588), .COUT(n15589), .S0(n94_adj_5854), 
          .S1(n91_adj_5853));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_31.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_31.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_29 (.A0(comb_d9[63]), .B0(comb9[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[64]), .B1(comb9[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15587), .COUT(n15588), .S0(n100_adj_5856), 
          .S1(n97_adj_5855));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_29.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_29.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_27 (.A0(comb_d9[61]), .B0(comb9[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[62]), .B1(comb9[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15586), .COUT(n15587), .S0(n106_adj_5858), 
          .S1(n103_adj_5857));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_27.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_27.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_25 (.A0(comb_d9[59]), .B0(comb9[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[60]), .B1(comb9[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15585), .COUT(n15586), .S0(n112_adj_5860), 
          .S1(n109_adj_5859));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_25.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_25.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_23 (.A0(comb_d9[57]), .B0(comb9[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[58]), .B1(comb9[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15584), .COUT(n15585), .S0(n118_adj_5862), 
          .S1(n115_adj_5861));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_23.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_23.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_21 (.A0(comb_d9[55]), .B0(comb9[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[56]), .B1(comb9[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15583), .COUT(n15584));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_21.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_21.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_19 (.A0(comb_d9[53]), .B0(comb9[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[54]), .B1(comb9[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15582), .COUT(n15583));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_19.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_19.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_17 (.A0(comb_d9[51]), .B0(comb9[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[52]), .B1(comb9[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15581), .COUT(n15582));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_17.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_17.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_15 (.A0(comb_d9[49]), .B0(comb9[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[50]), .B1(comb9[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15580), .COUT(n15581));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_15.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_15.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_13 (.A0(comb_d9[47]), .B0(comb9[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[48]), .B1(comb9[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15579), .COUT(n15580));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_13.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_13.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_11 (.A0(comb_d9[45]), .B0(comb9[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[46]), .B1(comb9[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15578), .COUT(n15579));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_9 (.A0(comb_d9[43]), .B0(comb9[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[44]), .B1(comb9[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15577), .COUT(n15578));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_7 (.A0(comb_d9[41]), .B0(comb9[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[42]), .B1(comb9[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15576), .COUT(n15577));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_5 (.A0(comb_d9[39]), .B0(comb9[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[40]), .B1(comb9[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15575), .COUT(n15576));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1076_add_4_3 (.A0(comb_d9[37]), .B0(comb9[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[38]), .B1(comb9[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15574), .COUT(n15575));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_1076_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_3.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_4_lut (.A(led_c_0), .B(led_c_1), .C(n17289), .D(led_c_2), 
         .Z(n16245)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'hfffd;
    CCU2C _add_1_1076_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[36]), .B1(comb9[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15574));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1076_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1076_add_4_1.INIT1 = 16'h9995;
    defparam _add_1_1076_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1076_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1232_add_4_16 (.A0(amdemod_d_11__N_1841[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15573), .S0(n34_adj_5835));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1232_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1232_add_4_16.INIT1 = 16'h0000;
    defparam _add_1_1232_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1232_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1232_add_4_14 (.A0(amdemod_d_11__N_1841[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1841[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15572), .COUT(n15573), .S0(n40_adj_5836));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1232_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_1232_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_1232_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1232_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1232_add_4_12 (.A0(amdemod_d_11__N_1841[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1841[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15571), .COUT(n15572), .S0(n46_adj_5838), 
          .S1(n43_adj_5837));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1232_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_1232_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_1232_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1232_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1232_add_4_10 (.A0(amdemod_d_11__N_1841[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1841[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15570), .COUT(n15571), .S0(n52_adj_5840), 
          .S1(n49_adj_5839));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1232_add_4_10.INIT0 = 16'h555f;
    defparam _add_1_1232_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_1232_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1232_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1232_add_4_8 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1841[3]), .D0(VCC_net), .A1(amdemod_d_11__N_1841[4]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n15569), .COUT(n15570), 
          .S0(n58_adj_5842), .S1(n55_adj_5841));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1232_add_4_8.INIT0 = 16'he1e1;
    defparam _add_1_1232_add_4_8.INIT1 = 16'h555f;
    defparam _add_1_1232_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1232_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1232_add_4_6 (.A0(n17134), .B0(amdemod_d_11__N_1841[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17137), .B1(amdemod_d_11__N_1841[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15568), .COUT(n15569), .S0(n64_adj_5844), 
          .S1(n61_adj_5843));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1232_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1232_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1232_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1232_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1232_add_4_4 (.A0(n17133), .B0(square_sum[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_d_11__N_1841[0]), .B1(amdemod_d_11__N_1841[11]), 
          .C1(n17134), .D1(amdemod_d_11__N_1840[11]), .CIN(n15567), .COUT(n15568), 
          .S0(n70_adj_5846), .S1(n67_adj_5845));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1232_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1232_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_1232_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1232_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1232_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15567), .S1(n73_adj_5847));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1232_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1232_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1232_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1232_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_38 (.A0(integrator3[71]), .B0(integrator2[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15566), .S0(n78_adj_5311));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1181_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_36 (.A0(integrator3[69]), .B0(integrator2[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[70]), .B1(integrator2[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15565), .COUT(n15566), .S0(n84_adj_5313), 
          .S1(n81_adj_5312));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_34 (.A0(integrator3[67]), .B0(integrator2[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[68]), .B1(integrator2[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15564), .COUT(n15565), .S0(n90_adj_5315), 
          .S1(n87_adj_5314));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_32 (.A0(integrator3[65]), .B0(integrator2[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[66]), .B1(integrator2[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15563), .COUT(n15564), .S0(n96_adj_5317), 
          .S1(n93_adj_5316));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_30 (.A0(integrator3[63]), .B0(integrator2[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[64]), .B1(integrator2[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15562), .COUT(n15563), .S0(n102_adj_5319), 
          .S1(n99_adj_5318));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_28 (.A0(integrator3[61]), .B0(integrator2[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[62]), .B1(integrator2[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15561), .COUT(n15562), .S0(n108_adj_5321), 
          .S1(n105_adj_5320));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_26 (.A0(integrator3[59]), .B0(integrator2[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[60]), .B1(integrator2[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15560), .COUT(n15561), .S0(n114_adj_5323), 
          .S1(n111_adj_5322));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_24 (.A0(integrator3[57]), .B0(integrator2[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[58]), .B1(integrator2[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15559), .COUT(n15560), .S0(n120_adj_5325), 
          .S1(n117_adj_5324));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_22 (.A0(integrator3[55]), .B0(integrator2[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[56]), .B1(integrator2[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15558), .COUT(n15559), .S0(n126_adj_5327), 
          .S1(n123_adj_5326));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_20 (.A0(integrator3[53]), .B0(integrator2[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[54]), .B1(integrator2[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15557), .COUT(n15558), .S0(n132_adj_5329), 
          .S1(n129_adj_5328));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_18 (.A0(integrator3[51]), .B0(integrator2[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[52]), .B1(integrator2[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15556), .COUT(n15557), .S0(n138_adj_5331), 
          .S1(n135_adj_5330));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1229_add_4_12 (.A0(amdemod_d_11__N_1850[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1850[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15741), .COUT(n15742), .S0(n46_adj_5978), 
          .S1(n43_adj_5977));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1229_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_1229_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_1229_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1229_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1229_add_4_10 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1850[5]), .D0(VCC_net), .A1(amdemod_d_11__N_1850[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n15740), .COUT(n15741), 
          .S0(n52_adj_5980), .S1(n49_adj_5979));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1229_add_4_10.INIT0 = 16'he1e1;
    defparam _add_1_1229_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_1229_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1229_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1262_add_4_12 (.A0(amdemod_d_11__N_2005), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(n17134), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15282), .COUT(n15283), .S0(amdemod_d_11__N_1840[9]), 
          .S1(amdemod_d_11__N_1840[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1262_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_1262_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_1262_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1262_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1262_add_4_10 (.A0(amdemod_d_11__N_2011), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2008), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15281), .COUT(n15282), .S0(amdemod_d_11__N_1840[7]), 
          .S1(amdemod_d_11__N_1840[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1262_add_4_10.INIT0 = 16'h555f;
    defparam _add_1_1262_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_1262_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1262_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1262_add_4_8 (.A0(amdemod_d_11__N_2017), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2014), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15280), .COUT(n15281), .S0(amdemod_d_11__N_1840[5]), 
          .S1(amdemod_d_11__N_1840[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1262_add_4_8.INIT0 = 16'h555f;
    defparam _add_1_1262_add_4_8.INIT1 = 16'h555f;
    defparam _add_1_1262_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1262_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1262_add_4_6 (.A0(n17137), .B0(amdemod_d_11__N_2023), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[23]), .B1(square_sum[22]), .C1(amdemod_d_11__N_2020), 
          .D1(VCC_net), .CIN(n15279), .COUT(n15280), .S0(amdemod_d_11__N_1840[3]), 
          .S1(amdemod_d_11__N_1840[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1262_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1262_add_4_6.INIT1 = 16'he1e1;
    defparam _add_1_1262_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1262_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1262_add_4_4 (.A0(n17134), .B0(square_sum[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(n17134), .B1(amdemod_d_11__N_2026), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15278), .COUT(n15279), .S0(amdemod_d_11__N_1840[1]), 
          .S1(amdemod_d_11__N_1840[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1262_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1262_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1262_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1262_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1262_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[16]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15278), .S1(amdemod_d_11__N_1840[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1262_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1262_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1262_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1262_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_38 (.A0(integrator4[71]), .B0(integrator3[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15277), .S0(n78_adj_5089));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1265_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_36 (.A0(integrator4[69]), .B0(integrator3[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[70]), .B1(integrator3[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15276), .COUT(n15277), .S0(n84_adj_5091), 
          .S1(n81_adj_5090));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_34 (.A0(integrator4[67]), .B0(integrator3[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[68]), .B1(integrator3[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15275), .COUT(n15276), .S0(n90_adj_5093), 
          .S1(n87_adj_5092));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_32 (.A0(integrator4[65]), .B0(integrator3[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[66]), .B1(integrator3[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15274), .COUT(n15275), .S0(n96_adj_5095), 
          .S1(n93_adj_5094));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_30 (.A0(integrator4[63]), .B0(integrator3[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[64]), .B1(integrator3[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15273), .COUT(n15274), .S0(n102_adj_5097), 
          .S1(n99_adj_5096));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_28 (.A0(integrator4[61]), .B0(integrator3[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[62]), .B1(integrator3[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15272), .COUT(n15273), .S0(n108_adj_5099), 
          .S1(n105_adj_5098));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_26 (.A0(integrator4[59]), .B0(integrator3[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[60]), .B1(integrator3[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15271), .COUT(n15272), .S0(n114_adj_5101), 
          .S1(n111_adj_5100));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_24 (.A0(integrator4[57]), .B0(integrator3[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[58]), .B1(integrator3[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15270), .COUT(n15271), .S0(n120_adj_5103), 
          .S1(n117_adj_5102));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_22 (.A0(integrator4[55]), .B0(integrator3[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[56]), .B1(integrator3[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15269), .COUT(n15270), .S0(n126_adj_5105), 
          .S1(n123_adj_5104));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_20 (.A0(integrator4[53]), .B0(integrator3[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[54]), .B1(integrator3[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15268), .COUT(n15269), .S0(n132_adj_5107), 
          .S1(n129_adj_5106));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_20.INJECT1_1 = "NO";
    FD1S3AX square_sum_e1_i0_i1 (.D(n79), .CK(cic_sine_clk), .Q(n46_adj_5700));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i1.GSR = "ENABLED";
    CCU2C _add_1_1014_add_4_7 (.A0(count_adj_6035[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_6035[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14869), .COUT(n14870), .S0(n46_adj_5173), 
          .S1(n43_adj_5172));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_1014_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1014_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1014_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1014_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1014_add_4_5 (.A0(count_adj_6035[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_6035[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14868), .COUT(n14869), .S0(n52_adj_5175), 
          .S1(n49_adj_5174));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_1014_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1014_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1014_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1014_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1014_add_4_3 (.A0(count_adj_6035[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count_adj_6035[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14867), .COUT(n14868), .S0(n58_adj_5177), 
          .S1(n55_adj_5176));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_1014_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1014_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1014_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1014_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1014_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_adj_6035[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14867), .S1(n61_adj_5178));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(83[25:34])
    defparam _add_1_1014_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1014_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1014_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1014_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_37 (.A0(integrator1[70]), .B0(cout_adj_5072), 
          .C0(n81), .D0(integrator2[70]), .A1(integrator1[71]), .B1(cout_adj_5072), 
          .C1(n78_adj_4984), .D1(integrator2[71]), .CIN(n14865), .S0(integrator2_71__N_490[70]), 
          .S1(integrator2_71__N_490[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_35 (.A0(integrator1[68]), .B0(cout_adj_5072), 
          .C0(n87), .D0(integrator2[68]), .A1(integrator1[69]), .B1(cout_adj_5072), 
          .C1(n84), .D1(integrator2[69]), .CIN(n14864), .COUT(n14865), 
          .S0(integrator2_71__N_490[68]), .S1(integrator2_71__N_490[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_33 (.A0(integrator1[66]), .B0(cout_adj_5072), 
          .C0(n93), .D0(integrator2[66]), .A1(integrator1[67]), .B1(cout_adj_5072), 
          .C1(n90), .D1(integrator2[67]), .CIN(n14863), .COUT(n14864), 
          .S0(integrator2_71__N_490[66]), .S1(integrator2_71__N_490[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_31 (.A0(integrator1[64]), .B0(cout_adj_5072), 
          .C0(n99), .D0(integrator2[64]), .A1(integrator1[65]), .B1(cout_adj_5072), 
          .C1(n96), .D1(integrator2[65]), .CIN(n14862), .COUT(n14863), 
          .S0(integrator2_71__N_490[64]), .S1(integrator2_71__N_490[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_29 (.A0(integrator1[62]), .B0(cout_adj_5072), 
          .C0(n105), .D0(integrator2[62]), .A1(integrator1[63]), .B1(cout_adj_5072), 
          .C1(n102), .D1(integrator2[63]), .CIN(n14861), .COUT(n14862), 
          .S0(integrator2_71__N_490[62]), .S1(integrator2_71__N_490[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_27 (.A0(integrator1[60]), .B0(cout_adj_5072), 
          .C0(n111), .D0(integrator2[60]), .A1(integrator1[61]), .B1(cout_adj_5072), 
          .C1(n108), .D1(integrator2[61]), .CIN(n14860), .COUT(n14861), 
          .S0(integrator2_71__N_490[60]), .S1(integrator2_71__N_490[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_25 (.A0(integrator1[58]), .B0(cout_adj_5072), 
          .C0(n117), .D0(integrator2[58]), .A1(integrator1[59]), .B1(cout_adj_5072), 
          .C1(n114), .D1(integrator2[59]), .CIN(n14859), .COUT(n14860), 
          .S0(integrator2_71__N_490[58]), .S1(integrator2_71__N_490[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_23 (.A0(integrator1[56]), .B0(cout_adj_5072), 
          .C0(n123), .D0(integrator2[56]), .A1(integrator1[57]), .B1(cout_adj_5072), 
          .C1(n120), .D1(integrator2[57]), .CIN(n14858), .COUT(n14859), 
          .S0(integrator2_71__N_490[56]), .S1(integrator2_71__N_490[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_21 (.A0(integrator1[54]), .B0(cout_adj_5072), 
          .C0(n129), .D0(integrator2[54]), .A1(integrator1[55]), .B1(cout_adj_5072), 
          .C1(n126), .D1(integrator2[55]), .CIN(n14857), .COUT(n14858), 
          .S0(integrator2_71__N_490[54]), .S1(integrator2_71__N_490[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_19 (.A0(integrator1[52]), .B0(cout_adj_5072), 
          .C0(n135), .D0(integrator2[52]), .A1(integrator1[53]), .B1(cout_adj_5072), 
          .C1(n132), .D1(integrator2[53]), .CIN(n14856), .COUT(n14857), 
          .S0(integrator2_71__N_490[52]), .S1(integrator2_71__N_490[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_17 (.A0(integrator1[50]), .B0(cout_adj_5072), 
          .C0(n141), .D0(integrator2[50]), .A1(integrator1[51]), .B1(cout_adj_5072), 
          .C1(n138), .D1(integrator2[51]), .CIN(n14855), .COUT(n14856), 
          .S0(integrator2_71__N_490[50]), .S1(integrator2_71__N_490[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_15 (.A0(integrator1[48]), .B0(cout_adj_5072), 
          .C0(n147), .D0(integrator2[48]), .A1(integrator1[49]), .B1(cout_adj_5072), 
          .C1(n144), .D1(integrator2[49]), .CIN(n14854), .COUT(n14855), 
          .S0(integrator2_71__N_490[48]), .S1(integrator2_71__N_490[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_13 (.A0(integrator1[46]), .B0(cout_adj_5072), 
          .C0(n153), .D0(integrator2[46]), .A1(integrator1[47]), .B1(cout_adj_5072), 
          .C1(n150), .D1(integrator2[47]), .CIN(n14853), .COUT(n14854), 
          .S0(integrator2_71__N_490[46]), .S1(integrator2_71__N_490[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_11 (.A0(integrator1[44]), .B0(cout_adj_5072), 
          .C0(n159), .D0(integrator2[44]), .A1(integrator1[45]), .B1(cout_adj_5072), 
          .C1(n156), .D1(integrator2[45]), .CIN(n14852), .COUT(n14853), 
          .S0(integrator2_71__N_490[44]), .S1(integrator2_71__N_490[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_9 (.A0(integrator1[42]), .B0(cout_adj_5072), 
          .C0(n165), .D0(integrator2[42]), .A1(integrator1[43]), .B1(cout_adj_5072), 
          .C1(n162), .D1(integrator2[43]), .CIN(n14851), .COUT(n14852), 
          .S0(integrator2_71__N_490[42]), .S1(integrator2_71__N_490[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_7 (.A0(integrator1[40]), .B0(cout_adj_5072), 
          .C0(n171), .D0(integrator2[40]), .A1(integrator1[41]), .B1(cout_adj_5072), 
          .C1(n168), .D1(integrator2[41]), .CIN(n14850), .COUT(n14851), 
          .S0(integrator2_71__N_490[40]), .S1(integrator2_71__N_490[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_5 (.A0(integrator1[38]), .B0(cout_adj_5072), 
          .C0(n177), .D0(integrator2[38]), .A1(integrator1[39]), .B1(cout_adj_5072), 
          .C1(n174), .D1(integrator2[39]), .CIN(n14849), .COUT(n14850), 
          .S0(integrator2_71__N_490[38]), .S1(integrator2_71__N_490[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_3 (.A0(integrator1[36]), .B0(cout_adj_5072), 
          .C0(n183), .D0(integrator2[36]), .A1(integrator1[37]), .B1(cout_adj_5072), 
          .C1(n180), .D1(integrator2[37]), .CIN(n14848), .COUT(n14849), 
          .S0(integrator2_71__N_490[36]), .S1(integrator2_71__N_490[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1017_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1017_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1017_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5072), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14848));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1017_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1017_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1017_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1017_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1049_add_4_9 (.A0(n17162), .B0(n17146), .C0(GND_net), 
          .D0(VCC_net), .A1(n17162), .B1(n17146), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14835), .S0(n25_adj_5180), .S1(n22_adj_5179));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1049_add_4_9.INIT0 = 16'h1111;
    defparam _add_1_1049_add_4_9.INIT1 = 16'h1111;
    defparam _add_1_1049_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1049_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1229_add_4_8 (.A0(n17134), .B0(amdemod_d_11__N_1850[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17137), .B1(amdemod_d_11__N_1850[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15739), .COUT(n15740), .S0(n58_adj_5982), 
          .S1(n55_adj_5981));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1229_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1229_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1229_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1229_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1229_add_4_6 (.A0(n17132), .B0(amdemod_d_11__N_1850[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1850[2]), .B1(amdemod_d_11__N_1841[11]), 
          .C1(n17134), .D1(amdemod_d_11__N_1840[11]), .CIN(n15738), .COUT(n15739), 
          .S0(n64_adj_5984), .S1(n61_adj_5983));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1229_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1229_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_1229_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1229_add_4_6.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_18 (.A0(phase_inc_gen1[16]), .B0(phase_accum[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[17]), .B1(phase_accum[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15477), .COUT(n15478), .S0(n273), 
          .S1(n270));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_18.INIT0 = 16'h666a;
    defparam phase_accum_add_4_18.INIT1 = 16'h666a;
    defparam phase_accum_add_4_18.INJECT1_0 = "NO";
    defparam phase_accum_add_4_18.INJECT1_1 = "NO";
    LUT4 i1888_4_lut (.A(n133_adj_5905), .B(n127), .C(led_c_3), .D(n17144), 
         .Z(n11622)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1888_4_lut.init = 16'hcac0;
    CCU2C _add_1_1229_add_4_4 (.A0(n17131), .B0(square_sum[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_d_11__N_1850[0]), .B1(amdemod_d_11__N_1851[13]), 
          .C1(n17132), .D1(amdemod_d_11__N_1850[13]), .CIN(n15737), .COUT(n15738), 
          .S0(n70_adj_5986), .S1(n67_adj_5985));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1229_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1229_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_1229_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1229_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1229_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15737), .S1(n73_adj_5987));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1229_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1229_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1229_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1229_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_37 (.A0(integrator_tmp[70]), .B0(cout), .C0(n81_adj_5426), 
          .D0(n3_adj_2961), .A1(integrator_tmp[71]), .B1(cout), .C1(n78_adj_5425), 
          .D1(n2_adj_2962), .CIN(n15735), .S0(comb6_71__N_1451[70]), .S1(comb6_71__N_1451[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_37.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_16 (.A0(phase_inc_gen1[14]), .B0(phase_accum[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[15]), .B1(phase_accum[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15476), .COUT(n15477), .S0(n279), 
          .S1(n276));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_16.INIT0 = 16'h666a;
    defparam phase_accum_add_4_16.INIT1 = 16'h666a;
    defparam phase_accum_add_4_16.INJECT1_0 = "NO";
    defparam phase_accum_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_35 (.A0(integrator_tmp[68]), .B0(cout), .C0(n87_adj_5428), 
          .D0(n5_adj_2959), .A1(integrator_tmp[69]), .B1(cout), .C1(n84_adj_5427), 
          .D1(n4_adj_2960), .CIN(n15734), .COUT(n15735), .S0(comb6_71__N_1451[68]), 
          .S1(comb6_71__N_1451[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_33 (.A0(integrator_tmp[66]), .B0(cout), .C0(n93_adj_5430), 
          .D0(n7_adj_2957), .A1(integrator_tmp[67]), .B1(cout), .C1(n90_adj_5429), 
          .D1(n6_adj_2958), .CIN(n15733), .COUT(n15734), .S0(comb6_71__N_1451[66]), 
          .S1(comb6_71__N_1451[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_31 (.A0(integrator_tmp[64]), .B0(cout), .C0(n99_adj_5432), 
          .D0(n9_adj_2955), .A1(integrator_tmp[65]), .B1(cout), .C1(n96_adj_5431), 
          .D1(n8_adj_2956), .CIN(n15732), .COUT(n15733), .S0(comb6_71__N_1451[64]), 
          .S1(comb6_71__N_1451[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_29 (.A0(integrator_tmp[62]), .B0(cout), .C0(n105_adj_5434), 
          .D0(n11_adj_2953), .A1(integrator_tmp[63]), .B1(cout), .C1(n102_adj_5433), 
          .D1(n10_adj_2954), .CIN(n15731), .COUT(n15732), .S0(comb6_71__N_1451[62]), 
          .S1(comb6_71__N_1451[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1250_add_4_5 (.A0(n17132), .B0(amdemod_d_11__N_1850[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17133), .B1(amdemod_d_11__N_1850[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15463), .COUT(n15464), .S0(n62), 
          .S1(n59));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1250_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1250_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1250_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1250_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_16 (.A0(integrator3[49]), .B0(integrator2[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[50]), .B1(integrator2[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15555), .COUT(n15556), .S0(n144_adj_5333), 
          .S1(n141_adj_5332));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_27 (.A0(integrator_tmp[60]), .B0(cout), .C0(n111_adj_5436), 
          .D0(n13_adj_2951), .A1(integrator_tmp[61]), .B1(cout), .C1(n108_adj_5435), 
          .D1(n12_adj_2952), .CIN(n15730), .COUT(n15731), .S0(comb6_71__N_1451[60]), 
          .S1(comb6_71__N_1451[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_25 (.A0(integrator_tmp[58]), .B0(cout), .C0(n117_adj_5438), 
          .D0(n15_adj_2949), .A1(integrator_tmp[59]), .B1(cout), .C1(n114_adj_5437), 
          .D1(n14_adj_2950), .CIN(n15729), .COUT(n15730), .S0(comb6_71__N_1451[58]), 
          .S1(comb6_71__N_1451[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_23 (.A0(integrator_tmp[56]), .B0(cout), .C0(n123_adj_5440), 
          .D0(n17_adj_4763), .A1(integrator_tmp[57]), .B1(cout), .C1(n120_adj_5439), 
          .D1(n16), .CIN(n15728), .COUT(n15729), .S0(comb6_71__N_1451[56]), 
          .S1(comb6_71__N_1451[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_21 (.A0(integrator_tmp[54]), .B0(cout), .C0(n129_adj_5442), 
          .D0(n19_adj_4748), .A1(integrator_tmp[55]), .B1(cout), .C1(n126_adj_5441), 
          .D1(n18_adj_4761), .CIN(n15727), .COUT(n15728), .S0(comb6_71__N_1451[54]), 
          .S1(comb6_71__N_1451[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1190_add_4_10 (.A0(amdemod_d_11__N_2083), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2080), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15341), .COUT(n15342), .S0(amdemod_d_11__N_1850[7]), 
          .S1(amdemod_d_11__N_1850[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1190_add_4_10.INIT0 = 16'h555f;
    defparam _add_1_1190_add_4_10.INIT1 = 16'h555f;
    defparam _add_1_1190_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1190_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_19 (.A0(integrator_tmp[52]), .B0(cout), .C0(n135_adj_5444), 
          .D0(n21_adj_4743), .A1(integrator_tmp[53]), .B1(cout), .C1(n132_adj_5443), 
          .D1(n20_adj_4744), .CIN(n15726), .COUT(n15727), .S0(comb6_71__N_1451[52]), 
          .S1(comb6_71__N_1451[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_17 (.A0(integrator_tmp[50]), .B0(cout), .C0(n141_adj_5446), 
          .D0(n23_adj_4727), .A1(integrator_tmp[51]), .B1(cout), .C1(n138_adj_5445), 
          .D1(n22_adj_4728), .CIN(n15725), .COUT(n15726), .S0(comb6_71__N_1451[50]), 
          .S1(comb6_71__N_1451[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_15 (.A0(integrator_tmp[48]), .B0(cout), .C0(n147_adj_5448), 
          .D0(n25_adj_2974), .A1(integrator_tmp[49]), .B1(cout), .C1(n144_adj_5447), 
          .D1(n24_adj_4716), .CIN(n15724), .COUT(n15725), .S0(comb6_71__N_1451[48]), 
          .S1(comb6_71__N_1451[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_13 (.A0(integrator_tmp[46]), .B0(cout), .C0(n153_adj_5450), 
          .D0(n27), .A1(integrator_tmp[47]), .B1(cout), .C1(n150_adj_5449), 
          .D1(n26_adj_2973), .CIN(n15723), .COUT(n15724), .S0(comb6_71__N_1451[46]), 
          .S1(comb6_71__N_1451[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_11 (.A0(integrator_tmp[44]), .B0(cout), .C0(n159_adj_5452), 
          .D0(n29_adj_2971), .A1(integrator_tmp[45]), .B1(cout), .C1(n156_adj_5451), 
          .D1(n28_adj_2972), .CIN(n15722), .COUT(n15723), .S0(comb6_71__N_1451[44]), 
          .S1(comb6_71__N_1451[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_9 (.A0(integrator_tmp[42]), .B0(cout), .C0(n165_adj_5454), 
          .D0(n31_adj_2969), .A1(integrator_tmp[43]), .B1(cout), .C1(n162_adj_5453), 
          .D1(n30_adj_2970), .CIN(n15721), .COUT(n15722), .S0(comb6_71__N_1451[42]), 
          .S1(comb6_71__N_1451[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_7 (.A0(integrator_tmp[40]), .B0(cout), .C0(n171_adj_5456), 
          .D0(n33_adj_2967), .A1(integrator_tmp[41]), .B1(cout), .C1(n168_adj_5455), 
          .D1(n32_adj_2968), .CIN(n15720), .COUT(n15721), .S0(comb6_71__N_1451[40]), 
          .S1(comb6_71__N_1451[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_5 (.A0(integrator_tmp[38]), .B0(cout), .C0(n177_adj_5458), 
          .D0(n35_adj_2965), .A1(integrator_tmp[39]), .B1(cout), .C1(n174_adj_5457), 
          .D1(n34_adj_2966), .CIN(n15719), .COUT(n15720), .S0(comb6_71__N_1451[38]), 
          .S1(comb6_71__N_1451[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_3 (.A0(integrator_tmp[36]), .B0(cout), .C0(n183_adj_5460), 
          .D0(n37_adj_2963), .A1(integrator_tmp[37]), .B1(cout), .C1(n180_adj_5459), 
          .D1(n36_adj_2964), .CIN(n15718), .COUT(n15719), .S0(comb6_71__N_1451[36]), 
          .S1(comb6_71__N_1451[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1040_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1040_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1190_add_4_12 (.A0(amdemod_d_11__N_2077), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2074), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15342), .COUT(n15343), .S0(amdemod_d_11__N_1850[9]), 
          .S1(amdemod_d_11__N_1850[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1190_add_4_12.INIT0 = 16'h555f;
    defparam _add_1_1190_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_1190_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1190_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1040_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15718));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1040_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1040_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1040_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1040_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1247_add_4_15 (.A0(amdemod_d_11__N_1851[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15714), .S0(n32_adj_5962));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1247_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1247_add_4_15.INIT1 = 16'h0000;
    defparam _add_1_1247_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1247_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1247_add_4_13 (.A0(amdemod_d_11__N_1851[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1851[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15713), .COUT(n15714), .S0(n38_adj_5963));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1247_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1247_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1247_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1247_add_4_13.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_14 (.A0(phase_inc_gen1[12]), .B0(phase_accum[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[13]), .B1(phase_accum[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15475), .COUT(n15476), .S0(n285), 
          .S1(n282));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_14.INIT0 = 16'h666a;
    defparam phase_accum_add_4_14.INIT1 = 16'h666a;
    defparam phase_accum_add_4_14.INJECT1_0 = "NO";
    defparam phase_accum_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1247_add_4_11 (.A0(amdemod_d_11__N_1851[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1851[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15712), .COUT(n15713), .S0(n44_adj_5965), 
          .S1(n41_adj_5964));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1247_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1247_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1247_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1247_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1247_add_4_9 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1851[5]), .D0(VCC_net), .A1(amdemod_d_11__N_1851[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n15711), .COUT(n15712), 
          .S0(n50_adj_5967), .S1(n47_adj_5966));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1247_add_4_9.INIT0 = 16'h1e1e;
    defparam _add_1_1247_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1247_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1247_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1247_add_4_7 (.A0(n17134), .B0(amdemod_d_11__N_1851[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1851[4]), .B1(n17162), 
          .C1(n17279), .D1(n17146), .CIN(n15710), .COUT(n15711), .S0(n56_adj_5969), 
          .S1(n53_adj_5968));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1247_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1247_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_1247_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1247_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1247_add_4_5 (.A0(n17132), .B0(amdemod_d_11__N_1851[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17133), .B1(amdemod_d_11__N_1851[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15709), .COUT(n15710), .S0(n62_adj_5971), 
          .S1(n59_adj_5970));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1247_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1247_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1247_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1247_add_4_5.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_12 (.A0(phase_inc_gen1[10]), .B0(phase_accum[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[11]), .B1(phase_accum[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15474), .COUT(n15475), .S0(n291), 
          .S1(n288));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_12.INIT0 = 16'h666a;
    defparam phase_accum_add_4_12.INIT1 = 16'h666a;
    defparam phase_accum_add_4_12.INJECT1_0 = "NO";
    defparam phase_accum_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1247_add_4_3 (.A0(square_sum[11]), .B0(amdemod_d_11__N_1851[13]), 
          .C0(n17132), .D0(amdemod_d_11__N_1850[13]), .A1(n17131), .B1(amdemod_d_11__N_1851[0]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15708), .COUT(n15709), .S0(n68_adj_5973), 
          .S1(n65_adj_5972));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1247_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_1247_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1247_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1247_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1247_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15708), .S1(n71_adj_5974));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1247_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1247_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1247_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1247_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_63 (.A0(phase_inc_gen[62]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[63]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15706), .S0(n133_adj_5905), .S1(n130_adj_5904));
    defparam _add_1_1244_add_4_63.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_63.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_63.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_63.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_61 (.A0(phase_inc_gen[60]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[61]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15705), .COUT(n15706), .S0(n139_adj_5907), 
          .S1(n136_adj_5906));
    defparam _add_1_1244_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_61.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_61.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_10 (.A0(phase_inc_gen1[8]), .B0(phase_accum[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[9]), .B1(phase_accum[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15473), .COUT(n15474), .S0(n297), 
          .S1(n294));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_10.INIT0 = 16'h666a;
    defparam phase_accum_add_4_10.INIT1 = 16'h666a;
    defparam phase_accum_add_4_10.INJECT1_0 = "NO";
    defparam phase_accum_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_59 (.A0(phase_inc_gen[58]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[59]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15704), .COUT(n15705), .S0(n145_adj_5909), 
          .S1(n142_adj_5908));
    defparam _add_1_1244_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_59.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_14 (.A0(integrator3[47]), .B0(integrator2[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[48]), .B1(integrator2[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15554), .COUT(n15555), .S0(n150_adj_5335), 
          .S1(n147_adj_5334));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_57 (.A0(phase_inc_gen[56]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[57]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15703), .COUT(n15704), .S0(n151_adj_5911), 
          .S1(n148_adj_5910));
    defparam _add_1_1244_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_55 (.A0(phase_inc_gen[54]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[55]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15702), .COUT(n15703), .S0(n157_adj_5913), 
          .S1(n154_adj_5912));
    defparam _add_1_1244_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_53 (.A0(phase_inc_gen[52]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[53]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15701), .COUT(n15702), .S0(n163_adj_5915), 
          .S1(n160_adj_5914));
    defparam _add_1_1244_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_51 (.A0(phase_inc_gen[50]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[51]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15700), .COUT(n15701), .S0(n169_adj_5917), 
          .S1(n166_adj_5916));
    defparam _add_1_1244_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_51.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_49 (.A0(phase_inc_gen[48]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[49]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15699), .COUT(n15700), .S0(n175_adj_5919), 
          .S1(n172_adj_5918));
    defparam _add_1_1244_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_49.INJECT1_1 = "NO";
    CCU2C _add_1_1250_add_4_11 (.A0(amdemod_d_11__N_1850[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1850[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15466), .COUT(n15467), .S0(n44), 
          .S1(n41));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1250_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1250_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1250_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1250_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_47 (.A0(phase_inc_gen[46]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[47]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15698), .COUT(n15699), .S0(n181_adj_5921), 
          .S1(n178_adj_5920));
    defparam _add_1_1244_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_1244_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_45 (.A0(phase_inc_gen[44]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[45]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15697), .COUT(n15698), .S0(n187_adj_5923), 
          .S1(n184_adj_5922));
    defparam _add_1_1244_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_45.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_43 (.A0(phase_inc_gen[42]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[43]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15696), .COUT(n15697), .S0(n193_adj_5925), 
          .S1(n190_adj_5924));
    defparam _add_1_1244_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_43.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_41 (.A0(phase_inc_gen[40]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[41]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15695), .COUT(n15696), .S0(n199_adj_5927), 
          .S1(n196_adj_5926));
    defparam _add_1_1244_add_4_41.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_1190_add_4_14 (.A0(amdemod_d_11__N_2071), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2068), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15343), .COUT(n15344), .S0(amdemod_d_11__N_1850[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1190_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_1190_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_1190_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1190_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_12 (.A0(integrator3[45]), .B0(integrator2[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[46]), .B1(integrator2[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15553), .COUT(n15554), .S0(n156_adj_5337), 
          .S1(n153_adj_5336));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_39 (.A0(phase_inc_gen[38]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[39]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15694), .COUT(n15695), .S0(n205_adj_5929), 
          .S1(n202_adj_5928));
    defparam _add_1_1244_add_4_39.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_39.INJECT1_1 = "NO";
    CCU2C _add_1_1190_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15338), .S1(amdemod_d_11__N_1850[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1190_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1190_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1190_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1190_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_18 (.A0(integrator4[51]), .B0(integrator3[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[52]), .B1(integrator3[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15267), .COUT(n15268), .S0(n138_adj_5109), 
          .S1(n135_adj_5108));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_18.INJECT1_1 = "NO";
    FD1S3AX square_sum_e1_i0_i2 (.D(n78), .CK(cic_sine_clk), .Q(n44_adj_5699));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i2.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i3 (.D(n77), .CK(cic_sine_clk), .Q(n42_adj_5698));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i3.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i4 (.D(n76), .CK(cic_sine_clk), .Q(n40_adj_5697));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i4.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i5 (.D(n75), .CK(cic_sine_clk), .Q(n38_adj_5696));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i5.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i6 (.D(n74), .CK(cic_sine_clk), .Q(n36_adj_5695));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i6.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i7 (.D(n73), .CK(cic_sine_clk), .Q(n34_adj_5694));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i7.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i8 (.D(n72), .CK(cic_sine_clk), .Q(n32_adj_5693));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i8.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i9 (.D(n71_adj_4749), .CK(cic_sine_clk), .Q(n30_adj_5692));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i9.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i10 (.D(n70), .CK(cic_sine_clk), .Q(n28_adj_5691));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i10.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i11 (.D(n69), .CK(cic_sine_clk), .Q(n26_adj_5690));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i11.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i12 (.D(n68_adj_4750), .CK(cic_sine_clk), .Q(n24_adj_5689));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i12.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i13 (.D(n67), .CK(cic_sine_clk), .Q(n22_adj_5688));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i13.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i14 (.D(n66_adj_4752), .CK(cic_sine_clk), .Q(n20_adj_5687));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i14.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i15 (.D(n65_adj_4753), .CK(cic_sine_clk), .Q(n18_adj_5686));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i15.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i16 (.D(n64_adj_4754), .CK(cic_sine_clk), .Q(n16_adj_5685));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i16.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i17 (.D(n63_adj_4755), .CK(cic_sine_clk), .Q(n14_adj_5684));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i17.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i18 (.D(n62_adj_4756), .CK(cic_sine_clk), .Q(n12_adj_5683));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i18.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i19 (.D(n61), .CK(cic_sine_clk), .Q(n10_adj_5682));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i19.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i20 (.D(n60), .CK(cic_sine_clk), .Q(n8_adj_5681));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i20.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i21 (.D(n59_adj_4758), .CK(cic_sine_clk), .Q(n6_adj_5680));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i21.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i22 (.D(n58), .CK(cic_sine_clk), .Q(n4_adj_5679));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i22.GSR = "ENABLED";
    FD1S3AX square_sum_e1_i0_i23 (.D(n57), .CK(cic_sine_clk), .Q(n2_adj_5678));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_e1_i0_i23.GSR = "ENABLED";
    CCU2C _add_1_1049_add_4_7 (.A0(n17157), .B0(n17163), .C0(GND_net), 
          .D0(VCC_net), .A1(n17162), .B1(n17146), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14834), .COUT(n14835), .S0(n31_adj_5182), .S1(n28_adj_5181));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1049_add_4_7.INIT0 = 16'h9999;
    defparam _add_1_1049_add_4_7.INIT1 = 16'h9999;
    defparam _add_1_1049_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1049_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1049_add_4_5 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1830[1]), .D0(VCC_net), .A1(n11179), .B1(n4_adj_4982), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14833), .COUT(n14834), .S0(n37_adj_5184), 
          .S1(n34_adj_5183));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1049_add_4_5.INIT0 = 16'he1ee;
    defparam _add_1_1049_add_4_5.INIT1 = 16'h6666;
    defparam _add_1_1049_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1049_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1049_add_4_3 (.A0(n17137), .B0(square_sum[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[20]), .B1(n17279), .C1(n17162), 
          .D1(n17146), .CIN(n14832), .COUT(n14833), .S0(n43_adj_5186), 
          .S1(n40_adj_5185));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1049_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_1049_add_4_3.INIT1 = 16'h9a95;
    defparam _add_1_1049_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1049_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1049_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[18]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14832), .S1(n46_adj_5187));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1049_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1049_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1049_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1049_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1199_add_4_16 (.A0(amdemod_d_11__N_2281), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14831), .S0(amdemod_d_11__N_1880[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1199_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1199_add_4_16.INIT1 = 16'h0000;
    defparam _add_1_1199_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1199_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1199_add_4_14 (.A0(n17137), .B0(amdemod_d_11__N_2287), 
          .C0(GND_net), .D0(VCC_net), .A1(square_sum[23]), .B1(square_sum[22]), 
          .C1(amdemod_d_11__N_2284), .D1(VCC_net), .CIN(n14830), .COUT(n14831));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1199_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1199_add_4_14.INIT1 = 16'he1e1;
    defparam _add_1_1199_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1199_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1199_add_4_12 (.A0(amdemod_d_11__N_2293), .B0(amdemod_d_11__N_1841[11]), 
          .C0(n17134), .D0(amdemod_d_11__N_1840[11]), .A1(n17134), .B1(amdemod_d_11__N_2290), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14829), .COUT(n14830));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1199_add_4_12.INIT0 = 16'h656a;
    defparam _add_1_1199_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1199_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1199_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1199_add_4_10 (.A0(amdemod_d_11__N_2299), .B0(amdemod_d_11__N_1851[13]), 
          .C0(n17132), .D0(amdemod_d_11__N_1850[13]), .A1(n17132), .B1(amdemod_d_11__N_2296), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14828), .COUT(n14829));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1199_add_4_10.INIT0 = 16'h656a;
    defparam _add_1_1199_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1199_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1199_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1199_add_4_8 (.A0(amdemod_d_11__N_2305), .B0(amdemod_d_11__N_1861[13]), 
          .C0(n17130), .D0(amdemod_d_11__N_1860[13]), .A1(n17130), .B1(amdemod_d_11__N_2302), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14827), .COUT(n14828));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1199_add_4_8.INIT0 = 16'h656a;
    defparam _add_1_1199_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1199_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1199_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1199_add_4_6 (.A0(amdemod_d_11__N_2311), .B0(amdemod_d_11__N_1871[13]), 
          .C0(n17128), .D0(amdemod_d_11__N_1870[13]), .A1(n17128), .B1(amdemod_d_11__N_2308), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14826), .COUT(n14827));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1199_add_4_6.INIT0 = 16'h656a;
    defparam _add_1_1199_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1199_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1199_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1199_add_4_4 (.A0(amdemod_d_11__N_1874), .B0(square_sum[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1874), .B1(amdemod_d_11__N_2314), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14825), .COUT(n14826));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1199_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1199_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1199_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1199_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1199_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14825));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1199_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1199_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1199_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1199_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_38 (.A0(integrator3_adj_6022[71]), .B0(integrator2_adj_6021[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14819), .S0(n78_adj_5188));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1130_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_36 (.A0(integrator3_adj_6022[69]), .B0(integrator2_adj_6021[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[70]), .B1(integrator2_adj_6021[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14818), .COUT(n14819), .S0(n84_adj_5190), 
          .S1(n81_adj_5189));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_34 (.A0(integrator3_adj_6022[67]), .B0(integrator2_adj_6021[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[68]), .B1(integrator2_adj_6021[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14817), .COUT(n14818), .S0(n90_adj_5192), 
          .S1(n87_adj_5191));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_32 (.A0(integrator3_adj_6022[65]), .B0(integrator2_adj_6021[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[66]), .B1(integrator2_adj_6021[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14816), .COUT(n14817), .S0(n96_adj_5194), 
          .S1(n93_adj_5193));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_30 (.A0(integrator3_adj_6022[63]), .B0(integrator2_adj_6021[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[64]), .B1(integrator2_adj_6021[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14815), .COUT(n14816), .S0(n102_adj_5196), 
          .S1(n99_adj_5195));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_28 (.A0(integrator3_adj_6022[61]), .B0(integrator2_adj_6021[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[62]), .B1(integrator2_adj_6021[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14814), .COUT(n14815), .S0(n108_adj_5198), 
          .S1(n105_adj_5197));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_26 (.A0(integrator3_adj_6022[59]), .B0(integrator2_adj_6021[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[60]), .B1(integrator2_adj_6021[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14813), .COUT(n14814), .S0(n114_adj_5200), 
          .S1(n111_adj_5199));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_24 (.A0(integrator3_adj_6022[57]), .B0(integrator2_adj_6021[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[58]), .B1(integrator2_adj_6021[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14812), .COUT(n14813), .S0(n120_adj_5202), 
          .S1(n117_adj_5201));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_22 (.A0(integrator3_adj_6022[55]), .B0(integrator2_adj_6021[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[56]), .B1(integrator2_adj_6021[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14811), .COUT(n14812), .S0(n126_adj_5204), 
          .S1(n123_adj_5203));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_20 (.A0(integrator3_adj_6022[53]), .B0(integrator2_adj_6021[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[54]), .B1(integrator2_adj_6021[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14810), .COUT(n14811), .S0(n132_adj_5206), 
          .S1(n129_adj_5205));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_18 (.A0(integrator3_adj_6022[51]), .B0(integrator2_adj_6021[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[52]), .B1(integrator2_adj_6021[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14809), .COUT(n14810), .S0(n138_adj_5208), 
          .S1(n135_adj_5207));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_16 (.A0(integrator3_adj_6022[49]), .B0(integrator2_adj_6021[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[50]), .B1(integrator2_adj_6021[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14808), .COUT(n14809), .S0(n144_adj_5210), 
          .S1(n141_adj_5209));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_14 (.A0(integrator3_adj_6022[47]), .B0(integrator2_adj_6021[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[48]), .B1(integrator2_adj_6021[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14807), .COUT(n14808), .S0(n150_adj_5212), 
          .S1(n147_adj_5211));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_12 (.A0(integrator3_adj_6022[45]), .B0(integrator2_adj_6021[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[46]), .B1(integrator2_adj_6021[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14806), .COUT(n14807), .S0(n156_adj_5214), 
          .S1(n153_adj_5213));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_10 (.A0(integrator3_adj_6022[43]), .B0(integrator2_adj_6021[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[44]), .B1(integrator2_adj_6021[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14805), .COUT(n14806), .S0(n162_adj_5216), 
          .S1(n159_adj_5215));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_8 (.A0(integrator3_adj_6022[41]), .B0(integrator2_adj_6021[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[42]), .B1(integrator2_adj_6021[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14804), .COUT(n14805), .S0(n168_adj_5218), 
          .S1(n165_adj_5217));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_6 (.A0(integrator3_adj_6022[39]), .B0(integrator2_adj_6021[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[40]), .B1(integrator2_adj_6021[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14803), .COUT(n14804), .S0(n174_adj_5220), 
          .S1(n171_adj_5219));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_4 (.A0(integrator3_adj_6022[37]), .B0(integrator2_adj_6021[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3_adj_6022[38]), .B1(integrator2_adj_6021[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14802), .COUT(n14803), .S0(n180_adj_5222), 
          .S1(n177_adj_5221));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1130_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1130_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator3_adj_6022[36]), .B1(integrator2_adj_6021[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14802), .S1(n183_adj_5223));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1130_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1130_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1130_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1130_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1052_add_4_9 (.A0(n17162), .B0(n17279), .C0(GND_net), 
          .D0(VCC_net), .A1(n17162), .B1(n17279), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14800), .S0(n25_adj_5225), .S1(n22_adj_5224));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1052_add_4_9.INIT0 = 16'h7777;
    defparam _add_1_1052_add_4_9.INIT1 = 16'h7777;
    defparam _add_1_1052_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1052_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1052_add_4_7 (.A0(n17157), .B0(n6_adj_4757), .C0(GND_net), 
          .D0(VCC_net), .A1(n17162), .B1(n17279), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14799), .COUT(n14800), .S0(n31_adj_5227), .S1(n28_adj_5226));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1052_add_4_7.INIT0 = 16'h6666;
    defparam _add_1_1052_add_4_7.INIT1 = 16'h6666;
    defparam _add_1_1052_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1052_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1052_add_4_5 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1830[1]), .D0(VCC_net), .A1(n17162), .B1(n4_adj_2948), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14798), .COUT(n14799), .S0(n37_adj_5229), 
          .S1(n34_adj_5228));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1052_add_4_5.INIT0 = 16'h1e1e;
    defparam _add_1_1052_add_4_5.INIT1 = 16'h6666;
    defparam _add_1_1052_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1052_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1052_add_4_3 (.A0(n17137), .B0(square_sum[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[20]), .B1(n17279), .C1(n17162), 
          .D1(n17146), .CIN(n14797), .COUT(n14798), .S0(n43_adj_5231), 
          .S1(n40_adj_5230));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1052_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_1052_add_4_3.INIT1 = 16'h9a95;
    defparam _add_1_1052_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1052_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1052_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[18]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14797), .S1(n46_adj_5232));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1052_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1052_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1052_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1052_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_38 (.A0(comb_d8[71]), .B0(comb8[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14796), .S0(n78_adj_5233));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1157_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_36 (.A0(comb_d8[69]), .B0(comb8[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[70]), .B1(comb8[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14795), .COUT(n14796), .S0(n84_adj_5235), 
          .S1(n81_adj_5234));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_34 (.A0(comb_d8[67]), .B0(comb8[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[68]), .B1(comb8[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14794), .COUT(n14795), .S0(n90_adj_5237), 
          .S1(n87_adj_5236));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_32 (.A0(comb_d8[65]), .B0(comb8[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[66]), .B1(comb8[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14793), .COUT(n14794), .S0(n96_adj_5239), 
          .S1(n93_adj_5238));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_30 (.A0(comb_d8[63]), .B0(comb8[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[64]), .B1(comb8[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14792), .COUT(n14793), .S0(n102_adj_5241), 
          .S1(n99_adj_5240));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_28 (.A0(comb_d8[61]), .B0(comb8[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[62]), .B1(comb8[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14791), .COUT(n14792), .S0(n108_adj_5243), 
          .S1(n105_adj_5242));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_26 (.A0(comb_d8[59]), .B0(comb8[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[60]), .B1(comb8[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14790), .COUT(n14791), .S0(n114_adj_5245), 
          .S1(n111_adj_5244));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_24 (.A0(comb_d8[57]), .B0(comb8[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[58]), .B1(comb8[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14789), .COUT(n14790), .S0(n120_adj_5247), 
          .S1(n117_adj_5246));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_22 (.A0(comb_d8[55]), .B0(comb8[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[56]), .B1(comb8[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14788), .COUT(n14789), .S0(n126_adj_5249), 
          .S1(n123_adj_5248));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_20 (.A0(comb_d8[53]), .B0(comb8[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[54]), .B1(comb8[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14787), .COUT(n14788), .S0(n132_adj_5251), 
          .S1(n129_adj_5250));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_18 (.A0(comb_d8[51]), .B0(comb8[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[52]), .B1(comb8[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14786), .COUT(n14787), .S0(n138_adj_5253), 
          .S1(n135_adj_5252));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_16 (.A0(comb_d8[49]), .B0(comb8[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[50]), .B1(comb8[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14785), .COUT(n14786), .S0(n144_adj_5255), 
          .S1(n141_adj_5254));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_14 (.A0(comb_d8[47]), .B0(comb8[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[48]), .B1(comb8[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14784), .COUT(n14785), .S0(n150_adj_5257), 
          .S1(n147_adj_5256));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_12 (.A0(comb_d8[45]), .B0(comb8[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[46]), .B1(comb8[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14783), .COUT(n14784), .S0(n156_adj_5259), 
          .S1(n153_adj_5258));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_10 (.A0(comb_d8[43]), .B0(comb8[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[44]), .B1(comb8[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14782), .COUT(n14783), .S0(n162_adj_5261), 
          .S1(n159_adj_5260));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_8 (.A0(comb_d8[41]), .B0(comb8[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[42]), .B1(comb8[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14781), .COUT(n14782), .S0(n168_adj_5263), 
          .S1(n165_adj_5262));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_6 (.A0(comb_d8[39]), .B0(comb8[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[40]), .B1(comb8[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14780), .COUT(n14781), .S0(n174_adj_5265), 
          .S1(n171_adj_5264));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_4 (.A0(comb_d8[37]), .B0(comb8[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[38]), .B1(comb8[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14779), .COUT(n14780), .S0(n180_adj_5267), 
          .S1(n177_adj_5266));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1157_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1157_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[36]), .B1(comb8[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14779), .S1(n183_adj_5268));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1157_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1157_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1157_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1157_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_38 (.A0(comb_d7[71]), .B0(comb7[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14778), .S0(n78_adj_5269));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1160_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_36 (.A0(comb_d7[69]), .B0(comb7[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[70]), .B1(comb7[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14777), .COUT(n14778), .S0(n84_adj_5271), 
          .S1(n81_adj_5270));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_34 (.A0(comb_d7[67]), .B0(comb7[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[68]), .B1(comb7[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14776), .COUT(n14777), .S0(n90_adj_5273), 
          .S1(n87_adj_5272));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_32 (.A0(comb_d7[65]), .B0(comb7[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[66]), .B1(comb7[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14775), .COUT(n14776), .S0(n96_adj_5275), 
          .S1(n93_adj_5274));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_30 (.A0(comb_d7[63]), .B0(comb7[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[64]), .B1(comb7[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14774), .COUT(n14775), .S0(n102_adj_5277), 
          .S1(n99_adj_5276));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_28 (.A0(comb_d7[61]), .B0(comb7[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[62]), .B1(comb7[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14773), .COUT(n14774), .S0(n108_adj_5279), 
          .S1(n105_adj_5278));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_26 (.A0(comb_d7[59]), .B0(comb7[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[60]), .B1(comb7[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14772), .COUT(n14773), .S0(n114_adj_5281), 
          .S1(n111_adj_5280));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_24 (.A0(comb_d7[57]), .B0(comb7[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[58]), .B1(comb7[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14771), .COUT(n14772), .S0(n120_adj_5283), 
          .S1(n117_adj_5282));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_22 (.A0(comb_d7[55]), .B0(comb7[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[56]), .B1(comb7[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14770), .COUT(n14771), .S0(n126_adj_5285), 
          .S1(n123_adj_5284));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_22.INJECT1_1 = "NO";
    LUT4 i2400_2_lut (.A(led_c_4), .B(n1827), .Z(n2545)) /* synthesis lut_function=(!(A+!(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i2400_2_lut.init = 16'h4444;
    LUT4 i1890_4_lut (.A(n130_adj_5904), .B(n124), .C(led_c_3), .D(n17144), 
         .Z(n11624)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1890_4_lut.init = 16'hcac0;
    LUT4 i273_2_lut_rep_339_3_lut_3_lut (.A(led_c_3), .B(n16220), .C(led_c_4), 
         .Z(n17136)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i273_2_lut_rep_339_3_lut_3_lut.init = 16'h4040;
    CCU2C _add_1_1160_add_4_20 (.A0(comb_d7[53]), .B0(comb7[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[54]), .B1(comb7[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14769), .COUT(n14770), .S0(n132_adj_5287), 
          .S1(n129_adj_5286));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_18 (.A0(comb_d7[51]), .B0(comb7[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[52]), .B1(comb7[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14768), .COUT(n14769), .S0(n138_adj_5289), 
          .S1(n135_adj_5288));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_16 (.A0(comb_d7[49]), .B0(comb7[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[50]), .B1(comb7[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14767), .COUT(n14768), .S0(n144_adj_5291), 
          .S1(n141_adj_5290));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_14 (.A0(comb_d7[47]), .B0(comb7[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[48]), .B1(comb7[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14766), .COUT(n14767), .S0(n150_adj_5293), 
          .S1(n147_adj_5292));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_12 (.A0(comb_d7[45]), .B0(comb7[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[46]), .B1(comb7[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14765), .COUT(n14766), .S0(n156_adj_5295), 
          .S1(n153_adj_5294));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_10 (.A0(comb_d7[43]), .B0(comb7[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[44]), .B1(comb7[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14764), .COUT(n14765), .S0(n162_adj_5297), 
          .S1(n159_adj_5296));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_8 (.A0(comb_d7[41]), .B0(comb7[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[42]), .B1(comb7[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14763), .COUT(n14764), .S0(n168_adj_5299), 
          .S1(n165_adj_5298));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_6 (.A0(comb_d7[39]), .B0(comb7[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[40]), .B1(comb7[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14762), .COUT(n14763), .S0(n174_adj_5301), 
          .S1(n171_adj_5300));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_4 (.A0(comb_d7[37]), .B0(comb7[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[38]), .B1(comb7[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14761), .COUT(n14762), .S0(n180_adj_5303), 
          .S1(n177_adj_5302));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1160_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1160_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[36]), .B1(comb7[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14761), .S1(n183_adj_5304));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1160_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1160_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1160_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1160_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_38 (.A0(comb_d8[35]), .B0(comb8[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14760), .S0(comb9_71__N_1667[35]), .S1(cout_adj_5305));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1163_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_36 (.A0(comb_d8[33]), .B0(comb8[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[34]), .B1(comb8[34]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14759), .COUT(n14760), .S0(comb9_71__N_1667[33]), 
          .S1(comb9_71__N_1667[34]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_34 (.A0(comb_d8[31]), .B0(comb8[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[32]), .B1(comb8[32]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14758), .COUT(n14759), .S0(comb9_71__N_1667[31]), 
          .S1(comb9_71__N_1667[32]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_32 (.A0(comb_d8[29]), .B0(comb8[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[30]), .B1(comb8[30]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14757), .COUT(n14758), .S0(comb9_71__N_1667[29]), 
          .S1(comb9_71__N_1667[30]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_30 (.A0(comb_d8[27]), .B0(comb8[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[28]), .B1(comb8[28]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14756), .COUT(n14757), .S0(comb9_71__N_1667[27]), 
          .S1(comb9_71__N_1667[28]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_28 (.A0(comb_d8[25]), .B0(comb8[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[26]), .B1(comb8[26]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14755), .COUT(n14756), .S0(comb9_71__N_1667[25]), 
          .S1(comb9_71__N_1667[26]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_26 (.A0(comb_d8[23]), .B0(comb8[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[24]), .B1(comb8[24]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14754), .COUT(n14755), .S0(comb9_71__N_1667[23]), 
          .S1(comb9_71__N_1667[24]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_24 (.A0(comb_d8[21]), .B0(comb8[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[22]), .B1(comb8[22]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14753), .COUT(n14754), .S0(comb9_71__N_1667[21]), 
          .S1(comb9_71__N_1667[22]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_22 (.A0(comb_d8[19]), .B0(comb8[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[20]), .B1(comb8[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14752), .COUT(n14753), .S0(comb9_71__N_1667[19]), 
          .S1(comb9_71__N_1667[20]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_20 (.A0(comb_d8[17]), .B0(comb8[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[18]), .B1(comb8[18]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14751), .COUT(n14752), .S0(comb9_71__N_1667[17]), 
          .S1(comb9_71__N_1667[18]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_18 (.A0(comb_d8[15]), .B0(comb8[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[16]), .B1(comb8[16]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14750), .COUT(n14751), .S0(comb9_71__N_1667[15]), 
          .S1(comb9_71__N_1667[16]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_16 (.A0(comb_d8[13]), .B0(comb8[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[14]), .B1(comb8[14]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14749), .COUT(n14750), .S0(comb9_71__N_1667[13]), 
          .S1(comb9_71__N_1667[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_14 (.A0(comb_d8[11]), .B0(comb8[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[12]), .B1(comb8[12]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14748), .COUT(n14749), .S0(comb9_71__N_1667[11]), 
          .S1(comb9_71__N_1667[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_12 (.A0(comb_d8[9]), .B0(comb8[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[10]), .B1(comb8[10]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14747), .COUT(n14748), .S0(comb9_71__N_1667[9]), 
          .S1(comb9_71__N_1667[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_10 (.A0(comb_d8[7]), .B0(comb8[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[8]), .B1(comb8[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14746), .COUT(n14747), .S0(comb9_71__N_1667[7]), 
          .S1(comb9_71__N_1667[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_8 (.A0(comb_d8[5]), .B0(comb8[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[6]), .B1(comb8[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14745), .COUT(n14746), .S0(comb9_71__N_1667[5]), 
          .S1(comb9_71__N_1667[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_6 (.A0(comb_d8[3]), .B0(comb8[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[4]), .B1(comb8[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14744), .COUT(n14745), .S0(comb9_71__N_1667[3]), 
          .S1(comb9_71__N_1667[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_4 (.A0(comb_d8[1]), .B0(comb8[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[2]), .B1(comb8[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14743), .COUT(n14744), .S0(comb9_71__N_1667[1]), 
          .S1(comb9_71__N_1667[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1163_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1163_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8[0]), .B1(comb8[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14743), .S1(comb9_71__N_1667[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1163_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1163_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1163_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1163_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_38 (.A0(comb_d9[35]), .B0(comb9[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14742), .S1(cout_adj_5306));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1166_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_36 (.A0(comb_d9[33]), .B0(comb9[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[34]), .B1(comb9[34]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14741), .COUT(n14742));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_34 (.A0(comb_d9[31]), .B0(comb9[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[32]), .B1(comb9[32]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14740), .COUT(n14741));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_32 (.A0(comb_d9[29]), .B0(comb9[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[30]), .B1(comb9[30]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14739), .COUT(n14740));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_30 (.A0(comb_d9[27]), .B0(comb9[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[28]), .B1(comb9[28]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14738), .COUT(n14739));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_28 (.A0(comb_d9[25]), .B0(comb9[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[26]), .B1(comb9[26]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14737), .COUT(n14738));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_26 (.A0(comb_d9[23]), .B0(comb9[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[24]), .B1(comb9[24]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14736), .COUT(n14737));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_24 (.A0(comb_d9[21]), .B0(comb9[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[22]), .B1(comb9[22]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14735), .COUT(n14736));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_22 (.A0(comb_d9[19]), .B0(comb9[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[20]), .B1(comb9[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14734), .COUT(n14735));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_20 (.A0(comb_d9[17]), .B0(comb9[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[18]), .B1(comb9[18]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14733), .COUT(n14734));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_18 (.A0(comb_d9[15]), .B0(comb9[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[16]), .B1(comb9[16]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14732), .COUT(n14733));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_16 (.A0(comb_d9[13]), .B0(comb9[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[14]), .B1(comb9[14]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14731), .COUT(n14732));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_14 (.A0(comb_d9[11]), .B0(comb9[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[12]), .B1(comb9[12]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14730), .COUT(n14731));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_12 (.A0(comb_d9[9]), .B0(comb9[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[10]), .B1(comb9[10]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14729), .COUT(n14730));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_10 (.A0(comb_d9[7]), .B0(comb9[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[8]), .B1(comb9[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14728), .COUT(n14729));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_8 (.A0(comb_d9[5]), .B0(comb9[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[6]), .B1(comb9[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14727), .COUT(n14728));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_6 (.A0(comb_d9[3]), .B0(comb9[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[4]), .B1(comb9[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14726), .COUT(n14727));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_4 (.A0(comb_d9[1]), .B0(comb9[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[2]), .B1(comb9[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14725), .COUT(n14726));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1166_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1166_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9[0]), .B1(comb9[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14725));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1166_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1166_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1166_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1166_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1202_add_4_10 (.A0(n17162), .B0(n17146), .C0(GND_net), 
          .D0(VCC_net), .A1(n17162), .B1(n17146), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14723), .S0(n27_adj_5349), .S1(n24_adj_5348));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1202_add_4_10.INIT0 = 16'heee1;
    defparam _add_1_1202_add_4_10.INIT1 = 16'heee1;
    defparam _add_1_1202_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1202_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1202_add_4_8 (.A0(n17157), .B0(n17163), .C0(GND_net), 
          .D0(VCC_net), .A1(n17162), .B1(n17146), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14722), .COUT(n14723), .S0(n33_adj_5351), .S1(n30_adj_5350));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1202_add_4_8.INIT0 = 16'h6669;
    defparam _add_1_1202_add_4_8.INIT1 = 16'h6669;
    defparam _add_1_1202_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1202_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1202_add_4_6 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1830[1]), .D0(VCC_net), .A1(n11179), .B1(n4_adj_4982), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14721), .COUT(n14722), .S0(n39), 
          .S1(n36_adj_5352));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1202_add_4_6.INIT0 = 16'h1e11;
    defparam _add_1_1202_add_4_6.INIT1 = 16'h9996;
    defparam _add_1_1202_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1202_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1202_add_4_4 (.A0(square_sum[19]), .B0(n17162), .C0(n17279), 
          .D0(n17146), .A1(n17137), .B1(square_sum[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14720), .COUT(n14721), .S0(n45), .S1(n42));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1202_add_4_4.INIT0 = 16'h596a;
    defparam _add_1_1202_add_4_4.INIT1 = 16'h6665;
    defparam _add_1_1202_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1202_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1202_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[18]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14720), .S1(n48));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1202_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1202_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1202_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1202_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_38 (.A0(integrator_d_tmp_adj_6019[35]), .B0(integrator_tmp_adj_6018[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14719), .S0(comb6_71__N_1451_adj_6052[35]), 
          .S1(cout_adj_5307));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1169_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_36 (.A0(integrator_d_tmp_adj_6019[33]), .B0(integrator_tmp_adj_6018[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[34]), 
          .B1(integrator_tmp_adj_6018[34]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14718), .COUT(n14719), .S0(comb6_71__N_1451_adj_6052[33]), 
          .S1(comb6_71__N_1451_adj_6052[34]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_34 (.A0(integrator_d_tmp_adj_6019[31]), .B0(integrator_tmp_adj_6018[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[32]), 
          .B1(integrator_tmp_adj_6018[32]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14717), .COUT(n14718), .S0(comb6_71__N_1451_adj_6052[31]), 
          .S1(comb6_71__N_1451_adj_6052[32]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_32 (.A0(integrator_d_tmp_adj_6019[29]), .B0(integrator_tmp_adj_6018[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[30]), 
          .B1(integrator_tmp_adj_6018[30]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14716), .COUT(n14717), .S0(comb6_71__N_1451_adj_6052[29]), 
          .S1(comb6_71__N_1451_adj_6052[30]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_30 (.A0(integrator_d_tmp_adj_6019[27]), .B0(integrator_tmp_adj_6018[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[28]), 
          .B1(integrator_tmp_adj_6018[28]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14715), .COUT(n14716), .S0(comb6_71__N_1451_adj_6052[27]), 
          .S1(comb6_71__N_1451_adj_6052[28]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_28 (.A0(integrator_d_tmp_adj_6019[25]), .B0(integrator_tmp_adj_6018[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[26]), 
          .B1(integrator_tmp_adj_6018[26]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14714), .COUT(n14715), .S0(comb6_71__N_1451_adj_6052[25]), 
          .S1(comb6_71__N_1451_adj_6052[26]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_26 (.A0(integrator_d_tmp_adj_6019[23]), .B0(integrator_tmp_adj_6018[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[24]), 
          .B1(integrator_tmp_adj_6018[24]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14713), .COUT(n14714), .S0(comb6_71__N_1451_adj_6052[23]), 
          .S1(comb6_71__N_1451_adj_6052[24]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_24 (.A0(integrator_d_tmp_adj_6019[21]), .B0(integrator_tmp_adj_6018[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[22]), 
          .B1(integrator_tmp_adj_6018[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14712), .COUT(n14713), .S0(comb6_71__N_1451_adj_6052[21]), 
          .S1(comb6_71__N_1451_adj_6052[22]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_22 (.A0(integrator_d_tmp_adj_6019[19]), .B0(integrator_tmp_adj_6018[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[20]), 
          .B1(integrator_tmp_adj_6018[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14711), .COUT(n14712), .S0(comb6_71__N_1451_adj_6052[19]), 
          .S1(comb6_71__N_1451_adj_6052[20]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_20 (.A0(integrator_d_tmp_adj_6019[17]), .B0(integrator_tmp_adj_6018[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[18]), 
          .B1(integrator_tmp_adj_6018[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14710), .COUT(n14711), .S0(comb6_71__N_1451_adj_6052[17]), 
          .S1(comb6_71__N_1451_adj_6052[18]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_18 (.A0(integrator_d_tmp_adj_6019[15]), .B0(integrator_tmp_adj_6018[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[16]), 
          .B1(integrator_tmp_adj_6018[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14709), .COUT(n14710), .S0(comb6_71__N_1451_adj_6052[15]), 
          .S1(comb6_71__N_1451_adj_6052[16]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_16 (.A0(integrator_d_tmp_adj_6019[13]), .B0(integrator_tmp_adj_6018[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[14]), 
          .B1(integrator_tmp_adj_6018[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14708), .COUT(n14709), .S0(comb6_71__N_1451_adj_6052[13]), 
          .S1(comb6_71__N_1451_adj_6052[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_14 (.A0(integrator_d_tmp_adj_6019[11]), .B0(integrator_tmp_adj_6018[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[12]), 
          .B1(integrator_tmp_adj_6018[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14707), .COUT(n14708), .S0(comb6_71__N_1451_adj_6052[11]), 
          .S1(comb6_71__N_1451_adj_6052[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_12 (.A0(integrator_d_tmp_adj_6019[9]), .B0(integrator_tmp_adj_6018[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[10]), 
          .B1(integrator_tmp_adj_6018[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14706), .COUT(n14707), .S0(comb6_71__N_1451_adj_6052[9]), 
          .S1(comb6_71__N_1451_adj_6052[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_10 (.A0(integrator_d_tmp_adj_6019[7]), .B0(integrator_tmp_adj_6018[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[8]), 
          .B1(integrator_tmp_adj_6018[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14705), .COUT(n14706), .S0(comb6_71__N_1451_adj_6052[7]), 
          .S1(comb6_71__N_1451_adj_6052[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_8 (.A0(integrator_d_tmp_adj_6019[5]), .B0(integrator_tmp_adj_6018[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[6]), 
          .B1(integrator_tmp_adj_6018[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14704), .COUT(n14705), .S0(comb6_71__N_1451_adj_6052[5]), 
          .S1(comb6_71__N_1451_adj_6052[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_6 (.A0(integrator_d_tmp_adj_6019[3]), .B0(integrator_tmp_adj_6018[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[4]), 
          .B1(integrator_tmp_adj_6018[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14703), .COUT(n14704), .S0(comb6_71__N_1451_adj_6052[3]), 
          .S1(comb6_71__N_1451_adj_6052[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_4 (.A0(integrator_d_tmp_adj_6019[1]), .B0(integrator_tmp_adj_6018[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[2]), 
          .B1(integrator_tmp_adj_6018[2]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14702), .COUT(n14703), .S0(comb6_71__N_1451_adj_6052[1]), 
          .S1(comb6_71__N_1451_adj_6052[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1169_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1169_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[0]), .B1(integrator_tmp_adj_6018[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14702), .S1(comb6_71__N_1451_adj_6052[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1169_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1169_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1169_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1169_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_38 (.A0(comb_d6_adj_6026[35]), .B0(comb6_adj_6025[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14701), .S0(comb7_71__N_1523_adj_6053[35]), 
          .S1(cout_adj_5308));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1172_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_36 (.A0(comb_d6_adj_6026[33]), .B0(comb6_adj_6025[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[34]), .B1(comb6_adj_6025[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14700), .COUT(n14701), .S0(comb7_71__N_1523_adj_6053[33]), 
          .S1(comb7_71__N_1523_adj_6053[34]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_34 (.A0(comb_d6_adj_6026[31]), .B0(comb6_adj_6025[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[32]), .B1(comb6_adj_6025[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14699), .COUT(n14700), .S0(comb7_71__N_1523_adj_6053[31]), 
          .S1(comb7_71__N_1523_adj_6053[32]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_32 (.A0(comb_d6_adj_6026[29]), .B0(comb6_adj_6025[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[30]), .B1(comb6_adj_6025[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14698), .COUT(n14699), .S0(comb7_71__N_1523_adj_6053[29]), 
          .S1(comb7_71__N_1523_adj_6053[30]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_30 (.A0(comb_d6_adj_6026[27]), .B0(comb6_adj_6025[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[28]), .B1(comb6_adj_6025[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14697), .COUT(n14698), .S0(comb7_71__N_1523_adj_6053[27]), 
          .S1(comb7_71__N_1523_adj_6053[28]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_28 (.A0(comb_d6_adj_6026[25]), .B0(comb6_adj_6025[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[26]), .B1(comb6_adj_6025[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14696), .COUT(n14697), .S0(comb7_71__N_1523_adj_6053[25]), 
          .S1(comb7_71__N_1523_adj_6053[26]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_26 (.A0(comb_d6_adj_6026[23]), .B0(comb6_adj_6025[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[24]), .B1(comb6_adj_6025[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14695), .COUT(n14696), .S0(comb7_71__N_1523_adj_6053[23]), 
          .S1(comb7_71__N_1523_adj_6053[24]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_24 (.A0(comb_d6_adj_6026[21]), .B0(comb6_adj_6025[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[22]), .B1(comb6_adj_6025[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14694), .COUT(n14695), .S0(comb7_71__N_1523_adj_6053[21]), 
          .S1(comb7_71__N_1523_adj_6053[22]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_22 (.A0(comb_d6_adj_6026[19]), .B0(comb6_adj_6025[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[20]), .B1(comb6_adj_6025[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14693), .COUT(n14694), .S0(comb7_71__N_1523_adj_6053[19]), 
          .S1(comb7_71__N_1523_adj_6053[20]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_20 (.A0(comb_d6_adj_6026[17]), .B0(comb6_adj_6025[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[18]), .B1(comb6_adj_6025[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14692), .COUT(n14693), .S0(comb7_71__N_1523_adj_6053[17]), 
          .S1(comb7_71__N_1523_adj_6053[18]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_18 (.A0(comb_d6_adj_6026[15]), .B0(comb6_adj_6025[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[16]), .B1(comb6_adj_6025[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14691), .COUT(n14692), .S0(comb7_71__N_1523_adj_6053[15]), 
          .S1(comb7_71__N_1523_adj_6053[16]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_16 (.A0(comb_d6_adj_6026[13]), .B0(comb6_adj_6025[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[14]), .B1(comb6_adj_6025[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14690), .COUT(n14691), .S0(comb7_71__N_1523_adj_6053[13]), 
          .S1(comb7_71__N_1523_adj_6053[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_14 (.A0(comb_d6_adj_6026[11]), .B0(comb6_adj_6025[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[12]), .B1(comb6_adj_6025[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14689), .COUT(n14690), .S0(comb7_71__N_1523_adj_6053[11]), 
          .S1(comb7_71__N_1523_adj_6053[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_12 (.A0(comb_d6_adj_6026[9]), .B0(comb6_adj_6025[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[10]), .B1(comb6_adj_6025[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14688), .COUT(n14689), .S0(comb7_71__N_1523_adj_6053[9]), 
          .S1(comb7_71__N_1523_adj_6053[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_10 (.A0(comb_d6_adj_6026[7]), .B0(comb6_adj_6025[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[8]), .B1(comb6_adj_6025[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14687), .COUT(n14688), .S0(comb7_71__N_1523_adj_6053[7]), 
          .S1(comb7_71__N_1523_adj_6053[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_8 (.A0(comb_d6_adj_6026[5]), .B0(comb6_adj_6025[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[6]), .B1(comb6_adj_6025[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14686), .COUT(n14687), .S0(comb7_71__N_1523_adj_6053[5]), 
          .S1(comb7_71__N_1523_adj_6053[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_6 (.A0(comb_d6_adj_6026[3]), .B0(comb6_adj_6025[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[4]), .B1(comb6_adj_6025[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14685), .COUT(n14686), .S0(comb7_71__N_1523_adj_6053[3]), 
          .S1(comb7_71__N_1523_adj_6053[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_4 (.A0(comb_d6_adj_6026[1]), .B0(comb6_adj_6025[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[2]), .B1(comb6_adj_6025[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14684), .COUT(n14685), .S0(comb7_71__N_1523_adj_6053[1]), 
          .S1(comb7_71__N_1523_adj_6053[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1172_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1172_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6_adj_6026[0]), .B1(comb6_adj_6025[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14684), .S1(comb7_71__N_1523_adj_6053[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1172_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1172_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1172_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1172_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_37 (.A0(integrator2_adj_6021[70]), .B0(cout_adj_5164), 
          .C0(n81_adj_5189), .D0(integrator3_adj_6022[70]), .A1(integrator2_adj_6021[71]), 
          .B1(cout_adj_5164), .C1(n78_adj_5188), .D1(integrator3_adj_6022[71]), 
          .CIN(n14682), .S0(integrator3_71__N_562_adj_6038[70]), .S1(integrator3_71__N_562_adj_6038[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_35 (.A0(integrator2_adj_6021[68]), .B0(cout_adj_5164), 
          .C0(n87_adj_5191), .D0(integrator3_adj_6022[68]), .A1(integrator2_adj_6021[69]), 
          .B1(cout_adj_5164), .C1(n84_adj_5190), .D1(integrator3_adj_6022[69]), 
          .CIN(n14681), .COUT(n14682), .S0(integrator3_71__N_562_adj_6038[68]), 
          .S1(integrator3_71__N_562_adj_6038[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_33 (.A0(integrator2_adj_6021[66]), .B0(cout_adj_5164), 
          .C0(n93_adj_5193), .D0(integrator3_adj_6022[66]), .A1(integrator2_adj_6021[67]), 
          .B1(cout_adj_5164), .C1(n90_adj_5192), .D1(integrator3_adj_6022[67]), 
          .CIN(n14680), .COUT(n14681), .S0(integrator3_71__N_562_adj_6038[66]), 
          .S1(integrator3_71__N_562_adj_6038[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_31 (.A0(integrator2_adj_6021[64]), .B0(cout_adj_5164), 
          .C0(n99_adj_5195), .D0(integrator3_adj_6022[64]), .A1(integrator2_adj_6021[65]), 
          .B1(cout_adj_5164), .C1(n96_adj_5194), .D1(integrator3_adj_6022[65]), 
          .CIN(n14679), .COUT(n14680), .S0(integrator3_71__N_562_adj_6038[64]), 
          .S1(integrator3_71__N_562_adj_6038[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_29 (.A0(integrator2_adj_6021[62]), .B0(cout_adj_5164), 
          .C0(n105_adj_5197), .D0(integrator3_adj_6022[62]), .A1(integrator2_adj_6021[63]), 
          .B1(cout_adj_5164), .C1(n102_adj_5196), .D1(integrator3_adj_6022[63]), 
          .CIN(n14678), .COUT(n14679), .S0(integrator3_71__N_562_adj_6038[62]), 
          .S1(integrator3_71__N_562_adj_6038[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_27 (.A0(integrator2_adj_6021[60]), .B0(cout_adj_5164), 
          .C0(n111_adj_5199), .D0(integrator3_adj_6022[60]), .A1(integrator2_adj_6021[61]), 
          .B1(cout_adj_5164), .C1(n108_adj_5198), .D1(integrator3_adj_6022[61]), 
          .CIN(n14677), .COUT(n14678), .S0(integrator3_71__N_562_adj_6038[60]), 
          .S1(integrator3_71__N_562_adj_6038[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_25 (.A0(integrator2_adj_6021[58]), .B0(cout_adj_5164), 
          .C0(n117_adj_5201), .D0(integrator3_adj_6022[58]), .A1(integrator2_adj_6021[59]), 
          .B1(cout_adj_5164), .C1(n114_adj_5200), .D1(integrator3_adj_6022[59]), 
          .CIN(n14676), .COUT(n14677), .S0(integrator3_71__N_562_adj_6038[58]), 
          .S1(integrator3_71__N_562_adj_6038[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_23 (.A0(integrator2_adj_6021[56]), .B0(cout_adj_5164), 
          .C0(n123_adj_5203), .D0(integrator3_adj_6022[56]), .A1(integrator2_adj_6021[57]), 
          .B1(cout_adj_5164), .C1(n120_adj_5202), .D1(integrator3_adj_6022[57]), 
          .CIN(n14675), .COUT(n14676), .S0(integrator3_71__N_562_adj_6038[56]), 
          .S1(integrator3_71__N_562_adj_6038[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_21 (.A0(integrator2_adj_6021[54]), .B0(cout_adj_5164), 
          .C0(n129_adj_5205), .D0(integrator3_adj_6022[54]), .A1(integrator2_adj_6021[55]), 
          .B1(cout_adj_5164), .C1(n126_adj_5204), .D1(integrator3_adj_6022[55]), 
          .CIN(n14674), .COUT(n14675), .S0(integrator3_71__N_562_adj_6038[54]), 
          .S1(integrator3_71__N_562_adj_6038[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_19 (.A0(integrator2_adj_6021[52]), .B0(cout_adj_5164), 
          .C0(n135_adj_5207), .D0(integrator3_adj_6022[52]), .A1(integrator2_adj_6021[53]), 
          .B1(cout_adj_5164), .C1(n132_adj_5206), .D1(integrator3_adj_6022[53]), 
          .CIN(n14673), .COUT(n14674), .S0(integrator3_71__N_562_adj_6038[52]), 
          .S1(integrator3_71__N_562_adj_6038[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_17 (.A0(integrator2_adj_6021[50]), .B0(cout_adj_5164), 
          .C0(n141_adj_5209), .D0(integrator3_adj_6022[50]), .A1(integrator2_adj_6021[51]), 
          .B1(cout_adj_5164), .C1(n138_adj_5208), .D1(integrator3_adj_6022[51]), 
          .CIN(n14672), .COUT(n14673), .S0(integrator3_71__N_562_adj_6038[50]), 
          .S1(integrator3_71__N_562_adj_6038[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_15 (.A0(integrator2_adj_6021[48]), .B0(cout_adj_5164), 
          .C0(n147_adj_5211), .D0(integrator3_adj_6022[48]), .A1(integrator2_adj_6021[49]), 
          .B1(cout_adj_5164), .C1(n144_adj_5210), .D1(integrator3_adj_6022[49]), 
          .CIN(n14671), .COUT(n14672), .S0(integrator3_71__N_562_adj_6038[48]), 
          .S1(integrator3_71__N_562_adj_6038[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_13 (.A0(integrator2_adj_6021[46]), .B0(cout_adj_5164), 
          .C0(n153_adj_5213), .D0(integrator3_adj_6022[46]), .A1(integrator2_adj_6021[47]), 
          .B1(cout_adj_5164), .C1(n150_adj_5212), .D1(integrator3_adj_6022[47]), 
          .CIN(n14670), .COUT(n14671), .S0(integrator3_71__N_562_adj_6038[46]), 
          .S1(integrator3_71__N_562_adj_6038[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_11 (.A0(integrator2_adj_6021[44]), .B0(cout_adj_5164), 
          .C0(n159_adj_5215), .D0(integrator3_adj_6022[44]), .A1(integrator2_adj_6021[45]), 
          .B1(cout_adj_5164), .C1(n156_adj_5214), .D1(integrator3_adj_6022[45]), 
          .CIN(n14669), .COUT(n14670), .S0(integrator3_71__N_562_adj_6038[44]), 
          .S1(integrator3_71__N_562_adj_6038[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_9 (.A0(integrator2_adj_6021[42]), .B0(cout_adj_5164), 
          .C0(n165_adj_5217), .D0(integrator3_adj_6022[42]), .A1(integrator2_adj_6021[43]), 
          .B1(cout_adj_5164), .C1(n162_adj_5216), .D1(integrator3_adj_6022[43]), 
          .CIN(n14668), .COUT(n14669), .S0(integrator3_71__N_562_adj_6038[42]), 
          .S1(integrator3_71__N_562_adj_6038[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_7 (.A0(integrator2_adj_6021[40]), .B0(cout_adj_5164), 
          .C0(n171_adj_5219), .D0(integrator3_adj_6022[40]), .A1(integrator2_adj_6021[41]), 
          .B1(cout_adj_5164), .C1(n168_adj_5218), .D1(integrator3_adj_6022[41]), 
          .CIN(n14667), .COUT(n14668), .S0(integrator3_71__N_562_adj_6038[40]), 
          .S1(integrator3_71__N_562_adj_6038[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_5 (.A0(integrator2_adj_6021[38]), .B0(cout_adj_5164), 
          .C0(n177_adj_5221), .D0(integrator3_adj_6022[38]), .A1(integrator2_adj_6021[39]), 
          .B1(cout_adj_5164), .C1(n174_adj_5220), .D1(integrator3_adj_6022[39]), 
          .CIN(n14666), .COUT(n14667), .S0(integrator3_71__N_562_adj_6038[38]), 
          .S1(integrator3_71__N_562_adj_6038[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_3 (.A0(integrator2_adj_6021[36]), .B0(cout_adj_5164), 
          .C0(n183_adj_5223), .D0(integrator3_adj_6022[36]), .A1(integrator2_adj_6021[37]), 
          .B1(cout_adj_5164), .C1(n180_adj_5222), .D1(integrator3_adj_6022[37]), 
          .CIN(n14665), .COUT(n14666), .S0(integrator3_71__N_562_adj_6038[36]), 
          .S1(integrator3_71__N_562_adj_6038[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1100_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1100_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1100_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5164), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14665));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1100_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1100_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1100_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1100_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_37 (.A0(integrator_tmp_adj_6018[70]), .B0(cout_adj_5307), 
          .C0(n81_adj_5800), .D0(n3_adj_4839), .A1(integrator_tmp_adj_6018[71]), 
          .B1(cout_adj_5307), .C1(n78_adj_5799), .D1(n2_adj_4838), .CIN(n14660), 
          .S0(comb6_71__N_1451_adj_6052[70]), .S1(comb6_71__N_1451_adj_6052[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_35 (.A0(integrator_tmp_adj_6018[68]), .B0(cout_adj_5307), 
          .C0(n87_adj_5802), .D0(n5_adj_4841), .A1(integrator_tmp_adj_6018[69]), 
          .B1(cout_adj_5307), .C1(n84_adj_5801), .D1(n4_adj_4840), .CIN(n14659), 
          .COUT(n14660), .S0(comb6_71__N_1451_adj_6052[68]), .S1(comb6_71__N_1451_adj_6052[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_33 (.A0(integrator_tmp_adj_6018[66]), .B0(cout_adj_5307), 
          .C0(n93_adj_5804), .D0(n7_adj_4843), .A1(integrator_tmp_adj_6018[67]), 
          .B1(cout_adj_5307), .C1(n90_adj_5803), .D1(n6_adj_4842), .CIN(n14658), 
          .COUT(n14659), .S0(comb6_71__N_1451_adj_6052[66]), .S1(comb6_71__N_1451_adj_6052[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_31 (.A0(integrator_tmp_adj_6018[64]), .B0(cout_adj_5307), 
          .C0(n99_adj_5806), .D0(n9_adj_4845), .A1(integrator_tmp_adj_6018[65]), 
          .B1(cout_adj_5307), .C1(n96_adj_5805), .D1(n8_adj_4844), .CIN(n14657), 
          .COUT(n14658), .S0(comb6_71__N_1451_adj_6052[64]), .S1(comb6_71__N_1451_adj_6052[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_29 (.A0(integrator_tmp_adj_6018[62]), .B0(cout_adj_5307), 
          .C0(n105_adj_5808), .D0(n11_adj_4847), .A1(integrator_tmp_adj_6018[63]), 
          .B1(cout_adj_5307), .C1(n102_adj_5807), .D1(n10_adj_4846), .CIN(n14656), 
          .COUT(n14657), .S0(comb6_71__N_1451_adj_6052[62]), .S1(comb6_71__N_1451_adj_6052[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_27 (.A0(integrator_tmp_adj_6018[60]), .B0(cout_adj_5307), 
          .C0(n111_adj_5810), .D0(n13_adj_4849), .A1(integrator_tmp_adj_6018[61]), 
          .B1(cout_adj_5307), .C1(n108_adj_5809), .D1(n12_adj_4848), .CIN(n14655), 
          .COUT(n14656), .S0(comb6_71__N_1451_adj_6052[60]), .S1(comb6_71__N_1451_adj_6052[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_25 (.A0(integrator_tmp_adj_6018[58]), .B0(cout_adj_5307), 
          .C0(n117_adj_5812), .D0(n15_adj_4851), .A1(integrator_tmp_adj_6018[59]), 
          .B1(cout_adj_5307), .C1(n114_adj_5811), .D1(n14_adj_4850), .CIN(n14654), 
          .COUT(n14655), .S0(comb6_71__N_1451_adj_6052[58]), .S1(comb6_71__N_1451_adj_6052[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_23 (.A0(integrator_tmp_adj_6018[56]), .B0(cout_adj_5307), 
          .C0(n123_adj_5814), .D0(n17_adj_4853), .A1(integrator_tmp_adj_6018[57]), 
          .B1(cout_adj_5307), .C1(n120_adj_5813), .D1(n16_adj_4852), .CIN(n14653), 
          .COUT(n14654), .S0(comb6_71__N_1451_adj_6052[56]), .S1(comb6_71__N_1451_adj_6052[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_21 (.A0(integrator_tmp_adj_6018[54]), .B0(cout_adj_5307), 
          .C0(n129_adj_5816), .D0(n19_adj_4855), .A1(integrator_tmp_adj_6018[55]), 
          .B1(cout_adj_5307), .C1(n126_adj_5815), .D1(n18_adj_4854), .CIN(n14652), 
          .COUT(n14653), .S0(comb6_71__N_1451_adj_6052[54]), .S1(comb6_71__N_1451_adj_6052[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_19 (.A0(integrator_tmp_adj_6018[52]), .B0(cout_adj_5307), 
          .C0(n135_adj_5818), .D0(n21_adj_4857), .A1(integrator_tmp_adj_6018[53]), 
          .B1(cout_adj_5307), .C1(n132_adj_5817), .D1(n20_adj_4856), .CIN(n14651), 
          .COUT(n14652), .S0(comb6_71__N_1451_adj_6052[52]), .S1(comb6_71__N_1451_adj_6052[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_17 (.A0(integrator_tmp_adj_6018[50]), .B0(cout_adj_5307), 
          .C0(n141_adj_5820), .D0(n23_adj_4859), .A1(integrator_tmp_adj_6018[51]), 
          .B1(cout_adj_5307), .C1(n138_adj_5819), .D1(n22_adj_4858), .CIN(n14650), 
          .COUT(n14651), .S0(comb6_71__N_1451_adj_6052[50]), .S1(comb6_71__N_1451_adj_6052[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_15 (.A0(integrator_tmp_adj_6018[48]), .B0(cout_adj_5307), 
          .C0(n147_adj_5822), .D0(n25_adj_4861), .A1(integrator_tmp_adj_6018[49]), 
          .B1(cout_adj_5307), .C1(n144_adj_5821), .D1(n24_adj_4860), .CIN(n14649), 
          .COUT(n14650), .S0(comb6_71__N_1451_adj_6052[48]), .S1(comb6_71__N_1451_adj_6052[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_13 (.A0(integrator_tmp_adj_6018[46]), .B0(cout_adj_5307), 
          .C0(n153_adj_5824), .D0(n27_adj_4863), .A1(integrator_tmp_adj_6018[47]), 
          .B1(cout_adj_5307), .C1(n150_adj_5823), .D1(n26_adj_4862), .CIN(n14648), 
          .COUT(n14649), .S0(comb6_71__N_1451_adj_6052[46]), .S1(comb6_71__N_1451_adj_6052[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_11 (.A0(integrator_tmp_adj_6018[44]), .B0(cout_adj_5307), 
          .C0(n159_adj_5826), .D0(n29_adj_4865), .A1(integrator_tmp_adj_6018[45]), 
          .B1(cout_adj_5307), .C1(n156_adj_5825), .D1(n28_adj_4864), .CIN(n14647), 
          .COUT(n14648), .S0(comb6_71__N_1451_adj_6052[44]), .S1(comb6_71__N_1451_adj_6052[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_9 (.A0(integrator_tmp_adj_6018[42]), .B0(cout_adj_5307), 
          .C0(n165_adj_5828), .D0(n31_adj_4867), .A1(integrator_tmp_adj_6018[43]), 
          .B1(cout_adj_5307), .C1(n162_adj_5827), .D1(n30_adj_4866), .CIN(n14646), 
          .COUT(n14647), .S0(comb6_71__N_1451_adj_6052[42]), .S1(comb6_71__N_1451_adj_6052[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_7 (.A0(integrator_tmp_adj_6018[40]), .B0(cout_adj_5307), 
          .C0(n171_adj_5830), .D0(n33_adj_4869), .A1(integrator_tmp_adj_6018[41]), 
          .B1(cout_adj_5307), .C1(n168_adj_5829), .D1(n32_adj_4868), .CIN(n14645), 
          .COUT(n14646), .S0(comb6_71__N_1451_adj_6052[40]), .S1(comb6_71__N_1451_adj_6052[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_5 (.A0(integrator_tmp_adj_6018[38]), .B0(cout_adj_5307), 
          .C0(n177_adj_5832), .D0(n35_adj_4871), .A1(integrator_tmp_adj_6018[39]), 
          .B1(cout_adj_5307), .C1(n174_adj_5831), .D1(n34_adj_4870), .CIN(n14644), 
          .COUT(n14645), .S0(comb6_71__N_1451_adj_6052[38]), .S1(comb6_71__N_1451_adj_6052[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_3 (.A0(integrator_tmp_adj_6018[36]), .B0(cout_adj_5307), 
          .C0(n183_adj_5834), .D0(n37_adj_4873), .A1(integrator_tmp_adj_6018[37]), 
          .B1(cout_adj_5307), .C1(n180_adj_5833), .D1(n36_adj_4872), .CIN(n14643), 
          .COUT(n14644), .S0(comb6_71__N_1451_adj_6052[36]), .S1(comb6_71__N_1451_adj_6052[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1079_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1079_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1079_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5307), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14643));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1079_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1079_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1079_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1079_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_37 (.A0(integrator1_adj_6020[70]), .B0(cout_adj_5163), 
          .C0(n81_adj_5024), .D0(integrator2_adj_6021[70]), .A1(integrator1_adj_6020[71]), 
          .B1(cout_adj_5163), .C1(n78_adj_5023), .D1(integrator2_adj_6021[71]), 
          .CIN(n14638), .S0(integrator2_71__N_490_adj_6037[70]), .S1(integrator2_71__N_490_adj_6037[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_35 (.A0(integrator1_adj_6020[68]), .B0(cout_adj_5163), 
          .C0(n87_adj_5026), .D0(integrator2_adj_6021[68]), .A1(integrator1_adj_6020[69]), 
          .B1(cout_adj_5163), .C1(n84_adj_5025), .D1(integrator2_adj_6021[69]), 
          .CIN(n14637), .COUT(n14638), .S0(integrator2_71__N_490_adj_6037[68]), 
          .S1(integrator2_71__N_490_adj_6037[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_33 (.A0(integrator1_adj_6020[66]), .B0(cout_adj_5163), 
          .C0(n93_adj_5028), .D0(integrator2_adj_6021[66]), .A1(integrator1_adj_6020[67]), 
          .B1(cout_adj_5163), .C1(n90_adj_5027), .D1(integrator2_adj_6021[67]), 
          .CIN(n14636), .COUT(n14637), .S0(integrator2_71__N_490_adj_6037[66]), 
          .S1(integrator2_71__N_490_adj_6037[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_31 (.A0(integrator1_adj_6020[64]), .B0(cout_adj_5163), 
          .C0(n99_adj_5030), .D0(integrator2_adj_6021[64]), .A1(integrator1_adj_6020[65]), 
          .B1(cout_adj_5163), .C1(n96_adj_5029), .D1(integrator2_adj_6021[65]), 
          .CIN(n14635), .COUT(n14636), .S0(integrator2_71__N_490_adj_6037[64]), 
          .S1(integrator2_71__N_490_adj_6037[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_29 (.A0(integrator1_adj_6020[62]), .B0(cout_adj_5163), 
          .C0(n105_adj_5032), .D0(integrator2_adj_6021[62]), .A1(integrator1_adj_6020[63]), 
          .B1(cout_adj_5163), .C1(n102_adj_5031), .D1(integrator2_adj_6021[63]), 
          .CIN(n14634), .COUT(n14635), .S0(integrator2_71__N_490_adj_6037[62]), 
          .S1(integrator2_71__N_490_adj_6037[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_27 (.A0(integrator1_adj_6020[60]), .B0(cout_adj_5163), 
          .C0(n111_adj_5034), .D0(integrator2_adj_6021[60]), .A1(integrator1_adj_6020[61]), 
          .B1(cout_adj_5163), .C1(n108_adj_5033), .D1(integrator2_adj_6021[61]), 
          .CIN(n14633), .COUT(n14634), .S0(integrator2_71__N_490_adj_6037[60]), 
          .S1(integrator2_71__N_490_adj_6037[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_27.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n17288), .B(n17153), .C(led_c_0), .D(led_c_1), 
         .Z(n16220)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i1_4_lut.init = 16'h0040;
    LUT4 i1645_3_lut_4_lut (.A(n17288), .B(n17150), .C(led_c_3), .D(n187), 
         .Z(n11367)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1645_3_lut_4_lut.init = 16'hf808;
    CCU2C _add_1_1103_add_4_25 (.A0(integrator1_adj_6020[58]), .B0(cout_adj_5163), 
          .C0(n117_adj_5036), .D0(integrator2_adj_6021[58]), .A1(integrator1_adj_6020[59]), 
          .B1(cout_adj_5163), .C1(n114_adj_5035), .D1(integrator2_adj_6021[59]), 
          .CIN(n14632), .COUT(n14633), .S0(integrator2_71__N_490_adj_6037[58]), 
          .S1(integrator2_71__N_490_adj_6037[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_23 (.A0(integrator1_adj_6020[56]), .B0(cout_adj_5163), 
          .C0(n123_adj_5038), .D0(integrator2_adj_6021[56]), .A1(integrator1_adj_6020[57]), 
          .B1(cout_adj_5163), .C1(n120_adj_5037), .D1(integrator2_adj_6021[57]), 
          .CIN(n14631), .COUT(n14632), .S0(integrator2_71__N_490_adj_6037[56]), 
          .S1(integrator2_71__N_490_adj_6037[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_21 (.A0(integrator1_adj_6020[54]), .B0(cout_adj_5163), 
          .C0(n129_adj_5040), .D0(integrator2_adj_6021[54]), .A1(integrator1_adj_6020[55]), 
          .B1(cout_adj_5163), .C1(n126_adj_5039), .D1(integrator2_adj_6021[55]), 
          .CIN(n14630), .COUT(n14631), .S0(integrator2_71__N_490_adj_6037[54]), 
          .S1(integrator2_71__N_490_adj_6037[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_19 (.A0(integrator1_adj_6020[52]), .B0(cout_adj_5163), 
          .C0(n135_adj_5042), .D0(integrator2_adj_6021[52]), .A1(integrator1_adj_6020[53]), 
          .B1(cout_adj_5163), .C1(n132_adj_5041), .D1(integrator2_adj_6021[53]), 
          .CIN(n14629), .COUT(n14630), .S0(integrator2_71__N_490_adj_6037[52]), 
          .S1(integrator2_71__N_490_adj_6037[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_17 (.A0(integrator1_adj_6020[50]), .B0(cout_adj_5163), 
          .C0(n141_adj_5044), .D0(integrator2_adj_6021[50]), .A1(integrator1_adj_6020[51]), 
          .B1(cout_adj_5163), .C1(n138_adj_5043), .D1(integrator2_adj_6021[51]), 
          .CIN(n14628), .COUT(n14629), .S0(integrator2_71__N_490_adj_6037[50]), 
          .S1(integrator2_71__N_490_adj_6037[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_15 (.A0(integrator1_adj_6020[48]), .B0(cout_adj_5163), 
          .C0(n147_adj_5046), .D0(integrator2_adj_6021[48]), .A1(integrator1_adj_6020[49]), 
          .B1(cout_adj_5163), .C1(n144_adj_5045), .D1(integrator2_adj_6021[49]), 
          .CIN(n14627), .COUT(n14628), .S0(integrator2_71__N_490_adj_6037[48]), 
          .S1(integrator2_71__N_490_adj_6037[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_13 (.A0(integrator1_adj_6020[46]), .B0(cout_adj_5163), 
          .C0(n153_adj_5048), .D0(integrator2_adj_6021[46]), .A1(integrator1_adj_6020[47]), 
          .B1(cout_adj_5163), .C1(n150_adj_5047), .D1(integrator2_adj_6021[47]), 
          .CIN(n14626), .COUT(n14627), .S0(integrator2_71__N_490_adj_6037[46]), 
          .S1(integrator2_71__N_490_adj_6037[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_11 (.A0(integrator1_adj_6020[44]), .B0(cout_adj_5163), 
          .C0(n159_adj_5050), .D0(integrator2_adj_6021[44]), .A1(integrator1_adj_6020[45]), 
          .B1(cout_adj_5163), .C1(n156_adj_5049), .D1(integrator2_adj_6021[45]), 
          .CIN(n14625), .COUT(n14626), .S0(integrator2_71__N_490_adj_6037[44]), 
          .S1(integrator2_71__N_490_adj_6037[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_9 (.A0(integrator1_adj_6020[42]), .B0(cout_adj_5163), 
          .C0(n165_adj_5052), .D0(integrator2_adj_6021[42]), .A1(integrator1_adj_6020[43]), 
          .B1(cout_adj_5163), .C1(n162_adj_5051), .D1(integrator2_adj_6021[43]), 
          .CIN(n14624), .COUT(n14625), .S0(integrator2_71__N_490_adj_6037[42]), 
          .S1(integrator2_71__N_490_adj_6037[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_7 (.A0(integrator1_adj_6020[40]), .B0(cout_adj_5163), 
          .C0(n171_adj_5054), .D0(integrator2_adj_6021[40]), .A1(integrator1_adj_6020[41]), 
          .B1(cout_adj_5163), .C1(n168_adj_5053), .D1(integrator2_adj_6021[41]), 
          .CIN(n14623), .COUT(n14624), .S0(integrator2_71__N_490_adj_6037[40]), 
          .S1(integrator2_71__N_490_adj_6037[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_5 (.A0(integrator1_adj_6020[38]), .B0(cout_adj_5163), 
          .C0(n177_adj_5056), .D0(integrator2_adj_6021[38]), .A1(integrator1_adj_6020[39]), 
          .B1(cout_adj_5163), .C1(n174_adj_5055), .D1(integrator2_adj_6021[39]), 
          .CIN(n14622), .COUT(n14623), .S0(integrator2_71__N_490_adj_6037[38]), 
          .S1(integrator2_71__N_490_adj_6037[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_3 (.A0(integrator1_adj_6020[36]), .B0(cout_adj_5163), 
          .C0(n183_adj_5058), .D0(integrator2_adj_6021[36]), .A1(integrator1_adj_6020[37]), 
          .B1(cout_adj_5163), .C1(n180_adj_5057), .D1(integrator2_adj_6021[37]), 
          .CIN(n14621), .COUT(n14622), .S0(integrator2_71__N_490_adj_6037[36]), 
          .S1(integrator2_71__N_490_adj_6037[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1103_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1103_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1103_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5163), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14621));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1103_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1103_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1103_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1103_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_37 (.A0(comb6_adj_6025[70]), .B0(cout_adj_5308), 
          .C0(n81_adj_5764), .D0(n3_adj_4875), .A1(comb6_adj_6025[71]), 
          .B1(cout_adj_5308), .C1(n78_adj_5763), .D1(n2_adj_4874), .CIN(n14616), 
          .S0(comb7_71__N_1523_adj_6053[70]), .S1(comb7_71__N_1523_adj_6053[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_35 (.A0(comb6_adj_6025[68]), .B0(cout_adj_5308), 
          .C0(n87_adj_5766), .D0(n5_adj_4877), .A1(comb6_adj_6025[69]), 
          .B1(cout_adj_5308), .C1(n84_adj_5765), .D1(n4_adj_4876), .CIN(n14615), 
          .COUT(n14616), .S0(comb7_71__N_1523_adj_6053[68]), .S1(comb7_71__N_1523_adj_6053[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_33 (.A0(comb6_adj_6025[66]), .B0(cout_adj_5308), 
          .C0(n93_adj_5768), .D0(n7_adj_4879), .A1(comb6_adj_6025[67]), 
          .B1(cout_adj_5308), .C1(n90_adj_5767), .D1(n6_adj_4878), .CIN(n14614), 
          .COUT(n14615), .S0(comb7_71__N_1523_adj_6053[66]), .S1(comb7_71__N_1523_adj_6053[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_31 (.A0(comb6_adj_6025[64]), .B0(cout_adj_5308), 
          .C0(n99_adj_5770), .D0(n9_adj_4881), .A1(comb6_adj_6025[65]), 
          .B1(cout_adj_5308), .C1(n96_adj_5769), .D1(n8_adj_4880), .CIN(n14613), 
          .COUT(n14614), .S0(comb7_71__N_1523_adj_6053[64]), .S1(comb7_71__N_1523_adj_6053[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_29 (.A0(comb6_adj_6025[62]), .B0(cout_adj_5308), 
          .C0(n105_adj_5772), .D0(n11_adj_4883), .A1(comb6_adj_6025[63]), 
          .B1(cout_adj_5308), .C1(n102_adj_5771), .D1(n10_adj_4882), .CIN(n14612), 
          .COUT(n14613), .S0(comb7_71__N_1523_adj_6053[62]), .S1(comb7_71__N_1523_adj_6053[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_27 (.A0(comb6_adj_6025[60]), .B0(cout_adj_5308), 
          .C0(n111_adj_5774), .D0(n13_adj_4885), .A1(comb6_adj_6025[61]), 
          .B1(cout_adj_5308), .C1(n108_adj_5773), .D1(n12_adj_4884), .CIN(n14611), 
          .COUT(n14612), .S0(comb7_71__N_1523_adj_6053[60]), .S1(comb7_71__N_1523_adj_6053[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_25 (.A0(comb6_adj_6025[58]), .B0(cout_adj_5308), 
          .C0(n117_adj_5776), .D0(n15_adj_4887), .A1(comb6_adj_6025[59]), 
          .B1(cout_adj_5308), .C1(n114_adj_5775), .D1(n14_adj_4886), .CIN(n14610), 
          .COUT(n14611), .S0(comb7_71__N_1523_adj_6053[58]), .S1(comb7_71__N_1523_adj_6053[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_23 (.A0(comb6_adj_6025[56]), .B0(cout_adj_5308), 
          .C0(n123_adj_5778), .D0(n17_adj_4889), .A1(comb6_adj_6025[57]), 
          .B1(cout_adj_5308), .C1(n120_adj_5777), .D1(n16_adj_4888), .CIN(n14609), 
          .COUT(n14610), .S0(comb7_71__N_1523_adj_6053[56]), .S1(comb7_71__N_1523_adj_6053[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_21 (.A0(comb6_adj_6025[54]), .B0(cout_adj_5308), 
          .C0(n129_adj_5780), .D0(n19_adj_4891), .A1(comb6_adj_6025[55]), 
          .B1(cout_adj_5308), .C1(n126_adj_5779), .D1(n18_adj_4890), .CIN(n14608), 
          .COUT(n14609), .S0(comb7_71__N_1523_adj_6053[54]), .S1(comb7_71__N_1523_adj_6053[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_19 (.A0(comb6_adj_6025[52]), .B0(cout_adj_5308), 
          .C0(n135_adj_5782), .D0(n21_adj_4893), .A1(comb6_adj_6025[53]), 
          .B1(cout_adj_5308), .C1(n132_adj_5781), .D1(n20_adj_4892), .CIN(n14607), 
          .COUT(n14608), .S0(comb7_71__N_1523_adj_6053[52]), .S1(comb7_71__N_1523_adj_6053[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_17 (.A0(comb6_adj_6025[50]), .B0(cout_adj_5308), 
          .C0(n141_adj_5784), .D0(n23_adj_4895), .A1(comb6_adj_6025[51]), 
          .B1(cout_adj_5308), .C1(n138_adj_5783), .D1(n22_adj_4894), .CIN(n14606), 
          .COUT(n14607), .S0(comb7_71__N_1523_adj_6053[50]), .S1(comb7_71__N_1523_adj_6053[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_15 (.A0(comb6_adj_6025[48]), .B0(cout_adj_5308), 
          .C0(n147_adj_5786), .D0(n25_adj_4897), .A1(comb6_adj_6025[49]), 
          .B1(cout_adj_5308), .C1(n144_adj_5785), .D1(n24_adj_4896), .CIN(n14605), 
          .COUT(n14606), .S0(comb7_71__N_1523_adj_6053[48]), .S1(comb7_71__N_1523_adj_6053[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_13 (.A0(comb6_adj_6025[46]), .B0(cout_adj_5308), 
          .C0(n153_adj_5788), .D0(n27_adj_4899), .A1(comb6_adj_6025[47]), 
          .B1(cout_adj_5308), .C1(n150_adj_5787), .D1(n26_adj_4898), .CIN(n14604), 
          .COUT(n14605), .S0(comb7_71__N_1523_adj_6053[46]), .S1(comb7_71__N_1523_adj_6053[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_11 (.A0(comb6_adj_6025[44]), .B0(cout_adj_5308), 
          .C0(n159_adj_5790), .D0(n29_adj_4901), .A1(comb6_adj_6025[45]), 
          .B1(cout_adj_5308), .C1(n156_adj_5789), .D1(n28_adj_4900), .CIN(n14603), 
          .COUT(n14604), .S0(comb7_71__N_1523_adj_6053[44]), .S1(comb7_71__N_1523_adj_6053[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_9 (.A0(comb6_adj_6025[42]), .B0(cout_adj_5308), 
          .C0(n165_adj_5792), .D0(n31_adj_4903), .A1(comb6_adj_6025[43]), 
          .B1(cout_adj_5308), .C1(n162_adj_5791), .D1(n30_adj_4902), .CIN(n14602), 
          .COUT(n14603), .S0(comb7_71__N_1523_adj_6053[42]), .S1(comb7_71__N_1523_adj_6053[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_7 (.A0(comb6_adj_6025[40]), .B0(cout_adj_5308), 
          .C0(n171_adj_5794), .D0(n33_adj_4905), .A1(comb6_adj_6025[41]), 
          .B1(cout_adj_5308), .C1(n168_adj_5793), .D1(n32_adj_4904), .CIN(n14601), 
          .COUT(n14602), .S0(comb7_71__N_1523_adj_6053[40]), .S1(comb7_71__N_1523_adj_6053[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_5 (.A0(comb6_adj_6025[38]), .B0(cout_adj_5308), 
          .C0(n177_adj_5796), .D0(n35_adj_4907), .A1(comb6_adj_6025[39]), 
          .B1(cout_adj_5308), .C1(n174_adj_5795), .D1(n34_adj_4906), .CIN(n14600), 
          .COUT(n14601), .S0(comb7_71__N_1523_adj_6053[38]), .S1(comb7_71__N_1523_adj_6053[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_3 (.A0(comb6_adj_6025[36]), .B0(cout_adj_5308), 
          .C0(n183_adj_5798), .D0(n37_adj_4909), .A1(comb6_adj_6025[37]), 
          .B1(cout_adj_5308), .C1(n180_adj_5797), .D1(n36_adj_4908), .CIN(n14599), 
          .COUT(n14600), .S0(comb7_71__N_1523_adj_6053[36]), .S1(comb7_71__N_1523_adj_6053[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1082_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1082_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1082_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5308), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14599));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1082_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1082_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1082_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1082_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_37 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n81_adj_4988), .D0(integrator1_adj_6020[70]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n78_adj_4987), .D1(integrator1_adj_6020[71]), 
          .CIN(n14594), .S0(integrator1_71__N_418_adj_6036[70]), .S1(integrator1_71__N_418_adj_6036[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_35 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n87_adj_4990), .D0(integrator1_adj_6020[68]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n84_adj_4989), .D1(integrator1_adj_6020[69]), 
          .CIN(n14593), .COUT(n14594), .S0(integrator1_71__N_418_adj_6036[68]), 
          .S1(integrator1_71__N_418_adj_6036[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_33 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n93_adj_4992), .D0(integrator1_adj_6020[66]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n90_adj_4991), .D1(integrator1_adj_6020[67]), 
          .CIN(n14592), .COUT(n14593), .S0(integrator1_71__N_418_adj_6036[66]), 
          .S1(integrator1_71__N_418_adj_6036[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_31 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n99_adj_4994), .D0(integrator1_adj_6020[64]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n96_adj_4993), .D1(integrator1_adj_6020[65]), 
          .CIN(n14591), .COUT(n14592), .S0(integrator1_71__N_418_adj_6036[64]), 
          .S1(integrator1_71__N_418_adj_6036[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_29 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n105_adj_4996), .D0(integrator1_adj_6020[62]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n102_adj_4995), .D1(integrator1_adj_6020[63]), 
          .CIN(n14590), .COUT(n14591), .S0(integrator1_71__N_418_adj_6036[62]), 
          .S1(integrator1_71__N_418_adj_6036[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_27 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n111_adj_4998), .D0(integrator1_adj_6020[60]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n108_adj_4997), .D1(integrator1_adj_6020[61]), 
          .CIN(n14589), .COUT(n14590), .S0(integrator1_71__N_418_adj_6036[60]), 
          .S1(integrator1_71__N_418_adj_6036[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_25 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n117_adj_5000), .D0(integrator1_adj_6020[58]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n114_adj_4999), .D1(integrator1_adj_6020[59]), 
          .CIN(n14588), .COUT(n14589), .S0(integrator1_71__N_418_adj_6036[58]), 
          .S1(integrator1_71__N_418_adj_6036[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_23 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n123_adj_5002), .D0(integrator1_adj_6020[56]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n120_adj_5001), .D1(integrator1_adj_6020[57]), 
          .CIN(n14587), .COUT(n14588), .S0(integrator1_71__N_418_adj_6036[56]), 
          .S1(integrator1_71__N_418_adj_6036[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_21 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n129_adj_5004), .D0(integrator1_adj_6020[54]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n126_adj_5003), .D1(integrator1_adj_6020[55]), 
          .CIN(n14586), .COUT(n14587), .S0(integrator1_71__N_418_adj_6036[54]), 
          .S1(integrator1_71__N_418_adj_6036[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_19 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n135_adj_5006), .D0(integrator1_adj_6020[52]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n132_adj_5005), .D1(integrator1_adj_6020[53]), 
          .CIN(n14585), .COUT(n14586), .S0(integrator1_71__N_418_adj_6036[52]), 
          .S1(integrator1_71__N_418_adj_6036[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_17 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n141_adj_5008), .D0(integrator1_adj_6020[50]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n138_adj_5007), .D1(integrator1_adj_6020[51]), 
          .CIN(n14584), .COUT(n14585), .S0(integrator1_71__N_418_adj_6036[50]), 
          .S1(integrator1_71__N_418_adj_6036[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_15 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n147_adj_5010), .D0(integrator1_adj_6020[48]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n144_adj_5009), .D1(integrator1_adj_6020[49]), 
          .CIN(n14583), .COUT(n14584), .S0(integrator1_71__N_418_adj_6036[48]), 
          .S1(integrator1_71__N_418_adj_6036[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_13 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n153_adj_5012), .D0(integrator1_adj_6020[46]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n150_adj_5011), .D1(integrator1_adj_6020[47]), 
          .CIN(n14582), .COUT(n14583), .S0(integrator1_71__N_418_adj_6036[46]), 
          .S1(integrator1_71__N_418_adj_6036[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_11 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n159_adj_5014), .D0(integrator1_adj_6020[44]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n156_adj_5013), .D1(integrator1_adj_6020[45]), 
          .CIN(n14581), .COUT(n14582), .S0(integrator1_71__N_418_adj_6036[44]), 
          .S1(integrator1_71__N_418_adj_6036[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_9 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n165_adj_5016), .D0(integrator1_adj_6020[42]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n162_adj_5015), .D1(integrator1_adj_6020[43]), 
          .CIN(n14580), .COUT(n14581), .S0(integrator1_71__N_418_adj_6036[42]), 
          .S1(integrator1_71__N_418_adj_6036[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_7 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n171_adj_5018), .D0(integrator1_adj_6020[40]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n168_adj_5017), .D1(integrator1_adj_6020[41]), 
          .CIN(n14579), .COUT(n14580), .S0(integrator1_71__N_418_adj_6036[40]), 
          .S1(integrator1_71__N_418_adj_6036[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_5 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n177_adj_5020), .D0(integrator1_adj_6020[38]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n174_adj_5019), .D1(integrator1_adj_6020[39]), 
          .CIN(n14578), .COUT(n14579), .S0(integrator1_71__N_418_adj_6036[38]), 
          .S1(integrator1_71__N_418_adj_6036[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_3 (.A0(mix_cosinewave[11]), .B0(cout_adj_5076), 
          .C0(n183_adj_5022), .D0(integrator1_adj_6020[36]), .A1(mix_cosinewave[11]), 
          .B1(cout_adj_5076), .C1(n180_adj_5021), .D1(integrator1_adj_6020[37]), 
          .CIN(n14577), .COUT(n14578), .S0(integrator1_71__N_418_adj_6036[36]), 
          .S1(integrator1_71__N_418_adj_6036[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1106_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1106_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1106_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5076), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14577));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1106_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1106_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1106_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1106_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_38 (.A0(comb_d7_adj_6028[35]), .B0(comb7_adj_6027[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14573), .S0(comb8_71__N_1595_adj_6054[35]), 
          .S1(cout_adj_5309));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1175_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_36 (.A0(comb_d7_adj_6028[33]), .B0(comb7_adj_6027[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[34]), .B1(comb7_adj_6027[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14572), .COUT(n14573), .S0(comb8_71__N_1595_adj_6054[33]), 
          .S1(comb8_71__N_1595_adj_6054[34]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_34 (.A0(comb_d7_adj_6028[31]), .B0(comb7_adj_6027[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[32]), .B1(comb7_adj_6027[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14571), .COUT(n14572), .S0(comb8_71__N_1595_adj_6054[31]), 
          .S1(comb8_71__N_1595_adj_6054[32]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_32 (.A0(comb_d7_adj_6028[29]), .B0(comb7_adj_6027[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[30]), .B1(comb7_adj_6027[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14570), .COUT(n14571), .S0(comb8_71__N_1595_adj_6054[29]), 
          .S1(comb8_71__N_1595_adj_6054[30]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_30 (.A0(comb_d7_adj_6028[27]), .B0(comb7_adj_6027[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[28]), .B1(comb7_adj_6027[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14569), .COUT(n14570), .S0(comb8_71__N_1595_adj_6054[27]), 
          .S1(comb8_71__N_1595_adj_6054[28]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_28 (.A0(comb_d7_adj_6028[25]), .B0(comb7_adj_6027[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[26]), .B1(comb7_adj_6027[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14568), .COUT(n14569), .S0(comb8_71__N_1595_adj_6054[25]), 
          .S1(comb8_71__N_1595_adj_6054[26]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_26 (.A0(comb_d7_adj_6028[23]), .B0(comb7_adj_6027[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[24]), .B1(comb7_adj_6027[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14567), .COUT(n14568), .S0(comb8_71__N_1595_adj_6054[23]), 
          .S1(comb8_71__N_1595_adj_6054[24]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_24 (.A0(comb_d7_adj_6028[21]), .B0(comb7_adj_6027[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[22]), .B1(comb7_adj_6027[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14566), .COUT(n14567), .S0(comb8_71__N_1595_adj_6054[21]), 
          .S1(comb8_71__N_1595_adj_6054[22]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_22 (.A0(comb_d7_adj_6028[19]), .B0(comb7_adj_6027[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[20]), .B1(comb7_adj_6027[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14565), .COUT(n14566), .S0(comb8_71__N_1595_adj_6054[19]), 
          .S1(comb8_71__N_1595_adj_6054[20]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_20 (.A0(comb_d7_adj_6028[17]), .B0(comb7_adj_6027[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[18]), .B1(comb7_adj_6027[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14564), .COUT(n14565), .S0(comb8_71__N_1595_adj_6054[17]), 
          .S1(comb8_71__N_1595_adj_6054[18]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_18 (.A0(comb_d7_adj_6028[15]), .B0(comb7_adj_6027[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[16]), .B1(comb7_adj_6027[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14563), .COUT(n14564), .S0(comb8_71__N_1595_adj_6054[15]), 
          .S1(comb8_71__N_1595_adj_6054[16]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_16 (.A0(comb_d7_adj_6028[13]), .B0(comb7_adj_6027[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[14]), .B1(comb7_adj_6027[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14562), .COUT(n14563), .S0(comb8_71__N_1595_adj_6054[13]), 
          .S1(comb8_71__N_1595_adj_6054[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_14 (.A0(comb_d7_adj_6028[11]), .B0(comb7_adj_6027[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[12]), .B1(comb7_adj_6027[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14561), .COUT(n14562), .S0(comb8_71__N_1595_adj_6054[11]), 
          .S1(comb8_71__N_1595_adj_6054[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_12 (.A0(comb_d7_adj_6028[9]), .B0(comb7_adj_6027[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[10]), .B1(comb7_adj_6027[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14560), .COUT(n14561), .S0(comb8_71__N_1595_adj_6054[9]), 
          .S1(comb8_71__N_1595_adj_6054[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_10 (.A0(comb_d7_adj_6028[7]), .B0(comb7_adj_6027[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[8]), .B1(comb7_adj_6027[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14559), .COUT(n14560), .S0(comb8_71__N_1595_adj_6054[7]), 
          .S1(comb8_71__N_1595_adj_6054[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_8 (.A0(comb_d7_adj_6028[5]), .B0(comb7_adj_6027[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[6]), .B1(comb7_adj_6027[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14558), .COUT(n14559), .S0(comb8_71__N_1595_adj_6054[5]), 
          .S1(comb8_71__N_1595_adj_6054[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_6 (.A0(comb_d7_adj_6028[3]), .B0(comb7_adj_6027[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[4]), .B1(comb7_adj_6027[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14557), .COUT(n14558), .S0(comb8_71__N_1595_adj_6054[3]), 
          .S1(comb8_71__N_1595_adj_6054[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_4 (.A0(comb_d7_adj_6028[1]), .B0(comb7_adj_6027[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[2]), .B1(comb7_adj_6027[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14556), .COUT(n14557), .S0(comb8_71__N_1595_adj_6054[1]), 
          .S1(comb8_71__N_1595_adj_6054[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1175_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1175_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7_adj_6028[0]), .B1(comb7_adj_6027[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14556), .S1(comb8_71__N_1595_adj_6054[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1175_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1175_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1175_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1175_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_38 (.A0(integrator_d_tmp[71]), .B0(integrator_tmp[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14555), .S0(n78_adj_5425));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1211_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_36 (.A0(integrator_d_tmp[69]), .B0(integrator_tmp[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[70]), .B1(integrator_tmp[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14554), .COUT(n14555), .S0(n84_adj_5427), 
          .S1(n81_adj_5426));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_34 (.A0(integrator_d_tmp[67]), .B0(integrator_tmp[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[68]), .B1(integrator_tmp[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14553), .COUT(n14554), .S0(n90_adj_5429), 
          .S1(n87_adj_5428));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_32 (.A0(integrator_d_tmp[65]), .B0(integrator_tmp[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[66]), .B1(integrator_tmp[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14552), .COUT(n14553), .S0(n96_adj_5431), 
          .S1(n93_adj_5430));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_30 (.A0(integrator_d_tmp[63]), .B0(integrator_tmp[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[64]), .B1(integrator_tmp[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14551), .COUT(n14552), .S0(n102_adj_5433), 
          .S1(n99_adj_5432));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_28 (.A0(integrator_d_tmp[61]), .B0(integrator_tmp[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[62]), .B1(integrator_tmp[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14550), .COUT(n14551), .S0(n108_adj_5435), 
          .S1(n105_adj_5434));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_26 (.A0(integrator_d_tmp[59]), .B0(integrator_tmp[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[60]), .B1(integrator_tmp[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14549), .COUT(n14550), .S0(n114_adj_5437), 
          .S1(n111_adj_5436));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_24 (.A0(integrator_d_tmp[57]), .B0(integrator_tmp[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[58]), .B1(integrator_tmp[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14548), .COUT(n14549), .S0(n120_adj_5439), 
          .S1(n117_adj_5438));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_22 (.A0(integrator_d_tmp[55]), .B0(integrator_tmp[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[56]), .B1(integrator_tmp[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14547), .COUT(n14548), .S0(n126_adj_5441), 
          .S1(n123_adj_5440));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_20 (.A0(integrator_d_tmp[53]), .B0(integrator_tmp[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[54]), .B1(integrator_tmp[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14546), .COUT(n14547), .S0(n132_adj_5443), 
          .S1(n129_adj_5442));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_18 (.A0(integrator_d_tmp[51]), .B0(integrator_tmp[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[52]), .B1(integrator_tmp[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14545), .COUT(n14546), .S0(n138_adj_5445), 
          .S1(n135_adj_5444));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_16 (.A0(integrator_d_tmp[49]), .B0(integrator_tmp[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[50]), .B1(integrator_tmp[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14544), .COUT(n14545), .S0(n144_adj_5447), 
          .S1(n141_adj_5446));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_14 (.A0(integrator_d_tmp[47]), .B0(integrator_tmp[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[48]), .B1(integrator_tmp[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14543), .COUT(n14544), .S0(n150_adj_5449), 
          .S1(n147_adj_5448));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_12 (.A0(integrator_d_tmp[45]), .B0(integrator_tmp[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[46]), .B1(integrator_tmp[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14542), .COUT(n14543), .S0(n156_adj_5451), 
          .S1(n153_adj_5450));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_10 (.A0(integrator_d_tmp[43]), .B0(integrator_tmp[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[44]), .B1(integrator_tmp[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14541), .COUT(n14542), .S0(n162_adj_5453), 
          .S1(n159_adj_5452));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_8 (.A0(integrator_d_tmp[41]), .B0(integrator_tmp[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[42]), .B1(integrator_tmp[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14540), .COUT(n14541), .S0(n168_adj_5455), 
          .S1(n165_adj_5454));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_6 (.A0(integrator_d_tmp[39]), .B0(integrator_tmp[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[40]), .B1(integrator_tmp[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14539), .COUT(n14540), .S0(n174_adj_5457), 
          .S1(n171_adj_5456));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_4 (.A0(integrator_d_tmp[37]), .B0(integrator_tmp[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[38]), .B1(integrator_tmp[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14538), .COUT(n14539), .S0(n180_adj_5459), 
          .S1(n177_adj_5458));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1211_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1211_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator_d_tmp[36]), .B1(integrator_tmp[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14538), .S1(n183_adj_5460));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1211_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1211_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1211_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1211_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_37 (.A0(integrator4[70]), .B0(cout_adj_5075), 
          .C0(n81_adj_5128), .D0(integrator5[70]), .A1(integrator4[71]), 
          .B1(cout_adj_5075), .C1(n78_adj_5127), .D1(integrator5[71]), 
          .CIN(n14536), .S0(integrator5_71__N_706[70]), .S1(integrator5_71__N_706[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_35 (.A0(integrator4[68]), .B0(cout_adj_5075), 
          .C0(n87_adj_5130), .D0(integrator5[68]), .A1(integrator4[69]), 
          .B1(cout_adj_5075), .C1(n84_adj_5129), .D1(integrator5[69]), 
          .CIN(n14535), .COUT(n14536), .S0(integrator5_71__N_706[68]), 
          .S1(integrator5_71__N_706[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_33 (.A0(integrator4[66]), .B0(cout_adj_5075), 
          .C0(n93_adj_5132), .D0(integrator5[66]), .A1(integrator4[67]), 
          .B1(cout_adj_5075), .C1(n90_adj_5131), .D1(integrator5[67]), 
          .CIN(n14534), .COUT(n14535), .S0(integrator5_71__N_706[66]), 
          .S1(integrator5_71__N_706[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_31 (.A0(integrator4[64]), .B0(cout_adj_5075), 
          .C0(n99_adj_5134), .D0(integrator5[64]), .A1(integrator4[65]), 
          .B1(cout_adj_5075), .C1(n96_adj_5133), .D1(integrator5[65]), 
          .CIN(n14533), .COUT(n14534), .S0(integrator5_71__N_706[64]), 
          .S1(integrator5_71__N_706[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_29 (.A0(integrator4[62]), .B0(cout_adj_5075), 
          .C0(n105_adj_5136), .D0(integrator5[62]), .A1(integrator4[63]), 
          .B1(cout_adj_5075), .C1(n102_adj_5135), .D1(integrator5[63]), 
          .CIN(n14532), .COUT(n14533), .S0(integrator5_71__N_706[62]), 
          .S1(integrator5_71__N_706[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_27 (.A0(integrator4[60]), .B0(cout_adj_5075), 
          .C0(n111_adj_5138), .D0(integrator5[60]), .A1(integrator4[61]), 
          .B1(cout_adj_5075), .C1(n108_adj_5137), .D1(integrator5[61]), 
          .CIN(n14531), .COUT(n14532), .S0(integrator5_71__N_706[60]), 
          .S1(integrator5_71__N_706[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_25 (.A0(integrator4[58]), .B0(cout_adj_5075), 
          .C0(n117_adj_5140), .D0(integrator5[58]), .A1(integrator4[59]), 
          .B1(cout_adj_5075), .C1(n114_adj_5139), .D1(integrator5[59]), 
          .CIN(n14530), .COUT(n14531), .S0(integrator5_71__N_706[58]), 
          .S1(integrator5_71__N_706[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_23 (.A0(integrator4[56]), .B0(cout_adj_5075), 
          .C0(n123_adj_5142), .D0(integrator5[56]), .A1(integrator4[57]), 
          .B1(cout_adj_5075), .C1(n120_adj_5141), .D1(integrator5[57]), 
          .CIN(n14529), .COUT(n14530), .S0(integrator5_71__N_706[56]), 
          .S1(integrator5_71__N_706[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_21 (.A0(integrator4[54]), .B0(cout_adj_5075), 
          .C0(n129_adj_5144), .D0(integrator5[54]), .A1(integrator4[55]), 
          .B1(cout_adj_5075), .C1(n126_adj_5143), .D1(integrator5[55]), 
          .CIN(n14528), .COUT(n14529), .S0(integrator5_71__N_706[54]), 
          .S1(integrator5_71__N_706[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_19 (.A0(integrator4[52]), .B0(cout_adj_5075), 
          .C0(n135_adj_5146), .D0(integrator5[52]), .A1(integrator4[53]), 
          .B1(cout_adj_5075), .C1(n132_adj_5145), .D1(integrator5[53]), 
          .CIN(n14527), .COUT(n14528), .S0(integrator5_71__N_706[52]), 
          .S1(integrator5_71__N_706[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_17 (.A0(integrator4[50]), .B0(cout_adj_5075), 
          .C0(n141_adj_5148), .D0(integrator5[50]), .A1(integrator4[51]), 
          .B1(cout_adj_5075), .C1(n138_adj_5147), .D1(integrator5[51]), 
          .CIN(n14526), .COUT(n14527), .S0(integrator5_71__N_706[50]), 
          .S1(integrator5_71__N_706[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_15 (.A0(integrator4[48]), .B0(cout_adj_5075), 
          .C0(n147_adj_5150), .D0(integrator5[48]), .A1(integrator4[49]), 
          .B1(cout_adj_5075), .C1(n144_adj_5149), .D1(integrator5[49]), 
          .CIN(n14525), .COUT(n14526), .S0(integrator5_71__N_706[48]), 
          .S1(integrator5_71__N_706[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_13 (.A0(integrator4[46]), .B0(cout_adj_5075), 
          .C0(n153_adj_5152), .D0(integrator5[46]), .A1(integrator4[47]), 
          .B1(cout_adj_5075), .C1(n150_adj_5151), .D1(integrator5[47]), 
          .CIN(n14524), .COUT(n14525), .S0(integrator5_71__N_706[46]), 
          .S1(integrator5_71__N_706[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_11 (.A0(integrator4[44]), .B0(cout_adj_5075), 
          .C0(n159_adj_5154), .D0(integrator5[44]), .A1(integrator4[45]), 
          .B1(cout_adj_5075), .C1(n156_adj_5153), .D1(integrator5[45]), 
          .CIN(n14523), .COUT(n14524), .S0(integrator5_71__N_706[44]), 
          .S1(integrator5_71__N_706[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_9 (.A0(integrator4[42]), .B0(cout_adj_5075), 
          .C0(n165_adj_5156), .D0(integrator5[42]), .A1(integrator4[43]), 
          .B1(cout_adj_5075), .C1(n162_adj_5155), .D1(integrator5[43]), 
          .CIN(n14522), .COUT(n14523), .S0(integrator5_71__N_706[42]), 
          .S1(integrator5_71__N_706[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_7 (.A0(integrator4[40]), .B0(cout_adj_5075), 
          .C0(n171_adj_5158), .D0(integrator5[40]), .A1(integrator4[41]), 
          .B1(cout_adj_5075), .C1(n168_adj_5157), .D1(integrator5[41]), 
          .CIN(n14521), .COUT(n14522), .S0(integrator5_71__N_706[40]), 
          .S1(integrator5_71__N_706[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_5 (.A0(integrator4[38]), .B0(cout_adj_5075), 
          .C0(n177_adj_5160), .D0(integrator5[38]), .A1(integrator4[39]), 
          .B1(cout_adj_5075), .C1(n174_adj_5159), .D1(integrator5[39]), 
          .CIN(n14520), .COUT(n14521), .S0(integrator5_71__N_706[38]), 
          .S1(integrator5_71__N_706[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_3 (.A0(integrator4[36]), .B0(cout_adj_5075), 
          .C0(n183_adj_5162), .D0(integrator5[36]), .A1(integrator4[37]), 
          .B1(cout_adj_5075), .C1(n180_adj_5161), .D1(integrator5[37]), 
          .CIN(n14519), .COUT(n14520), .S0(integrator5_71__N_706[36]), 
          .S1(integrator5_71__N_706[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1043_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1043_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1043_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5075), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14519));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1043_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1043_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1043_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1043_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_38 (.A0(integrator1[71]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14513), .S0(n78_adj_5353));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1205_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_36 (.A0(integrator1[69]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[70]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14512), .COUT(n14513), .S0(n84_adj_5355), 
          .S1(n81_adj_5354));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_34 (.A0(integrator1[67]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[68]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14511), .COUT(n14512), .S0(n90_adj_5357), 
          .S1(n87_adj_5356));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_32 (.A0(integrator1[65]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[66]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14510), .COUT(n14511), .S0(n96_adj_5359), 
          .S1(n93_adj_5358));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_30 (.A0(integrator1[63]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[64]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14509), .COUT(n14510), .S0(n102_adj_5361), 
          .S1(n99_adj_5360));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_28 (.A0(integrator1[61]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[62]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14508), .COUT(n14509), .S0(n108_adj_5363), 
          .S1(n105_adj_5362));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_26 (.A0(integrator1[59]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[60]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14507), .COUT(n14508), .S0(n114_adj_5365), 
          .S1(n111_adj_5364));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_24 (.A0(integrator1[57]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[58]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14506), .COUT(n14507), .S0(n120_adj_5367), 
          .S1(n117_adj_5366));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_22 (.A0(integrator1[55]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[56]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14505), .COUT(n14506), .S0(n126_adj_5369), 
          .S1(n123_adj_5368));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_20 (.A0(integrator1[53]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[54]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14504), .COUT(n14505), .S0(n132_adj_5371), 
          .S1(n129_adj_5370));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_18 (.A0(integrator1[51]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[52]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14503), .COUT(n14504), .S0(n138_adj_5373), 
          .S1(n135_adj_5372));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_16 (.A0(integrator1[49]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[50]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14502), .COUT(n14503), .S0(n144_adj_5375), 
          .S1(n141_adj_5374));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_14 (.A0(integrator1[47]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[48]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14501), .COUT(n14502), .S0(n150_adj_5377), 
          .S1(n147_adj_5376));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_12 (.A0(integrator1[45]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[46]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14500), .COUT(n14501), .S0(n156_adj_5379), 
          .S1(n153_adj_5378));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_10 (.A0(integrator1[43]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[44]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14499), .COUT(n14500), .S0(n162_adj_5381), 
          .S1(n159_adj_5380));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_8 (.A0(integrator1[41]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[42]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14498), .COUT(n14499), .S0(n168_adj_5383), 
          .S1(n165_adj_5382));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_6 (.A0(integrator1[39]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[40]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14497), .COUT(n14498), .S0(n174_adj_5385), 
          .S1(n171_adj_5384));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_4 (.A0(integrator1[37]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[38]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14496), .COUT(n14497), .S0(n180_adj_5387), 
          .S1(n177_adj_5386));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1205_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1205_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator1[36]), .B1(mix_sinewave[11]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14496), .S1(n183_adj_5388));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1205_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1205_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1205_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1205_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1220_add_4_16 (.A0(amdemod_d_11__N_1861[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14495), .S0(n34_adj_5483));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1220_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1220_add_4_16.INIT1 = 16'h0000;
    defparam _add_1_1220_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1220_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1220_add_4_14 (.A0(amdemod_d_11__N_1861[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1861[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14494), .COUT(n14495), .S0(n40_adj_5484));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1220_add_4_14.INIT0 = 16'h555f;
    defparam _add_1_1220_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_1220_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1220_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1220_add_4_12 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1861[7]), .D0(VCC_net), .A1(amdemod_d_11__N_1861[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n14493), .COUT(n14494), 
          .S0(n46_adj_5486), .S1(n43_adj_5485));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1220_add_4_12.INIT0 = 16'he1e1;
    defparam _add_1_1220_add_4_12.INIT1 = 16'h555f;
    defparam _add_1_1220_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1220_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1220_add_4_10 (.A0(n17134), .B0(amdemod_d_11__N_1861[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17137), .B1(amdemod_d_11__N_1861[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14492), .COUT(n14493), .S0(n52_adj_5488), 
          .S1(n49_adj_5487));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1220_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1220_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1220_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1220_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1220_add_4_8 (.A0(n17132), .B0(amdemod_d_11__N_1861[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1861[4]), .B1(amdemod_d_11__N_1841[11]), 
          .C1(n17134), .D1(amdemod_d_11__N_1840[11]), .CIN(n14491), .COUT(n14492), 
          .S0(n58_adj_5490), .S1(n55_adj_5489));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1220_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1220_add_4_8.INIT1 = 16'h656a;
    defparam _add_1_1220_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1220_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1220_add_4_6 (.A0(n17130), .B0(amdemod_d_11__N_1861[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1861[2]), .B1(amdemod_d_11__N_1851[13]), 
          .C1(n17132), .D1(amdemod_d_11__N_1850[13]), .CIN(n14490), .COUT(n14491), 
          .S0(n64_adj_5492), .S1(n61_adj_5491));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1220_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1220_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_1220_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1220_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1220_add_4_4 (.A0(n17129), .B0(square_sum[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_d_11__N_1861[0]), .B1(amdemod_d_11__N_1861[13]), 
          .C1(n17130), .D1(amdemod_d_11__N_1860[13]), .CIN(n14489), .COUT(n14490), 
          .S0(n70_adj_5494), .S1(n67_adj_5493));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1220_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1220_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_1220_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1220_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1220_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14489), .S1(n73_adj_5495));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1220_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1220_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1220_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1220_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_38 (.A0(comb_d8_adj_6030[35]), .B0(comb8_adj_6029[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14488), .S0(comb9_71__N_1667_adj_6055[35]), 
          .S1(cout_adj_5310));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1178_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_36 (.A0(comb_d8_adj_6030[33]), .B0(comb8_adj_6029[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[34]), .B1(comb8_adj_6029[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14487), .COUT(n14488), .S0(comb9_71__N_1667_adj_6055[33]), 
          .S1(comb9_71__N_1667_adj_6055[34]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_34 (.A0(comb_d8_adj_6030[31]), .B0(comb8_adj_6029[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[32]), .B1(comb8_adj_6029[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14486), .COUT(n14487), .S0(comb9_71__N_1667_adj_6055[31]), 
          .S1(comb9_71__N_1667_adj_6055[32]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_32 (.A0(comb_d8_adj_6030[29]), .B0(comb8_adj_6029[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[30]), .B1(comb8_adj_6029[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14485), .COUT(n14486), .S0(comb9_71__N_1667_adj_6055[29]), 
          .S1(comb9_71__N_1667_adj_6055[30]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_30 (.A0(comb_d8_adj_6030[27]), .B0(comb8_adj_6029[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[28]), .B1(comb8_adj_6029[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14484), .COUT(n14485), .S0(comb9_71__N_1667_adj_6055[27]), 
          .S1(comb9_71__N_1667_adj_6055[28]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_28 (.A0(comb_d8_adj_6030[25]), .B0(comb8_adj_6029[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[26]), .B1(comb8_adj_6029[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14483), .COUT(n14484), .S0(comb9_71__N_1667_adj_6055[25]), 
          .S1(comb9_71__N_1667_adj_6055[26]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_26 (.A0(comb_d8_adj_6030[23]), .B0(comb8_adj_6029[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[24]), .B1(comb8_adj_6029[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14482), .COUT(n14483), .S0(comb9_71__N_1667_adj_6055[23]), 
          .S1(comb9_71__N_1667_adj_6055[24]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_24 (.A0(comb_d8_adj_6030[21]), .B0(comb8_adj_6029[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[22]), .B1(comb8_adj_6029[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14481), .COUT(n14482), .S0(comb9_71__N_1667_adj_6055[21]), 
          .S1(comb9_71__N_1667_adj_6055[22]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_22 (.A0(comb_d8_adj_6030[19]), .B0(comb8_adj_6029[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[20]), .B1(comb8_adj_6029[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14480), .COUT(n14481), .S0(comb9_71__N_1667_adj_6055[19]), 
          .S1(comb9_71__N_1667_adj_6055[20]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_20 (.A0(comb_d8_adj_6030[17]), .B0(comb8_adj_6029[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[18]), .B1(comb8_adj_6029[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14479), .COUT(n14480), .S0(comb9_71__N_1667_adj_6055[17]), 
          .S1(comb9_71__N_1667_adj_6055[18]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_18 (.A0(comb_d8_adj_6030[15]), .B0(comb8_adj_6029[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[16]), .B1(comb8_adj_6029[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14478), .COUT(n14479), .S0(comb9_71__N_1667_adj_6055[15]), 
          .S1(comb9_71__N_1667_adj_6055[16]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_16 (.A0(comb_d8_adj_6030[13]), .B0(comb8_adj_6029[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[14]), .B1(comb8_adj_6029[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14477), .COUT(n14478), .S0(comb9_71__N_1667_adj_6055[13]), 
          .S1(comb9_71__N_1667_adj_6055[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_14 (.A0(comb_d8_adj_6030[11]), .B0(comb8_adj_6029[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[12]), .B1(comb8_adj_6029[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14476), .COUT(n14477), .S0(comb9_71__N_1667_adj_6055[11]), 
          .S1(comb9_71__N_1667_adj_6055[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_12 (.A0(comb_d8_adj_6030[9]), .B0(comb8_adj_6029[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[10]), .B1(comb8_adj_6029[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14475), .COUT(n14476), .S0(comb9_71__N_1667_adj_6055[9]), 
          .S1(comb9_71__N_1667_adj_6055[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_10 (.A0(comb_d8_adj_6030[7]), .B0(comb8_adj_6029[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[8]), .B1(comb8_adj_6029[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14474), .COUT(n14475), .S0(comb9_71__N_1667_adj_6055[7]), 
          .S1(comb9_71__N_1667_adj_6055[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_8 (.A0(comb_d8_adj_6030[5]), .B0(comb8_adj_6029[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[6]), .B1(comb8_adj_6029[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14473), .COUT(n14474), .S0(comb9_71__N_1667_adj_6055[5]), 
          .S1(comb9_71__N_1667_adj_6055[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_6 (.A0(comb_d8_adj_6030[3]), .B0(comb8_adj_6029[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[4]), .B1(comb8_adj_6029[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14472), .COUT(n14473), .S0(comb9_71__N_1667_adj_6055[3]), 
          .S1(comb9_71__N_1667_adj_6055[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_4 (.A0(comb_d8_adj_6030[1]), .B0(comb8_adj_6029[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[2]), .B1(comb8_adj_6029[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14471), .COUT(n14472), .S0(comb9_71__N_1667_adj_6055[1]), 
          .S1(comb9_71__N_1667_adj_6055[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1178_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1178_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8_adj_6030[0]), .B1(comb8_adj_6029[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14471), .S1(comb9_71__N_1667_adj_6055[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1178_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1178_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1178_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1178_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_37 (.A0(comb_d9_adj_6032[71]), .B0(comb9_adj_6031[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14470), .S0(n76_adj_5496));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_37.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_37.INIT1 = 16'h0000;
    defparam _add_1_1091_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_35 (.A0(comb_d9_adj_6032[69]), .B0(comb9_adj_6031[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[70]), .B1(comb9_adj_6031[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14469), .COUT(n14470), .S0(n82), 
          .S1(n79_adj_5497));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_35.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_35.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_33 (.A0(comb_d9_adj_6032[67]), .B0(comb9_adj_6031[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[68]), .B1(comb9_adj_6031[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14468), .COUT(n14469), .S0(n88), 
          .S1(n85));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_33.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_33.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_31 (.A0(comb_d9_adj_6032[65]), .B0(comb9_adj_6031[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[66]), .B1(comb9_adj_6031[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14467), .COUT(n14468), .S0(n94), 
          .S1(n91));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_31.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_31.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_29 (.A0(comb_d9_adj_6032[63]), .B0(comb9_adj_6031[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[64]), .B1(comb9_adj_6031[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14466), .COUT(n14467), .S0(n100), 
          .S1(n97));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_29.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_29.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_27 (.A0(comb_d9_adj_6032[61]), .B0(comb9_adj_6031[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[62]), .B1(comb9_adj_6031[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14465), .COUT(n14466), .S0(n106), 
          .S1(n103));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_27.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_27.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_25 (.A0(comb_d9_adj_6032[59]), .B0(comb9_adj_6031[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[60]), .B1(comb9_adj_6031[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14464), .COUT(n14465), .S0(n112), 
          .S1(n109));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_25.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_25.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_23 (.A0(comb_d9_adj_6032[57]), .B0(comb9_adj_6031[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[58]), .B1(comb9_adj_6031[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14463), .COUT(n14464), .S0(n118), 
          .S1(n115));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_23.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_23.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_21 (.A0(comb_d9_adj_6032[55]), .B0(comb9_adj_6031[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[56]), .B1(comb9_adj_6031[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14462), .COUT(n14463));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_21.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_21.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_19 (.A0(comb_d9_adj_6032[53]), .B0(comb9_adj_6031[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[54]), .B1(comb9_adj_6031[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14461), .COUT(n14462));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_19.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_19.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_17 (.A0(comb_d9_adj_6032[51]), .B0(comb9_adj_6031[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[52]), .B1(comb9_adj_6031[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14460), .COUT(n14461));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_17.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_17.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_15 (.A0(comb_d9_adj_6032[49]), .B0(comb9_adj_6031[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[50]), .B1(comb9_adj_6031[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14459), .COUT(n14460));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_15.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_15.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_13 (.A0(comb_d9_adj_6032[47]), .B0(comb9_adj_6031[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[48]), .B1(comb9_adj_6031[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14458), .COUT(n14459));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_13.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_13.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_11 (.A0(comb_d9_adj_6032[45]), .B0(comb9_adj_6031[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[46]), .B1(comb9_adj_6031[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14457), .COUT(n14458));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_11.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_9 (.A0(comb_d9_adj_6032[43]), .B0(comb9_adj_6031[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[44]), .B1(comb9_adj_6031[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14456), .COUT(n14457));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_7 (.A0(comb_d9_adj_6032[41]), .B0(comb9_adj_6031[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[42]), .B1(comb9_adj_6031[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14455), .COUT(n14456));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_5 (.A0(comb_d9_adj_6032[39]), .B0(comb9_adj_6031[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[40]), .B1(comb9_adj_6031[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14454), .COUT(n14455));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_3 (.A0(comb_d9_adj_6032[37]), .B0(comb9_adj_6031[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[38]), .B1(comb9_adj_6031[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14453), .COUT(n14454));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_3.INIT0 = 16'h9995;
    defparam _add_1_1091_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1091_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9_adj_6032[36]), .B1(comb9_adj_6031[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14453));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1091_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1091_add_4_1.INIT1 = 16'h9995;
    defparam _add_1_1091_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1091_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_38 (.A0(integrator4_adj_6023[71]), .B0(integrator3_adj_6022[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14452), .S0(n78_adj_5498));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1133_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_36 (.A0(integrator4_adj_6023[69]), .B0(integrator3_adj_6022[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[70]), .B1(integrator3_adj_6022[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14451), .COUT(n14452), .S0(n84_adj_5500), 
          .S1(n81_adj_5499));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_34 (.A0(integrator4_adj_6023[67]), .B0(integrator3_adj_6022[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[68]), .B1(integrator3_adj_6022[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14450), .COUT(n14451), .S0(n90_adj_5502), 
          .S1(n87_adj_5501));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_32 (.A0(integrator4_adj_6023[65]), .B0(integrator3_adj_6022[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[66]), .B1(integrator3_adj_6022[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14449), .COUT(n14450), .S0(n96_adj_5504), 
          .S1(n93_adj_5503));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_30 (.A0(integrator4_adj_6023[63]), .B0(integrator3_adj_6022[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[64]), .B1(integrator3_adj_6022[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14448), .COUT(n14449), .S0(n102_adj_5506), 
          .S1(n99_adj_5505));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_28 (.A0(integrator4_adj_6023[61]), .B0(integrator3_adj_6022[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[62]), .B1(integrator3_adj_6022[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14447), .COUT(n14448), .S0(n108_adj_5508), 
          .S1(n105_adj_5507));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_26 (.A0(integrator4_adj_6023[59]), .B0(integrator3_adj_6022[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[60]), .B1(integrator3_adj_6022[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14446), .COUT(n14447), .S0(n114_adj_5510), 
          .S1(n111_adj_5509));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_24 (.A0(integrator4_adj_6023[57]), .B0(integrator3_adj_6022[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[58]), .B1(integrator3_adj_6022[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14445), .COUT(n14446), .S0(n120_adj_5512), 
          .S1(n117_adj_5511));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_22 (.A0(integrator4_adj_6023[55]), .B0(integrator3_adj_6022[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[56]), .B1(integrator3_adj_6022[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14444), .COUT(n14445), .S0(n126_adj_5514), 
          .S1(n123_adj_5513));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_20 (.A0(integrator4_adj_6023[53]), .B0(integrator3_adj_6022[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[54]), .B1(integrator3_adj_6022[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14443), .COUT(n14444), .S0(n132_adj_5516), 
          .S1(n129_adj_5515));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_18 (.A0(integrator4_adj_6023[51]), .B0(integrator3_adj_6022[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[52]), .B1(integrator3_adj_6022[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14442), .COUT(n14443), .S0(n138_adj_5518), 
          .S1(n135_adj_5517));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_16 (.A0(integrator4_adj_6023[49]), .B0(integrator3_adj_6022[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[50]), .B1(integrator3_adj_6022[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14441), .COUT(n14442), .S0(n144_adj_5520), 
          .S1(n141_adj_5519));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_14 (.A0(integrator4_adj_6023[47]), .B0(integrator3_adj_6022[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[48]), .B1(integrator3_adj_6022[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14440), .COUT(n14441), .S0(n150_adj_5522), 
          .S1(n147_adj_5521));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_12 (.A0(integrator4_adj_6023[45]), .B0(integrator3_adj_6022[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[46]), .B1(integrator3_adj_6022[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14439), .COUT(n14440), .S0(n156_adj_5524), 
          .S1(n153_adj_5523));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_10 (.A0(integrator4_adj_6023[43]), .B0(integrator3_adj_6022[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[44]), .B1(integrator3_adj_6022[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14438), .COUT(n14439), .S0(n162_adj_5526), 
          .S1(n159_adj_5525));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_8 (.A0(integrator4_adj_6023[41]), .B0(integrator3_adj_6022[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[42]), .B1(integrator3_adj_6022[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14437), .COUT(n14438), .S0(n168_adj_5528), 
          .S1(n165_adj_5527));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_6 (.A0(integrator4_adj_6023[39]), .B0(integrator3_adj_6022[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[40]), .B1(integrator3_adj_6022[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14436), .COUT(n14437), .S0(n174_adj_5530), 
          .S1(n171_adj_5529));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_4 (.A0(integrator4_adj_6023[37]), .B0(integrator3_adj_6022[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4_adj_6023[38]), .B1(integrator3_adj_6022[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14435), .COUT(n14436), .S0(n180_adj_5532), 
          .S1(n177_adj_5531));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1133_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1133_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator4_adj_6023[36]), .B1(integrator3_adj_6022[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14435), .S1(n183_adj_5533));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1133_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1133_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1133_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1133_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1055_add_4_15 (.A0(amdemod_d_11__N_1871[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14434), .S0(n32_adj_5534));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1055_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1055_add_4_15.INIT1 = 16'h0000;
    defparam _add_1_1055_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1055_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1055_add_4_13 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1871[9]), .D0(VCC_net), .A1(amdemod_d_11__N_1871[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n14433), .COUT(n14434), 
          .S0(n38_adj_5535));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1055_add_4_13.INIT0 = 16'h1e1e;
    defparam _add_1_1055_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1055_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1055_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1055_add_4_11 (.A0(n17134), .B0(amdemod_d_11__N_1871[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1871[8]), .B1(n17162), 
          .C1(n17279), .D1(n17146), .CIN(n14432), .COUT(n14433), .S0(n44_adj_5537), 
          .S1(n41_adj_5536));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1055_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_1055_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_1055_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1055_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1055_add_4_9 (.A0(n17132), .B0(amdemod_d_11__N_1871[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17133), .B1(amdemod_d_11__N_1871[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14431), .COUT(n14432), .S0(n50_adj_5539), 
          .S1(n47_adj_5538));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1055_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1055_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1055_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1055_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1055_add_4_7 (.A0(n17130), .B0(amdemod_d_11__N_1871[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17131), .B1(amdemod_d_11__N_1871[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14430), .COUT(n14431), .S0(n56_adj_5541), 
          .S1(n53_adj_5540));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1055_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1055_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1055_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1055_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1055_add_4_5 (.A0(n17128), .B0(amdemod_d_11__N_1871[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17129), .B1(amdemod_d_11__N_1871[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14429), .COUT(n14430), .S0(n62_adj_5543), 
          .S1(n59_adj_5542));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1055_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1055_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1055_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1055_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1055_add_4_3 (.A0(square_sum[3]), .B0(amdemod_d_11__N_1871[13]), 
          .C0(n17128), .D0(amdemod_d_11__N_1870[13]), .A1(n17127), .B1(amdemod_d_11__N_1871[0]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14428), .COUT(n14429), .S0(n68_adj_5545), 
          .S1(n65_adj_5544));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1055_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_1055_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1055_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1055_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1055_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14428), .S1(n71_adj_5546));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1055_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1055_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1055_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1055_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_15 (.A0(amdemod_d_11__N_2065), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14427), .S0(amdemod_d_11__N_1851[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1020_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1020_add_4_15.INIT1 = 16'h0000;
    defparam _add_1_1020_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_13 (.A0(amdemod_d_11__N_2071), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2068), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14426), .COUT(n14427), .S0(amdemod_d_11__N_1851[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1020_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1020_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1020_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_11 (.A0(amdemod_d_11__N_2077), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2074), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14425), .COUT(n14426), .S0(amdemod_d_11__N_1851[9]), 
          .S1(amdemod_d_11__N_1851[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1020_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1020_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1020_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_9 (.A0(amdemod_d_11__N_2083), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2080), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14424), .COUT(n14425), .S0(amdemod_d_11__N_1851[7]), 
          .S1(amdemod_d_11__N_1851[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1020_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1020_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1020_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_7 (.A0(amdemod_d_11__N_2089), .B0(n17162), .C0(n17279), 
          .D0(n17146), .A1(square_sum[23]), .B1(square_sum[22]), .C1(amdemod_d_11__N_2086), 
          .D1(VCC_net), .CIN(n14423), .COUT(n14424), .S0(amdemod_d_11__N_1851[5]), 
          .S1(amdemod_d_11__N_1851[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1020_add_4_7.INIT0 = 16'h596a;
    defparam _add_1_1020_add_4_7.INIT1 = 16'h1e1e;
    defparam _add_1_1020_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_5 (.A0(n17133), .B0(amdemod_d_11__N_2095), .C0(GND_net), 
          .D0(VCC_net), .A1(n17134), .B1(amdemod_d_11__N_2092), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14422), .COUT(n14423), .S0(amdemod_d_11__N_1851[3]), 
          .S1(amdemod_d_11__N_1851[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1020_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1020_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1020_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_3 (.A0(n17132), .B0(square_sum[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(n17132), .B1(amdemod_d_11__N_2098), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14421), .COUT(n14422), .S0(amdemod_d_11__N_1851[1]), 
          .S1(amdemod_d_11__N_1851[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1020_add_4_3.INIT0 = 16'h666a;
    defparam _add_1_1020_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1020_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1020_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14421), .S1(amdemod_d_11__N_1851[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1020_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1020_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1020_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1020_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_38 (.A0(integrator5_adj_6024[71]), .B0(integrator4_adj_6023[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14420), .S0(n78_adj_5547));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1136_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_36 (.A0(integrator5_adj_6024[69]), .B0(integrator4_adj_6023[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[70]), .B1(integrator4_adj_6023[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14419), .COUT(n14420), .S0(n84_adj_5549), 
          .S1(n81_adj_5548));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_34 (.A0(integrator5_adj_6024[67]), .B0(integrator4_adj_6023[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[68]), .B1(integrator4_adj_6023[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14418), .COUT(n14419), .S0(n90_adj_5551), 
          .S1(n87_adj_5550));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_32 (.A0(integrator5_adj_6024[65]), .B0(integrator4_adj_6023[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[66]), .B1(integrator4_adj_6023[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14417), .COUT(n14418), .S0(n96_adj_5553), 
          .S1(n93_adj_5552));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_30 (.A0(integrator5_adj_6024[63]), .B0(integrator4_adj_6023[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[64]), .B1(integrator4_adj_6023[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14416), .COUT(n14417), .S0(n102_adj_5555), 
          .S1(n99_adj_5554));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_28 (.A0(integrator5_adj_6024[61]), .B0(integrator4_adj_6023[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[62]), .B1(integrator4_adj_6023[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14415), .COUT(n14416), .S0(n108_adj_5557), 
          .S1(n105_adj_5556));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_26 (.A0(integrator5_adj_6024[59]), .B0(integrator4_adj_6023[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[60]), .B1(integrator4_adj_6023[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14414), .COUT(n14415), .S0(n114_adj_5559), 
          .S1(n111_adj_5558));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_24 (.A0(integrator5_adj_6024[57]), .B0(integrator4_adj_6023[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[58]), .B1(integrator4_adj_6023[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14413), .COUT(n14414), .S0(n120_adj_5561), 
          .S1(n117_adj_5560));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_22 (.A0(integrator5_adj_6024[55]), .B0(integrator4_adj_6023[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[56]), .B1(integrator4_adj_6023[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14412), .COUT(n14413), .S0(n126_adj_5563), 
          .S1(n123_adj_5562));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_20 (.A0(integrator5_adj_6024[53]), .B0(integrator4_adj_6023[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[54]), .B1(integrator4_adj_6023[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14411), .COUT(n14412), .S0(n132_adj_5565), 
          .S1(n129_adj_5564));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_18 (.A0(integrator5_adj_6024[51]), .B0(integrator4_adj_6023[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[52]), .B1(integrator4_adj_6023[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14410), .COUT(n14411), .S0(n138_adj_5567), 
          .S1(n135_adj_5566));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_16 (.A0(integrator5_adj_6024[49]), .B0(integrator4_adj_6023[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[50]), .B1(integrator4_adj_6023[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14409), .COUT(n14410), .S0(n144_adj_5569), 
          .S1(n141_adj_5568));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_14 (.A0(integrator5_adj_6024[47]), .B0(integrator4_adj_6023[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[48]), .B1(integrator4_adj_6023[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14408), .COUT(n14409), .S0(n150_adj_5571), 
          .S1(n147_adj_5570));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_12 (.A0(integrator5_adj_6024[45]), .B0(integrator4_adj_6023[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[46]), .B1(integrator4_adj_6023[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14407), .COUT(n14408), .S0(n156_adj_5573), 
          .S1(n153_adj_5572));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_10 (.A0(integrator5_adj_6024[43]), .B0(integrator4_adj_6023[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[44]), .B1(integrator4_adj_6023[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14406), .COUT(n14407), .S0(n162_adj_5575), 
          .S1(n159_adj_5574));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_8 (.A0(integrator5_adj_6024[41]), .B0(integrator4_adj_6023[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[42]), .B1(integrator4_adj_6023[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14405), .COUT(n14406), .S0(n168_adj_5577), 
          .S1(n165_adj_5576));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_6 (.A0(integrator5_adj_6024[39]), .B0(integrator4_adj_6023[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[40]), .B1(integrator4_adj_6023[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14404), .COUT(n14405), .S0(n174_adj_5579), 
          .S1(n171_adj_5578));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_4 (.A0(integrator5_adj_6024[37]), .B0(integrator4_adj_6023[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator5_adj_6024[38]), .B1(integrator4_adj_6023[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14403), .COUT(n14404), .S0(n180_adj_5581), 
          .S1(n177_adj_5580));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1136_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1136_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5_adj_6024[36]), .B1(integrator4_adj_6023[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14403), .S1(n183_adj_5582));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_1136_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1136_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1136_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1136_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_38 (.A0(comb_d9_adj_6032[71]), .B0(comb9_adj_6031[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14402), .S0(n78_adj_5583));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1139_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_36 (.A0(comb_d9_adj_6032[69]), .B0(comb9_adj_6031[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[70]), .B1(comb9_adj_6031[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14401), .COUT(n14402), .S0(n84_adj_5585), 
          .S1(n81_adj_5584));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_34 (.A0(comb_d9_adj_6032[67]), .B0(comb9_adj_6031[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[68]), .B1(comb9_adj_6031[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14400), .COUT(n14401), .S0(n90_adj_5587), 
          .S1(n87_adj_5586));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_32 (.A0(comb_d9_adj_6032[65]), .B0(comb9_adj_6031[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[66]), .B1(comb9_adj_6031[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14399), .COUT(n14400), .S0(n96_adj_5589), 
          .S1(n93_adj_5588));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_30 (.A0(comb_d9_adj_6032[63]), .B0(comb9_adj_6031[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[64]), .B1(comb9_adj_6031[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14398), .COUT(n14399), .S0(n102_adj_5591), 
          .S1(n99_adj_5590));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_28 (.A0(comb_d9_adj_6032[61]), .B0(comb9_adj_6031[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[62]), .B1(comb9_adj_6031[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14397), .COUT(n14398), .S0(n108_adj_5593), 
          .S1(n105_adj_5592));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_26 (.A0(comb_d9_adj_6032[59]), .B0(comb9_adj_6031[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[60]), .B1(comb9_adj_6031[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14396), .COUT(n14397), .S0(n114_adj_5595), 
          .S1(n111_adj_5594));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_24 (.A0(comb_d9_adj_6032[57]), .B0(comb9_adj_6031[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[58]), .B1(comb9_adj_6031[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14395), .COUT(n14396), .S0(n120_adj_5597), 
          .S1(n117_adj_5596));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_22 (.A0(comb_d9_adj_6032[55]), .B0(comb9_adj_6031[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[56]), .B1(comb9_adj_6031[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14394), .COUT(n14395));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_20 (.A0(comb_d9_adj_6032[53]), .B0(comb9_adj_6031[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[54]), .B1(comb9_adj_6031[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14393), .COUT(n14394));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_18 (.A0(comb_d9_adj_6032[51]), .B0(comb9_adj_6031[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[52]), .B1(comb9_adj_6031[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14392), .COUT(n14393));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_16 (.A0(comb_d9_adj_6032[49]), .B0(comb9_adj_6031[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[50]), .B1(comb9_adj_6031[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14391), .COUT(n14392));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_14 (.A0(comb_d9_adj_6032[47]), .B0(comb9_adj_6031[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[48]), .B1(comb9_adj_6031[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14390), .COUT(n14391));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_12 (.A0(comb_d9_adj_6032[45]), .B0(comb9_adj_6031[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[46]), .B1(comb9_adj_6031[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14389), .COUT(n14390));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_10 (.A0(comb_d9_adj_6032[43]), .B0(comb9_adj_6031[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[44]), .B1(comb9_adj_6031[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14388), .COUT(n14389));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_8 (.A0(comb_d9_adj_6032[41]), .B0(comb9_adj_6031[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[42]), .B1(comb9_adj_6031[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14387), .COUT(n14388));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_6 (.A0(comb_d9_adj_6032[39]), .B0(comb9_adj_6031[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[40]), .B1(comb9_adj_6031[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14386), .COUT(n14387));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_4 (.A0(comb_d9_adj_6032[37]), .B0(comb9_adj_6031[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[38]), .B1(comb9_adj_6031[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14385), .COUT(n14386));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1139_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1139_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9_adj_6032[36]), .B1(comb9_adj_6031[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14385));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1139_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1139_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1139_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1139_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_38 (.A0(comb_d6[71]), .B0(comb6[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14384), .S0(n78_adj_5389));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1208_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_36 (.A0(comb_d6[69]), .B0(comb6[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[70]), .B1(comb6[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14383), .COUT(n14384), .S0(n84_adj_5391), 
          .S1(n81_adj_5390));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_34 (.A0(comb_d6[67]), .B0(comb6[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[68]), .B1(comb6[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14382), .COUT(n14383), .S0(n90_adj_5393), 
          .S1(n87_adj_5392));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_32 (.A0(comb_d6[65]), .B0(comb6[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[66]), .B1(comb6[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14381), .COUT(n14382), .S0(n96_adj_5395), 
          .S1(n93_adj_5394));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_30 (.A0(comb_d6[63]), .B0(comb6[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[64]), .B1(comb6[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14380), .COUT(n14381), .S0(n102_adj_5397), 
          .S1(n99_adj_5396));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_28 (.A0(comb_d6[61]), .B0(comb6[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[62]), .B1(comb6[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14379), .COUT(n14380), .S0(n108_adj_5399), 
          .S1(n105_adj_5398));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_26 (.A0(comb_d6[59]), .B0(comb6[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[60]), .B1(comb6[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14378), .COUT(n14379), .S0(n114_adj_5401), 
          .S1(n111_adj_5400));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_24 (.A0(comb_d6[57]), .B0(comb6[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[58]), .B1(comb6[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14377), .COUT(n14378), .S0(n120_adj_5403), 
          .S1(n117_adj_5402));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_22 (.A0(comb_d6[55]), .B0(comb6[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[56]), .B1(comb6[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14376), .COUT(n14377), .S0(n126_adj_5405), 
          .S1(n123_adj_5404));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_20 (.A0(comb_d6[53]), .B0(comb6[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[54]), .B1(comb6[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14375), .COUT(n14376), .S0(n132_adj_5407), 
          .S1(n129_adj_5406));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_18 (.A0(comb_d6[51]), .B0(comb6[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[52]), .B1(comb6[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14374), .COUT(n14375), .S0(n138_adj_5409), 
          .S1(n135_adj_5408));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_16 (.A0(comb_d6[49]), .B0(comb6[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[50]), .B1(comb6[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14373), .COUT(n14374), .S0(n144_adj_5411), 
          .S1(n141_adj_5410));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_14 (.A0(comb_d6[47]), .B0(comb6[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[48]), .B1(comb6[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14372), .COUT(n14373), .S0(n150_adj_5413), 
          .S1(n147_adj_5412));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_12 (.A0(comb_d6[45]), .B0(comb6[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[46]), .B1(comb6[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14371), .COUT(n14372), .S0(n156_adj_5415), 
          .S1(n153_adj_5414));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_10 (.A0(comb_d6[43]), .B0(comb6[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[44]), .B1(comb6[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14370), .COUT(n14371), .S0(n162_adj_5417), 
          .S1(n159_adj_5416));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_8 (.A0(comb_d6[41]), .B0(comb6[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[42]), .B1(comb6[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14369), .COUT(n14370), .S0(n168_adj_5419), 
          .S1(n165_adj_5418));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_6 (.A0(comb_d6[39]), .B0(comb6[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[40]), .B1(comb6[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14368), .COUT(n14369), .S0(n174_adj_5421), 
          .S1(n171_adj_5420));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_4 (.A0(comb_d6[37]), .B0(comb6[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[38]), .B1(comb6[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14367), .COUT(n14368), .S0(n180_adj_5423), 
          .S1(n177_adj_5422));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1208_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_4.INJECT1_1 = "NO";
    FD1S3AX phase_accum_e3_i0_i1 (.D(n318), .CK(clk_80mhz), .Q(phase_accum[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i1.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i2 (.D(n315), .CK(clk_80mhz), .Q(phase_accum[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i2.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i3 (.D(n312), .CK(clk_80mhz), .Q(phase_accum[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i3.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i4 (.D(n309), .CK(clk_80mhz), .Q(phase_accum[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i4.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i5 (.D(n306), .CK(clk_80mhz), .Q(phase_accum[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i5.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i6 (.D(n303), .CK(clk_80mhz), .Q(phase_accum[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i6.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i7 (.D(n300), .CK(clk_80mhz), .Q(phase_accum[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i7.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i8 (.D(n297), .CK(clk_80mhz), .Q(phase_accum[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i8.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i9 (.D(n294), .CK(clk_80mhz), .Q(phase_accum[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i9.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i10 (.D(n291), .CK(clk_80mhz), .Q(phase_accum[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i10.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i11 (.D(n288), .CK(clk_80mhz), .Q(phase_accum[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i11.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i12 (.D(n285), .CK(clk_80mhz), .Q(phase_accum[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i12.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i13 (.D(n282), .CK(clk_80mhz), .Q(phase_accum[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i13.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i14 (.D(n279), .CK(clk_80mhz), .Q(phase_accum[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i14.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i15 (.D(n276), .CK(clk_80mhz), .Q(phase_accum[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i15.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i16 (.D(n273), .CK(clk_80mhz), .Q(phase_accum[16]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i16.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i17 (.D(n270), .CK(clk_80mhz), .Q(phase_accum[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i17.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i18 (.D(n267), .CK(clk_80mhz), .Q(phase_accum[18]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i18.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i19 (.D(n264), .CK(clk_80mhz), .Q(phase_accum[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i19.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i20 (.D(n261), .CK(clk_80mhz), .Q(phase_accum[20]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i20.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i21 (.D(n258), .CK(clk_80mhz), .Q(phase_accum[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i21.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i22 (.D(n255), .CK(clk_80mhz), .Q(phase_accum[22]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i22.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i23 (.D(n252), .CK(clk_80mhz), .Q(phase_accum[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i23.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i24 (.D(n249), .CK(clk_80mhz), .Q(phase_accum[24]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i24.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i25 (.D(n246), .CK(clk_80mhz), .Q(phase_accum[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i25.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i26 (.D(n243), .CK(clk_80mhz), .Q(phase_accum[26]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i26.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i27 (.D(n240), .CK(clk_80mhz), .Q(phase_accum[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i27.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i28 (.D(n237), .CK(clk_80mhz), .Q(phase_accum[28]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i28.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i29 (.D(n234), .CK(clk_80mhz), .Q(phase_accum[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i29.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i30 (.D(n231), .CK(clk_80mhz), .Q(phase_accum[30]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i30.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i31 (.D(n228), .CK(clk_80mhz), .Q(phase_accum[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i31.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i32 (.D(n225), .CK(clk_80mhz), .Q(phase_accum[32]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i32.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i33 (.D(n222), .CK(clk_80mhz), .Q(phase_accum[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i33.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i34 (.D(n219), .CK(clk_80mhz), .Q(phase_accum[34]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i34.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i35 (.D(n216), .CK(clk_80mhz), .Q(phase_accum[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i35.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i36 (.D(n213), .CK(clk_80mhz), .Q(phase_accum[36]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i36.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i37 (.D(n210), .CK(clk_80mhz), .Q(phase_accum[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i37.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i38 (.D(n207), .CK(clk_80mhz), .Q(phase_accum[38]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i38.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i39 (.D(n204), .CK(clk_80mhz), .Q(phase_accum[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i39.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i40 (.D(n201), .CK(clk_80mhz), .Q(phase_accum[40]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i40.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i41 (.D(n198), .CK(clk_80mhz), .Q(phase_accum[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i41.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i42 (.D(n195), .CK(clk_80mhz), .Q(phase_accum[42]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i42.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i43 (.D(n192), .CK(clk_80mhz), .Q(phase_accum[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i43.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i44 (.D(n189), .CK(clk_80mhz), .Q(phase_accum[44]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i44.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i45 (.D(n186), .CK(clk_80mhz), .Q(phase_accum[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i45.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i46 (.D(n183_adj_5677), .CK(clk_80mhz), .Q(phase_accum[46]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i46.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i47 (.D(n180_adj_5676), .CK(clk_80mhz), .Q(phase_accum[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i47.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i48 (.D(n177_adj_5675), .CK(clk_80mhz), .Q(phase_accum[48]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i48.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i49 (.D(n174_adj_5674), .CK(clk_80mhz), .Q(phase_accum[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i49.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i50 (.D(n171_adj_5673), .CK(clk_80mhz), .Q(phase_accum[50]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i50.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i51 (.D(n168_adj_5672), .CK(clk_80mhz), .Q(phase_accum[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i51.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i52 (.D(n165_adj_5671), .CK(clk_80mhz), .Q(phase_accum[52]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i52.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i53 (.D(n162_adj_5670), .CK(clk_80mhz), .Q(phase_accum[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i53.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i54 (.D(n159_adj_5669), .CK(clk_80mhz), .Q(phase_accum[54]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i54.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i55 (.D(n156_adj_5668), .CK(clk_80mhz), .Q(phase_accum[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i55.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i56 (.D(n153_adj_5667), .CK(clk_80mhz), .Q(phase_acc[56]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i56.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i57 (.D(n150_adj_5666), .CK(clk_80mhz), .Q(phase_acc[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i57.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i58 (.D(n147_adj_5665), .CK(clk_80mhz), .Q(phase_acc[58]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i58.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i59 (.D(n144_adj_5664), .CK(clk_80mhz), .Q(phase_acc[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i59.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i60 (.D(n141_adj_5663), .CK(clk_80mhz), .Q(phase_acc[60]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i60.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i61 (.D(n138_adj_5662), .CK(clk_80mhz), .Q(phase_acc[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i61.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i62 (.D(n135_adj_5661), .CK(clk_80mhz), .Q(phase_acc[62]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i62.GSR = "ENABLED";
    FD1S3AX phase_accum_e3_i0_i63 (.D(n132_adj_5660), .CK(clk_80mhz), .Q(phase_acc[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_e3_i0_i63.GSR = "ENABLED";
    CCU2C _add_1_1244_add_4_37 (.A0(phase_inc_gen[36]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[37]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15693), .COUT(n15694), .S0(n211_adj_5931), 
          .S1(n208_adj_5930));
    defparam _add_1_1244_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_35 (.A0(phase_inc_gen[34]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[35]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15692), .COUT(n15693), .S0(n217_adj_5933), 
          .S1(n214_adj_5932));
    defparam _add_1_1244_add_4_35.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_33 (.A0(phase_inc_gen[32]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[33]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15691), .COUT(n15692), .S0(n223_adj_5935), 
          .S1(n220_adj_5934));
    defparam _add_1_1244_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_31 (.A0(phase_inc_gen[30]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[31]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15690), .COUT(n15691), .S0(n229_adj_5937), 
          .S1(n226_adj_5936));
    defparam _add_1_1244_add_4_31.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_29 (.A0(phase_inc_gen[28]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[29]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15689), .COUT(n15690), .S0(n235_adj_5939), 
          .S1(n232_adj_5938));
    defparam _add_1_1244_add_4_29.INIT0 = 16'haaa0;
    defparam _add_1_1244_add_4_29.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_27 (.A0(phase_inc_gen[26]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[27]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15688), .COUT(n15689), .S0(n241_adj_5941), 
          .S1(n238_adj_5940));
    defparam _add_1_1244_add_4_27.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_25 (.A0(phase_inc_gen[24]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[25]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15687), .COUT(n15688), .S0(n247_adj_5943), 
          .S1(n244_adj_5942));
    defparam _add_1_1244_add_4_25.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_25.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_23 (.A0(phase_inc_gen[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[23]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15686), .COUT(n15687), .S0(n253_adj_5945), 
          .S1(n250_adj_5944));
    defparam _add_1_1244_add_4_23.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_23.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_21 (.A0(phase_inc_gen[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[21]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15685), .COUT(n15686), .S0(n259_adj_5947), 
          .S1(n256_adj_5946));
    defparam _add_1_1244_add_4_21.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_21.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_19 (.A0(phase_inc_gen[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15684), .COUT(n15685), .S0(n265_adj_5949), 
          .S1(n262_adj_5948));
    defparam _add_1_1244_add_4_19.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_16 (.A0(integrator4[49]), .B0(integrator3[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[50]), .B1(integrator3[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15266), .COUT(n15267), .S0(n144_adj_5111), 
          .S1(n141_adj_5110));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1208_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[36]), .B1(comb6[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14367), .S1(n183_adj_5424));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1208_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1208_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1208_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1208_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1214_add_4_10 (.A0(n17162), .B0(n17279), .C0(GND_net), 
          .D0(VCC_net), .A1(n17162), .B1(n17279), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14365), .S0(n27_adj_5462), .S1(n24_adj_5461));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1214_add_4_10.INIT0 = 16'h8887;
    defparam _add_1_1214_add_4_10.INIT1 = 16'h8887;
    defparam _add_1_1214_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1214_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1214_add_4_8 (.A0(n17157), .B0(n6_adj_4757), .C0(GND_net), 
          .D0(VCC_net), .A1(n17162), .B1(n17279), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14364), .COUT(n14365), .S0(n33_adj_5464), .S1(n30_adj_5463));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1214_add_4_8.INIT0 = 16'h9996;
    defparam _add_1_1214_add_4_8.INIT1 = 16'h9996;
    defparam _add_1_1214_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1214_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1214_add_4_6 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1830[1]), .D0(VCC_net), .A1(n17162), .B1(n4_adj_2948), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14363), .COUT(n14364), .S0(n39_adj_5466), 
          .S1(n36_adj_5465));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1214_add_4_6.INIT0 = 16'he1e1;
    defparam _add_1_1214_add_4_6.INIT1 = 16'h9996;
    defparam _add_1_1214_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1214_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1214_add_4_4 (.A0(square_sum[19]), .B0(n17162), .C0(n17279), 
          .D0(n17146), .A1(n17137), .B1(square_sum[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14362), .COUT(n14363), .S0(n45_adj_5468), 
          .S1(n42_adj_5467));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1214_add_4_4.INIT0 = 16'h596a;
    defparam _add_1_1214_add_4_4.INIT1 = 16'h6665;
    defparam _add_1_1214_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1214_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1214_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[18]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14362), .S1(n48_adj_5469));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1214_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1214_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1214_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1214_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_37 (.A0(integrator3[70]), .B0(cout_adj_5074), 
          .C0(n81_adj_5090), .D0(integrator4[70]), .A1(integrator3[71]), 
          .B1(cout_adj_5074), .C1(n78_adj_5089), .D1(integrator4[71]), 
          .CIN(n14360), .S0(integrator4_71__N_634[70]), .S1(integrator4_71__N_634[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_35 (.A0(integrator3[68]), .B0(cout_adj_5074), 
          .C0(n87_adj_5092), .D0(integrator4[68]), .A1(integrator3[69]), 
          .B1(cout_adj_5074), .C1(n84_adj_5091), .D1(integrator4[69]), 
          .CIN(n14359), .COUT(n14360), .S0(integrator4_71__N_634[68]), 
          .S1(integrator4_71__N_634[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_33 (.A0(integrator3[66]), .B0(cout_adj_5074), 
          .C0(n93_adj_5094), .D0(integrator4[66]), .A1(integrator3[67]), 
          .B1(cout_adj_5074), .C1(n90_adj_5093), .D1(integrator4[67]), 
          .CIN(n14358), .COUT(n14359), .S0(integrator4_71__N_634[66]), 
          .S1(integrator4_71__N_634[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_31 (.A0(integrator3[64]), .B0(cout_adj_5074), 
          .C0(n99_adj_5096), .D0(integrator4[64]), .A1(integrator3[65]), 
          .B1(cout_adj_5074), .C1(n96_adj_5095), .D1(integrator4[65]), 
          .CIN(n14357), .COUT(n14358), .S0(integrator4_71__N_634[64]), 
          .S1(integrator4_71__N_634[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_29 (.A0(integrator3[62]), .B0(cout_adj_5074), 
          .C0(n105_adj_5098), .D0(integrator4[62]), .A1(integrator3[63]), 
          .B1(cout_adj_5074), .C1(n102_adj_5097), .D1(integrator4[63]), 
          .CIN(n14356), .COUT(n14357), .S0(integrator4_71__N_634[62]), 
          .S1(integrator4_71__N_634[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_27 (.A0(integrator3[60]), .B0(cout_adj_5074), 
          .C0(n111_adj_5100), .D0(integrator4[60]), .A1(integrator3[61]), 
          .B1(cout_adj_5074), .C1(n108_adj_5099), .D1(integrator4[61]), 
          .CIN(n14355), .COUT(n14356), .S0(integrator4_71__N_634[60]), 
          .S1(integrator4_71__N_634[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_25 (.A0(integrator3[58]), .B0(cout_adj_5074), 
          .C0(n117_adj_5102), .D0(integrator4[58]), .A1(integrator3[59]), 
          .B1(cout_adj_5074), .C1(n114_adj_5101), .D1(integrator4[59]), 
          .CIN(n14354), .COUT(n14355), .S0(integrator4_71__N_634[58]), 
          .S1(integrator4_71__N_634[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_23 (.A0(integrator3[56]), .B0(cout_adj_5074), 
          .C0(n123_adj_5104), .D0(integrator4[56]), .A1(integrator3[57]), 
          .B1(cout_adj_5074), .C1(n120_adj_5103), .D1(integrator4[57]), 
          .CIN(n14353), .COUT(n14354), .S0(integrator4_71__N_634[56]), 
          .S1(integrator4_71__N_634[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_21 (.A0(integrator3[54]), .B0(cout_adj_5074), 
          .C0(n129_adj_5106), .D0(integrator4[54]), .A1(integrator3[55]), 
          .B1(cout_adj_5074), .C1(n126_adj_5105), .D1(integrator4[55]), 
          .CIN(n14352), .COUT(n14353), .S0(integrator4_71__N_634[54]), 
          .S1(integrator4_71__N_634[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_19 (.A0(integrator3[52]), .B0(cout_adj_5074), 
          .C0(n135_adj_5108), .D0(integrator4[52]), .A1(integrator3[53]), 
          .B1(cout_adj_5074), .C1(n132_adj_5107), .D1(integrator4[53]), 
          .CIN(n14351), .COUT(n14352), .S0(integrator4_71__N_634[52]), 
          .S1(integrator4_71__N_634[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_17 (.A0(integrator3[50]), .B0(cout_adj_5074), 
          .C0(n141_adj_5110), .D0(integrator4[50]), .A1(integrator3[51]), 
          .B1(cout_adj_5074), .C1(n138_adj_5109), .D1(integrator4[51]), 
          .CIN(n14350), .COUT(n14351), .S0(integrator4_71__N_634[50]), 
          .S1(integrator4_71__N_634[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_15 (.A0(integrator3[48]), .B0(cout_adj_5074), 
          .C0(n147_adj_5112), .D0(integrator4[48]), .A1(integrator3[49]), 
          .B1(cout_adj_5074), .C1(n144_adj_5111), .D1(integrator4[49]), 
          .CIN(n14349), .COUT(n14350), .S0(integrator4_71__N_634[48]), 
          .S1(integrator4_71__N_634[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_13 (.A0(integrator3[46]), .B0(cout_adj_5074), 
          .C0(n153_adj_5114), .D0(integrator4[46]), .A1(integrator3[47]), 
          .B1(cout_adj_5074), .C1(n150_adj_5113), .D1(integrator4[47]), 
          .CIN(n14348), .COUT(n14349), .S0(integrator4_71__N_634[46]), 
          .S1(integrator4_71__N_634[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_11 (.A0(integrator3[44]), .B0(cout_adj_5074), 
          .C0(n159_adj_5116), .D0(integrator4[44]), .A1(integrator3[45]), 
          .B1(cout_adj_5074), .C1(n156_adj_5115), .D1(integrator4[45]), 
          .CIN(n14347), .COUT(n14348), .S0(integrator4_71__N_634[44]), 
          .S1(integrator4_71__N_634[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_9 (.A0(integrator3[42]), .B0(cout_adj_5074), 
          .C0(n165_adj_5118), .D0(integrator4[42]), .A1(integrator3[43]), 
          .B1(cout_adj_5074), .C1(n162_adj_5117), .D1(integrator4[43]), 
          .CIN(n14346), .COUT(n14347), .S0(integrator4_71__N_634[42]), 
          .S1(integrator4_71__N_634[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_7 (.A0(integrator3[40]), .B0(cout_adj_5074), 
          .C0(n171_adj_5120), .D0(integrator4[40]), .A1(integrator3[41]), 
          .B1(cout_adj_5074), .C1(n168_adj_5119), .D1(integrator4[41]), 
          .CIN(n14345), .COUT(n14346), .S0(integrator4_71__N_634[40]), 
          .S1(integrator4_71__N_634[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_5 (.A0(integrator3[38]), .B0(cout_adj_5074), 
          .C0(n177_adj_5122), .D0(integrator4[38]), .A1(integrator3[39]), 
          .B1(cout_adj_5074), .C1(n174_adj_5121), .D1(integrator4[39]), 
          .CIN(n14344), .COUT(n14345), .S0(integrator4_71__N_634[38]), 
          .S1(integrator4_71__N_634[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_3 (.A0(integrator3[36]), .B0(cout_adj_5074), 
          .C0(n183_adj_5124), .D0(integrator4[36]), .A1(integrator3[37]), 
          .B1(cout_adj_5074), .C1(n180_adj_5123), .D1(integrator4[37]), 
          .CIN(n14343), .COUT(n14344), .S0(integrator4_71__N_634[36]), 
          .S1(integrator4_71__N_634[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1046_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1046_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1046_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5074), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14343));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1046_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1046_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1046_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1046_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1217_add_4_16 (.A0(amdemod_d_11__N_1870[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14339), .S0(n34_adj_5470));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1217_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1217_add_4_16.INIT1 = 16'h0000;
    defparam _add_1_1217_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1217_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1217_add_4_14 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1870[9]), .D0(VCC_net), .A1(amdemod_d_11__N_1870[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n14338), .COUT(n14339), 
          .S0(n40_adj_5471));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1217_add_4_14.INIT0 = 16'he1e1;
    defparam _add_1_1217_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_1217_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1217_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1217_add_4_12 (.A0(n17134), .B0(amdemod_d_11__N_1870[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17137), .B1(amdemod_d_11__N_1870[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14337), .COUT(n14338), .S0(n46_adj_5473), 
          .S1(n43_adj_5472));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1217_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1217_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1217_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1217_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1217_add_4_10 (.A0(n17132), .B0(amdemod_d_11__N_1870[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1870[6]), .B1(amdemod_d_11__N_1841[11]), 
          .C1(n17134), .D1(amdemod_d_11__N_1840[11]), .CIN(n14336), .COUT(n14337), 
          .S0(n52_adj_5475), .S1(n49_adj_5474));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1217_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1217_add_4_10.INIT1 = 16'h656a;
    defparam _add_1_1217_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1217_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1217_add_4_8 (.A0(n17130), .B0(amdemod_d_11__N_1870[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1870[4]), .B1(amdemod_d_11__N_1851[13]), 
          .C1(n17132), .D1(amdemod_d_11__N_1850[13]), .CIN(n14335), .COUT(n14336), 
          .S0(n58_adj_5477), .S1(n55_adj_5476));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1217_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1217_add_4_8.INIT1 = 16'h656a;
    defparam _add_1_1217_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1217_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1217_add_4_6 (.A0(n17128), .B0(amdemod_d_11__N_1870[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1870[2]), .B1(amdemod_d_11__N_1861[13]), 
          .C1(n17130), .D1(amdemod_d_11__N_1860[13]), .CIN(n14334), .COUT(n14335), 
          .S0(n64_adj_5479), .S1(n61_adj_5478));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1217_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1217_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_1217_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1217_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1217_add_4_4 (.A0(n17127), .B0(square_sum[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_d_11__N_1870[0]), .B1(amdemod_d_11__N_1871[13]), 
          .C1(n17128), .D1(amdemod_d_11__N_1870[13]), .CIN(n14333), .COUT(n14334), 
          .S0(n70_adj_5481), .S1(n67_adj_5480));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1217_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1217_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_1217_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1217_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1217_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14333), .S1(n73_adj_5482));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1217_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1217_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1217_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1217_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_978_add_4_15 (.A0(amdemod_d_11__N_1840[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14332), .S0(n32_adj_5059));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_978_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_978_add_4_15.INIT1 = 16'h0000;
    defparam _add_1_978_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_978_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_978_add_4_13 (.A0(amdemod_d_11__N_1840[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1840[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14331), .COUT(n14332), .S0(n38_adj_5060));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_978_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_978_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_978_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_978_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_978_add_4_11 (.A0(amdemod_d_11__N_1840[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1840[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14330), .COUT(n14331), .S0(n44_adj_5062), 
          .S1(n41_adj_5061));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_978_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_978_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_978_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_978_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_978_add_4_9 (.A0(amdemod_d_11__N_1840[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1840[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14329), .COUT(n14330), .S0(n50_adj_5064), 
          .S1(n47_adj_5063));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_978_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_978_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_978_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_978_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_978_add_4_7 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1840[3]), .D0(VCC_net), .A1(amdemod_d_11__N_1840[4]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n14328), .COUT(n14329), 
          .S0(n56_adj_5066), .S1(n53_adj_5065));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_978_add_4_7.INIT0 = 16'h1e1e;
    defparam _add_1_978_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_978_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_978_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_978_add_4_5 (.A0(n17134), .B0(amdemod_d_11__N_1840[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1840[2]), .B1(n17162), 
          .C1(n17279), .D1(n17146), .CIN(n14327), .COUT(n14328), .S0(n62_adj_5068), 
          .S1(n59_adj_5067));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_978_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_978_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_978_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_978_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_978_add_4_3 (.A0(square_sum[15]), .B0(amdemod_d_11__N_1841[11]), 
          .C0(n17134), .D0(amdemod_d_11__N_1840[11]), .A1(n17133), .B1(amdemod_d_11__N_1840[0]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14326), .COUT(n14327), .S0(n68_adj_5070), 
          .S1(n65_adj_5069));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_978_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_978_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_978_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_978_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_978_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14326), .S1(n71_adj_5071));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_978_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_978_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_978_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_978_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_38 (.A0(integrator_d_tmp_adj_6019[71]), .B0(integrator_tmp_adj_6018[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14325), .S0(n78_adj_5799));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1151_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_36 (.A0(integrator_d_tmp_adj_6019[69]), .B0(integrator_tmp_adj_6018[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[70]), 
          .B1(integrator_tmp_adj_6018[70]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14324), .COUT(n14325), .S0(n84_adj_5801), .S1(n81_adj_5800));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_34 (.A0(integrator_d_tmp_adj_6019[67]), .B0(integrator_tmp_adj_6018[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[68]), 
          .B1(integrator_tmp_adj_6018[68]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14323), .COUT(n14324), .S0(n90_adj_5803), .S1(n87_adj_5802));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_32 (.A0(integrator_d_tmp_adj_6019[65]), .B0(integrator_tmp_adj_6018[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[66]), 
          .B1(integrator_tmp_adj_6018[66]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14322), .COUT(n14323), .S0(n96_adj_5805), .S1(n93_adj_5804));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_30 (.A0(integrator_d_tmp_adj_6019[63]), .B0(integrator_tmp_adj_6018[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[64]), 
          .B1(integrator_tmp_adj_6018[64]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14321), .COUT(n14322), .S0(n102_adj_5807), .S1(n99_adj_5806));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_28 (.A0(integrator_d_tmp_adj_6019[61]), .B0(integrator_tmp_adj_6018[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[62]), 
          .B1(integrator_tmp_adj_6018[62]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14320), .COUT(n14321), .S0(n108_adj_5809), .S1(n105_adj_5808));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_26 (.A0(integrator_d_tmp_adj_6019[59]), .B0(integrator_tmp_adj_6018[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[60]), 
          .B1(integrator_tmp_adj_6018[60]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14319), .COUT(n14320), .S0(n114_adj_5811), .S1(n111_adj_5810));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_24 (.A0(integrator_d_tmp_adj_6019[57]), .B0(integrator_tmp_adj_6018[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[58]), 
          .B1(integrator_tmp_adj_6018[58]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14318), .COUT(n14319), .S0(n120_adj_5813), .S1(n117_adj_5812));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_22 (.A0(integrator_d_tmp_adj_6019[55]), .B0(integrator_tmp_adj_6018[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[56]), 
          .B1(integrator_tmp_adj_6018[56]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14317), .COUT(n14318), .S0(n126_adj_5815), .S1(n123_adj_5814));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_20 (.A0(integrator_d_tmp_adj_6019[53]), .B0(integrator_tmp_adj_6018[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[54]), 
          .B1(integrator_tmp_adj_6018[54]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14316), .COUT(n14317), .S0(n132_adj_5817), .S1(n129_adj_5816));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_18 (.A0(integrator_d_tmp_adj_6019[51]), .B0(integrator_tmp_adj_6018[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[52]), 
          .B1(integrator_tmp_adj_6018[52]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14315), .COUT(n14316), .S0(n138_adj_5819), .S1(n135_adj_5818));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_16 (.A0(integrator_d_tmp_adj_6019[49]), .B0(integrator_tmp_adj_6018[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[50]), 
          .B1(integrator_tmp_adj_6018[50]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14314), .COUT(n14315), .S0(n144_adj_5821), .S1(n141_adj_5820));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_14 (.A0(integrator_d_tmp_adj_6019[47]), .B0(integrator_tmp_adj_6018[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[48]), 
          .B1(integrator_tmp_adj_6018[48]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14313), .COUT(n14314), .S0(n150_adj_5823), .S1(n147_adj_5822));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_12 (.A0(integrator_d_tmp_adj_6019[45]), .B0(integrator_tmp_adj_6018[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[46]), 
          .B1(integrator_tmp_adj_6018[46]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14312), .COUT(n14313), .S0(n156_adj_5825), .S1(n153_adj_5824));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_10 (.A0(integrator_d_tmp_adj_6019[43]), .B0(integrator_tmp_adj_6018[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[44]), 
          .B1(integrator_tmp_adj_6018[44]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14311), .COUT(n14312), .S0(n162_adj_5827), .S1(n159_adj_5826));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_8 (.A0(integrator_d_tmp_adj_6019[41]), .B0(integrator_tmp_adj_6018[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[42]), 
          .B1(integrator_tmp_adj_6018[42]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14310), .COUT(n14311), .S0(n168_adj_5829), .S1(n165_adj_5828));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_6 (.A0(integrator_d_tmp_adj_6019[39]), .B0(integrator_tmp_adj_6018[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[40]), 
          .B1(integrator_tmp_adj_6018[40]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14309), .COUT(n14310), .S0(n174_adj_5831), .S1(n171_adj_5830));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_4 (.A0(integrator_d_tmp_adj_6019[37]), .B0(integrator_tmp_adj_6018[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[38]), 
          .B1(integrator_tmp_adj_6018[38]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14308), .COUT(n14309), .S0(n180_adj_5833), .S1(n177_adj_5832));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1151_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1151_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator_d_tmp_adj_6019[36]), .B1(integrator_tmp_adj_6018[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n14308), .S1(n183_adj_5834));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1151_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1151_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1151_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1151_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1058_add_4_15 (.A0(amdemod_d_11__N_1870[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14307), .S0(n32_adj_5598));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1058_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1058_add_4_15.INIT1 = 16'h0000;
    defparam _add_1_1058_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1058_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1058_add_4_13 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1870[9]), .D0(VCC_net), .A1(amdemod_d_11__N_1870[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n14306), .COUT(n14307), 
          .S0(n38_adj_5599));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1058_add_4_13.INIT0 = 16'h1e1e;
    defparam _add_1_1058_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1058_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1058_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1058_add_4_11 (.A0(n17134), .B0(amdemod_d_11__N_1870[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1870[8]), .B1(n17162), 
          .C1(n17279), .D1(n17146), .CIN(n14305), .COUT(n14306), .S0(n44_adj_5601), 
          .S1(n41_adj_5600));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1058_add_4_11.INIT0 = 16'h9995;
    defparam _add_1_1058_add_4_11.INIT1 = 16'h596a;
    defparam _add_1_1058_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1058_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1058_add_4_9 (.A0(n17132), .B0(amdemod_d_11__N_1870[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17133), .B1(amdemod_d_11__N_1870[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14304), .COUT(n14305), .S0(n50_adj_5603), 
          .S1(n47_adj_5602));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1058_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1058_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1058_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1058_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1058_add_4_7 (.A0(n17130), .B0(amdemod_d_11__N_1870[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17131), .B1(amdemod_d_11__N_1870[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14303), .COUT(n14304), .S0(n56_adj_5605), 
          .S1(n53_adj_5604));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1058_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1058_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1058_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1058_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1058_add_4_5 (.A0(n17128), .B0(amdemod_d_11__N_1870[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17129), .B1(amdemod_d_11__N_1870[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14302), .COUT(n14303), .S0(n62_adj_5607), 
          .S1(n59_adj_5606));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1058_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1058_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1058_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1058_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1058_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14301), .S1(n71_adj_5610));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1058_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1058_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1058_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1058_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1058_add_4_3 (.A0(square_sum[3]), .B0(amdemod_d_11__N_1871[13]), 
          .C0(n17128), .D0(amdemod_d_11__N_1870[13]), .A1(n17127), .B1(amdemod_d_11__N_1870[0]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14301), .COUT(n14302), .S0(n68_adj_5609), 
          .S1(n65_adj_5608));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1058_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_1058_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1058_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1058_add_4_3.INJECT1_1 = "NO";
    FD1P3AX cic_gain__i2 (.D(led_c_1), .SP(clk_80mhz_enable_1445), .CK(clk_80mhz), 
            .Q(cic_gain[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam cic_gain__i2.GSR = "ENABLED";
    LUT4 mux_251_i61_4_lut (.A(n11397), .B(n139_adj_5907), .C(n17136), 
         .D(n2244), .Z(n1984)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i61_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1244_add_4_17 (.A0(phase_inc_gen[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15683), .COUT(n15684), .S0(n271_adj_5951), 
          .S1(n268_adj_5950));
    defparam _add_1_1244_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1244_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_17.INJECT1_1 = "NO";
    LUT4 i1886_4_lut (.A(n136_adj_5906), .B(n130), .C(led_c_3), .D(n17144), 
         .Z(n11620)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1886_4_lut.init = 16'hcac0;
    LUT4 i27_3_lut_3_lut (.A(led_c_3), .B(n17150), .C(n247), .Z(n13_adj_4747)) /* synthesis lut_function=(!(A (C)+!A !(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i27_3_lut_3_lut.init = 16'h4e4e;
    CCU2C _add_1_1244_add_4_15 (.A0(phase_inc_gen[14]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15682), .COUT(n15683), .S0(n277_adj_5953), 
          .S1(n274_adj_5952));
    defparam _add_1_1244_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_13 (.A0(phase_inc_gen[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[13]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15681), .COUT(n15682), .S0(n283_adj_5955), 
          .S1(n280_adj_5954));
    defparam _add_1_1244_add_4_13.INIT0 = 16'h555f;
    defparam _add_1_1244_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_13.INJECT1_1 = "NO";
    LUT4 i1545_2_lut_3_lut_4_lut_4_lut (.A(led_c_3), .B(n17150), .C(n16220), 
         .D(led_c_4), .Z(n11259)) /* synthesis lut_function=(!(A+!(B+!((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i1545_2_lut_3_lut_4_lut_4_lut.init = 16'h4454;
    LUT4 i1_3_lut_3_lut (.A(led_c_3), .B(led_c_0), .C(led_c_4), .Z(n16451)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i1_3_lut_3_lut.init = 16'h5454;
    LUT4 mux_251_i59_4_lut (.A(n11393), .B(n145_adj_5909), .C(n17136), 
         .D(n2244), .Z(n1986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i59_4_lut.init = 16'hcfca;
    LUT4 i1637_3_lut_4_lut (.A(n17288), .B(n17150), .C(led_c_3), .D(n202), 
         .Z(n11359)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1637_3_lut_4_lut.init = 16'hf707;
    LUT4 i2507_2_lut_2_lut (.A(led_c_3), .B(n268), .Z(n2094)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i2507_2_lut_2_lut.init = 16'hdddd;
    LUT4 mux_251_i60_4_lut (.A(n11395), .B(n142_adj_5908), .C(n17136), 
         .D(n2244), .Z(n1985)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i60_4_lut.init = 16'hc0ca;
    LUT4 i4698_2_lut (.A(integrator1[0]), .B(mix_sinewave[0]), .Z(integrator1_71__N_418[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4698_2_lut.init = 16'h6666;
    CCU2C _add_1_1244_add_4_11 (.A0(phase_inc_gen[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15680), .COUT(n15681), .S0(n289_adj_5957), 
          .S1(n286_adj_5956));
    defparam _add_1_1244_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1244_add_4_11.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_11.INJECT1_1 = "NO";
    LUT4 i1631_3_lut_4_lut (.A(n17288), .B(n17150), .C(n17289), .D(n211), 
         .Z(n11353)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1631_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_251_i57_4_lut (.A(n2187), .B(n151_adj_5911), .C(n17136), 
         .D(n2244), .Z(n1988)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i57_4_lut.init = 16'hc0ca;
    LUT4 i2525_2_lut_2_lut (.A(led_c_3), .B(n295), .Z(n2237)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i2525_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1884_4_lut (.A(n148_adj_5910), .B(n142), .C(led_c_3), .D(n17144), 
         .Z(n11618)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1884_4_lut.init = 16'hcac0;
    LUT4 mux_251_i55_4_lut (.A(n11387), .B(n157_adj_5913), .C(n17136), 
         .D(n2244), .Z(n1990)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i55_4_lut.init = 16'hcfca;
    LUT4 i2545_2_lut_2_lut (.A(led_c_3), .B(n145), .Z(n2187)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i2545_2_lut_2_lut.init = 16'hdddd;
    LUT4 mux_251_i56_4_lut (.A(n2054), .B(n154_adj_5912), .C(n17136), 
         .D(n11259), .Z(n1989)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i56_4_lut.init = 16'hcfca;
    CCU2C _add_1_1244_add_4_9 (.A0(phase_inc_gen[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15679), .COUT(n15680), .S0(n295_adj_5959), 
          .S1(n292_adj_5958));
    defparam _add_1_1244_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1244_add_4_9.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_9.INJECT1_1 = "NO";
    LUT4 i2510_2_lut_2_lut (.A(led_c_3), .B(n181), .Z(n2065)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i2510_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2512_2_lut (.A(n148), .B(n17289), .Z(n2054)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i2512_2_lut.init = 16'h8888;
    LUT4 i27_3_lut_3_lut_adj_199 (.A(led_c_3), .B(n17150), .C(n193), .Z(n13_adj_5726)) /* synthesis lut_function=(!(A (C)+!A !(B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i27_3_lut_3_lut_adj_199.init = 16'h4e4e;
    CCU2C _add_1_1244_add_4_7 (.A0(phase_inc_gen[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15678), .COUT(n15679), .S0(n301_adj_5961), 
          .S1(n298_adj_5960));
    defparam _add_1_1244_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1244_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_7.INJECT1_1 = "NO";
    LUT4 i2537_2_lut_2_lut (.A(led_c_3), .B(n226), .Z(n2214)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i2537_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1882_4_lut (.A(n163_adj_5915), .B(n157), .C(led_c_3), .D(n17144), 
         .Z(n11616)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1882_4_lut.init = 16'hcac0;
    CCU2C _add_1_1244_add_4_5 (.A0(phase_inc_gen[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15677), .COUT(n15678), .S0(n307), .S1(n304));
    defparam _add_1_1244_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1244_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_3 (.A0(phase_inc_gen[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15676), .COUT(n15677), .S0(n313), .S1(n310));
    defparam _add_1_1244_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1244_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1244_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1244_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(phase_inc_gen[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15676), .S1(n316));
    defparam _add_1_1244_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1244_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1244_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1244_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_14 (.A0(integrator4[47]), .B0(integrator3[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[48]), .B1(integrator3[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15265), .COUT(n15266), .S0(n150_adj_5113), 
          .S1(n147_adj_5112));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_12 (.A0(integrator4[45]), .B0(integrator3[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[46]), .B1(integrator3[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15264), .COUT(n15265), .S0(n156_adj_5115), 
          .S1(n153_adj_5114));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_10 (.A0(integrator4[43]), .B0(integrator3[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[44]), .B1(integrator3[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15263), .COUT(n15264), .S0(n162_adj_5117), 
          .S1(n159_adj_5116));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_8 (.A0(integrator4[41]), .B0(integrator3[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[42]), .B1(integrator3[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15262), .COUT(n15263), .S0(n168_adj_5119), 
          .S1(n165_adj_5118));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_6 (.A0(integrator4[39]), .B0(integrator3[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[40]), .B1(integrator3[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15261), .COUT(n15262), .S0(n174_adj_5121), 
          .S1(n171_adj_5120));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_4 (.A0(integrator4[37]), .B0(integrator3[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator4[38]), .B1(integrator3[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15260), .COUT(n15261), .S0(n180_adj_5123), 
          .S1(n177_adj_5122));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1265_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1265_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator4[36]), .B1(integrator3[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15260), .S1(n183_adj_5124));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1265_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1265_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1265_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1265_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_38 (.A0(comb_d9_adj_6032[35]), .B0(comb9_adj_6031[35]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15259), .S1(cout_adj_5125));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1268_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_36 (.A0(comb_d9_adj_6032[33]), .B0(comb9_adj_6031[33]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[34]), .B1(comb9_adj_6031[34]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15258), .COUT(n15259));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_34 (.A0(comb_d9_adj_6032[31]), .B0(comb9_adj_6031[31]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[32]), .B1(comb9_adj_6031[32]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15257), .COUT(n15258));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_32 (.A0(comb_d9_adj_6032[29]), .B0(comb9_adj_6031[29]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[30]), .B1(comb9_adj_6031[30]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15256), .COUT(n15257));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_30 (.A0(comb_d9_adj_6032[27]), .B0(comb9_adj_6031[27]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[28]), .B1(comb9_adj_6031[28]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15255), .COUT(n15256));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_28 (.A0(comb_d9_adj_6032[25]), .B0(comb9_adj_6031[25]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[26]), .B1(comb9_adj_6031[26]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15254), .COUT(n15255));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_26 (.A0(comb_d9_adj_6032[23]), .B0(comb9_adj_6031[23]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[24]), .B1(comb9_adj_6031[24]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15253), .COUT(n15254));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_24 (.A0(comb_d9_adj_6032[21]), .B0(comb9_adj_6031[21]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[22]), .B1(comb9_adj_6031[22]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15252), .COUT(n15253));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_22 (.A0(comb_d9_adj_6032[19]), .B0(comb9_adj_6031[19]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[20]), .B1(comb9_adj_6031[20]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15251), .COUT(n15252));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_20 (.A0(comb_d9_adj_6032[17]), .B0(comb9_adj_6031[17]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[18]), .B1(comb9_adj_6031[18]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15250), .COUT(n15251));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_18 (.A0(comb_d9_adj_6032[15]), .B0(comb9_adj_6031[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[16]), .B1(comb9_adj_6031[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15249), .COUT(n15250));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_16 (.A0(comb_d9_adj_6032[13]), .B0(comb9_adj_6031[13]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[14]), .B1(comb9_adj_6031[14]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15248), .COUT(n15249));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_14 (.A0(comb_d9_adj_6032[11]), .B0(comb9_adj_6031[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[12]), .B1(comb9_adj_6031[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15247), .COUT(n15248));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_12 (.A0(comb_d9_adj_6032[9]), .B0(comb9_adj_6031[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[10]), .B1(comb9_adj_6031[10]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15246), .COUT(n15247));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_10 (.A0(comb_d9_adj_6032[7]), .B0(comb9_adj_6031[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[8]), .B1(comb9_adj_6031[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15245), .COUT(n15246));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_8 (.A0(comb_d9_adj_6032[5]), .B0(comb9_adj_6031[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[6]), .B1(comb9_adj_6031[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15244), .COUT(n15245));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_6 (.A0(comb_d9_adj_6032[3]), .B0(comb9_adj_6031[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[4]), .B1(comb9_adj_6031[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15243), .COUT(n15244));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_4 (.A0(comb_d9_adj_6032[1]), .B0(comb9_adj_6031[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d9_adj_6032[2]), .B1(comb9_adj_6031[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15242), .COUT(n15243));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1268_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1268_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d9_adj_6032[0]), .B1(comb9_adj_6031[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15242));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam _add_1_1268_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1268_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1268_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1268_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15241), .S0(cout_adj_5126));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_1271_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_1271_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_36 (.A0(integrator1[34]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[35]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15240), .COUT(n15241), .S0(integrator1_71__N_418[34]), 
          .S1(integrator1_71__N_418[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_34 (.A0(integrator1[32]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[33]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15239), .COUT(n15240), .S0(integrator1_71__N_418[32]), 
          .S1(integrator1_71__N_418[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_32 (.A0(integrator1[30]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[31]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15238), .COUT(n15239), .S0(integrator1_71__N_418[30]), 
          .S1(integrator1_71__N_418[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_30 (.A0(integrator1[28]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[29]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15237), .COUT(n15238), .S0(integrator1_71__N_418[28]), 
          .S1(integrator1_71__N_418[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_28 (.A0(integrator1[26]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[27]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15236), .COUT(n15237), .S0(integrator1_71__N_418[26]), 
          .S1(integrator1_71__N_418[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_26 (.A0(integrator1[24]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[25]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15235), .COUT(n15236), .S0(integrator1_71__N_418[24]), 
          .S1(integrator1_71__N_418[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_24 (.A0(integrator1[22]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[23]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15234), .COUT(n15235), .S0(integrator1_71__N_418[22]), 
          .S1(integrator1_71__N_418[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_22 (.A0(integrator1[20]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[21]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15233), .COUT(n15234), .S0(integrator1_71__N_418[20]), 
          .S1(integrator1_71__N_418[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_20 (.A0(integrator1[18]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[19]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15232), .COUT(n15233), .S0(integrator1_71__N_418[18]), 
          .S1(integrator1_71__N_418[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_18 (.A0(integrator1[16]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[17]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15231), .COUT(n15232), .S0(integrator1_71__N_418[16]), 
          .S1(integrator1_71__N_418[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_16 (.A0(integrator1[14]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[15]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15230), .COUT(n15231), .S0(integrator1_71__N_418[14]), 
          .S1(integrator1_71__N_418[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_14 (.A0(integrator1[12]), .B0(mix_sinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[13]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15229), .COUT(n15230), .S0(integrator1_71__N_418[12]), 
          .S1(integrator1_71__N_418[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_12 (.A0(integrator1[10]), .B0(mix_sinewave[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[11]), .B1(mix_sinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15228), .COUT(n15229), .S0(integrator1_71__N_418[10]), 
          .S1(integrator1_71__N_418[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_10 (.A0(integrator1[8]), .B0(mix_sinewave[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[9]), .B1(mix_sinewave[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15227), .COUT(n15228), .S0(integrator1_71__N_418[8]), 
          .S1(integrator1_71__N_418[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_8 (.A0(integrator1[6]), .B0(mix_sinewave[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[7]), .B1(mix_sinewave[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15226), .COUT(n15227), .S0(integrator1_71__N_418[6]), 
          .S1(integrator1_71__N_418[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_6 (.A0(integrator1[4]), .B0(mix_sinewave[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[5]), .B1(mix_sinewave[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15225), .COUT(n15226), .S0(integrator1_71__N_418[4]), 
          .S1(integrator1_71__N_418[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_4 (.A0(integrator1[2]), .B0(mix_sinewave[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[3]), .B1(mix_sinewave[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15224), .COUT(n15225), .S0(integrator1_71__N_418[2]), 
          .S1(integrator1_71__N_418[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1271_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1271_add_4_2 (.A0(integrator1[0]), .B0(mix_sinewave[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1[1]), .B1(mix_sinewave[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15224), .S1(integrator1_71__N_418[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1271_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_1271_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1271_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1271_add_4_2.INJECT1_1 = "NO";
    LUT4 i1623_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(led_c_3), .D(n223), 
         .Z(n11345)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1623_3_lut_4_lut.init = 16'hf808;
    CCU2C _add_1_add_4_38 (.A0(integrator5[71]), .B0(integrator4[71]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15222), .S0(n78_adj_5127));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_36 (.A0(integrator5[69]), .B0(integrator4[69]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[70]), .B1(integrator4[70]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15221), .COUT(n15222), .S0(n84_adj_5129), 
          .S1(n81_adj_5128));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_34 (.A0(integrator5[67]), .B0(integrator4[67]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[68]), .B1(integrator4[68]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15220), .COUT(n15221), .S0(n90_adj_5131), 
          .S1(n87_adj_5130));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_32 (.A0(integrator5[65]), .B0(integrator4[65]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[66]), .B1(integrator4[66]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15219), .COUT(n15220), .S0(n96_adj_5133), 
          .S1(n93_adj_5132));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_30 (.A0(integrator5[63]), .B0(integrator4[63]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[64]), .B1(integrator4[64]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15218), .COUT(n15219), .S0(n102_adj_5135), 
          .S1(n99_adj_5134));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_28 (.A0(integrator5[61]), .B0(integrator4[61]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[62]), .B1(integrator4[62]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15217), .COUT(n15218), .S0(n108_adj_5137), 
          .S1(n105_adj_5136));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_26 (.A0(integrator5[59]), .B0(integrator4[59]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[60]), .B1(integrator4[60]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15216), .COUT(n15217), .S0(n114_adj_5139), 
          .S1(n111_adj_5138));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_24 (.A0(integrator5[57]), .B0(integrator4[57]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[58]), .B1(integrator4[58]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15215), .COUT(n15216), .S0(n120_adj_5141), 
          .S1(n117_adj_5140));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_22 (.A0(integrator5[55]), .B0(integrator4[55]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[56]), .B1(integrator4[56]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15214), .COUT(n15215), .S0(n126_adj_5143), 
          .S1(n123_adj_5142));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_20 (.A0(integrator5[53]), .B0(integrator4[53]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[54]), .B1(integrator4[54]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15213), .COUT(n15214), .S0(n132_adj_5145), 
          .S1(n129_adj_5144));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_18 (.A0(integrator5[51]), .B0(integrator4[51]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[52]), .B1(integrator4[52]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15212), .COUT(n15213), .S0(n138_adj_5147), 
          .S1(n135_adj_5146));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_16 (.A0(integrator5[49]), .B0(integrator4[49]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[50]), .B1(integrator4[50]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15211), .COUT(n15212), .S0(n144_adj_5149), 
          .S1(n141_adj_5148));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_14 (.A0(integrator5[47]), .B0(integrator4[47]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[48]), .B1(integrator4[48]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15210), .COUT(n15211), .S0(n150_adj_5151), 
          .S1(n147_adj_5150));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_12 (.A0(integrator5[45]), .B0(integrator4[45]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[46]), .B1(integrator4[46]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15209), .COUT(n15210), .S0(n156_adj_5153), 
          .S1(n153_adj_5152));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_10 (.A0(integrator5[43]), .B0(integrator4[43]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[44]), .B1(integrator4[44]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15208), .COUT(n15209), .S0(n162_adj_5155), 
          .S1(n159_adj_5154));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_8 (.A0(integrator5[41]), .B0(integrator4[41]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[42]), .B1(integrator4[42]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15207), .COUT(n15208), .S0(n168_adj_5157), 
          .S1(n165_adj_5156));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_6 (.A0(integrator5[39]), .B0(integrator4[39]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[40]), .B1(integrator4[40]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15206), .COUT(n15207), .S0(n174_adj_5159), 
          .S1(n171_adj_5158));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_4 (.A0(integrator5[37]), .B0(integrator4[37]), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator5[38]), .B1(integrator4[38]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15205), .COUT(n15206), .S0(n180_adj_5161), 
          .S1(n177_adj_5160));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(integrator5[36]), .B1(integrator4[36]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n15205), .S1(n183_adj_5162));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(70[20:45])
    defparam _add_1_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15204), .S0(cout_adj_5163));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_999_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_999_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_36 (.A0(integrator2_adj_6021[34]), .B0(integrator1_adj_6020[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[35]), .B1(integrator1_adj_6020[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15203), .COUT(n15204), .S0(integrator2_71__N_490_adj_6037[34]), 
          .S1(integrator2_71__N_490_adj_6037[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_34 (.A0(integrator2_adj_6021[32]), .B0(integrator1_adj_6020[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[33]), .B1(integrator1_adj_6020[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15202), .COUT(n15203), .S0(integrator2_71__N_490_adj_6037[32]), 
          .S1(integrator2_71__N_490_adj_6037[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_32 (.A0(integrator2_adj_6021[30]), .B0(integrator1_adj_6020[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[31]), .B1(integrator1_adj_6020[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15201), .COUT(n15202), .S0(integrator2_71__N_490_adj_6037[30]), 
          .S1(integrator2_71__N_490_adj_6037[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_30 (.A0(integrator2_adj_6021[28]), .B0(integrator1_adj_6020[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[29]), .B1(integrator1_adj_6020[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15200), .COUT(n15201), .S0(integrator2_71__N_490_adj_6037[28]), 
          .S1(integrator2_71__N_490_adj_6037[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_28 (.A0(integrator2_adj_6021[26]), .B0(integrator1_adj_6020[26]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[27]), .B1(integrator1_adj_6020[27]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15199), .COUT(n15200), .S0(integrator2_71__N_490_adj_6037[26]), 
          .S1(integrator2_71__N_490_adj_6037[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_26 (.A0(integrator2_adj_6021[24]), .B0(integrator1_adj_6020[24]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[25]), .B1(integrator1_adj_6020[25]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15198), .COUT(n15199), .S0(integrator2_71__N_490_adj_6037[24]), 
          .S1(integrator2_71__N_490_adj_6037[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_24 (.A0(integrator2_adj_6021[22]), .B0(integrator1_adj_6020[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[23]), .B1(integrator1_adj_6020[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15197), .COUT(n15198), .S0(integrator2_71__N_490_adj_6037[22]), 
          .S1(integrator2_71__N_490_adj_6037[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_22 (.A0(integrator2_adj_6021[20]), .B0(integrator1_adj_6020[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[21]), .B1(integrator1_adj_6020[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15196), .COUT(n15197), .S0(integrator2_71__N_490_adj_6037[20]), 
          .S1(integrator2_71__N_490_adj_6037[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_20 (.A0(integrator2_adj_6021[18]), .B0(integrator1_adj_6020[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[19]), .B1(integrator1_adj_6020[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15195), .COUT(n15196), .S0(integrator2_71__N_490_adj_6037[18]), 
          .S1(integrator2_71__N_490_adj_6037[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_18 (.A0(integrator2_adj_6021[16]), .B0(integrator1_adj_6020[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[17]), .B1(integrator1_adj_6020[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15194), .COUT(n15195), .S0(integrator2_71__N_490_adj_6037[16]), 
          .S1(integrator2_71__N_490_adj_6037[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_16 (.A0(integrator2_adj_6021[14]), .B0(integrator1_adj_6020[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[15]), .B1(integrator1_adj_6020[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15193), .COUT(n15194), .S0(integrator2_71__N_490_adj_6037[14]), 
          .S1(integrator2_71__N_490_adj_6037[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_14 (.A0(integrator2_adj_6021[12]), .B0(integrator1_adj_6020[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[13]), .B1(integrator1_adj_6020[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15192), .COUT(n15193), .S0(integrator2_71__N_490_adj_6037[12]), 
          .S1(integrator2_71__N_490_adj_6037[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_12 (.A0(integrator2_adj_6021[10]), .B0(integrator1_adj_6020[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[11]), .B1(integrator1_adj_6020[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15191), .COUT(n15192), .S0(integrator2_71__N_490_adj_6037[10]), 
          .S1(integrator2_71__N_490_adj_6037[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_10 (.A0(integrator2_adj_6021[8]), .B0(integrator1_adj_6020[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[9]), .B1(integrator1_adj_6020[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15190), .COUT(n15191), .S0(integrator2_71__N_490_adj_6037[8]), 
          .S1(integrator2_71__N_490_adj_6037[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_8 (.A0(integrator2_adj_6021[6]), .B0(integrator1_adj_6020[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[7]), .B1(integrator1_adj_6020[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15189), .COUT(n15190), .S0(integrator2_71__N_490_adj_6037[6]), 
          .S1(integrator2_71__N_490_adj_6037[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_6 (.A0(integrator2_adj_6021[4]), .B0(integrator1_adj_6020[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[5]), .B1(integrator1_adj_6020[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15188), .COUT(n15189), .S0(integrator2_71__N_490_adj_6037[4]), 
          .S1(integrator2_71__N_490_adj_6037[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_4 (.A0(integrator2_adj_6021[2]), .B0(integrator1_adj_6020[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[3]), .B1(integrator1_adj_6020[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15187), .COUT(n15188), .S0(integrator2_71__N_490_adj_6037[2]), 
          .S1(integrator2_71__N_490_adj_6037[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_999_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_999_add_4_2 (.A0(integrator2_adj_6021[0]), .B0(integrator1_adj_6020[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[1]), .B1(integrator1_adj_6020[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15187), .S1(integrator2_71__N_490_adj_6037[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_999_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_999_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_999_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_999_add_4_2.INJECT1_1 = "NO";
    LUT4 mux_251_i54_4_lut (.A(n11385), .B(n160_adj_5914), .C(n17136), 
         .D(n2244), .Z(n1991)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i54_4_lut.init = 16'hc0ca;
    CCU2C _add_1_1118_add_4_38 (.A0(comb_d6[35]), .B0(comb6[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15185), .S0(comb7_71__N_1523[35]), .S1(cout_adj_4985));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1118_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_36 (.A0(comb_d6[33]), .B0(comb6[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[34]), .B1(comb6[34]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15184), .COUT(n15185), .S0(comb7_71__N_1523[33]), 
          .S1(comb7_71__N_1523[34]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_34 (.A0(comb_d6[31]), .B0(comb6[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[32]), .B1(comb6[32]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15183), .COUT(n15184), .S0(comb7_71__N_1523[31]), 
          .S1(comb7_71__N_1523[32]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_32 (.A0(comb_d6[29]), .B0(comb6[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[30]), .B1(comb6[30]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15182), .COUT(n15183), .S0(comb7_71__N_1523[29]), 
          .S1(comb7_71__N_1523[30]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_30 (.A0(comb_d6[27]), .B0(comb6[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[28]), .B1(comb6[28]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15181), .COUT(n15182), .S0(comb7_71__N_1523[27]), 
          .S1(comb7_71__N_1523[28]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_28 (.A0(comb_d6[25]), .B0(comb6[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[26]), .B1(comb6[26]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15180), .COUT(n15181), .S0(comb7_71__N_1523[25]), 
          .S1(comb7_71__N_1523[26]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_26 (.A0(comb_d6[23]), .B0(comb6[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[24]), .B1(comb6[24]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15179), .COUT(n15180), .S0(comb7_71__N_1523[23]), 
          .S1(comb7_71__N_1523[24]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_24 (.A0(comb_d6[21]), .B0(comb6[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[22]), .B1(comb6[22]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15178), .COUT(n15179), .S0(comb7_71__N_1523[21]), 
          .S1(comb7_71__N_1523[22]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_22 (.A0(comb_d6[19]), .B0(comb6[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[20]), .B1(comb6[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15177), .COUT(n15178), .S0(comb7_71__N_1523[19]), 
          .S1(comb7_71__N_1523[20]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_20 (.A0(comb_d6[17]), .B0(comb6[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[18]), .B1(comb6[18]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15176), .COUT(n15177), .S0(comb7_71__N_1523[17]), 
          .S1(comb7_71__N_1523[18]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_18 (.A0(comb_d6[15]), .B0(comb6[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[16]), .B1(comb6[16]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15175), .COUT(n15176), .S0(comb7_71__N_1523[15]), 
          .S1(comb7_71__N_1523[16]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_16 (.A0(comb_d6[13]), .B0(comb6[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[14]), .B1(comb6[14]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15174), .COUT(n15175), .S0(comb7_71__N_1523[13]), 
          .S1(comb7_71__N_1523[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_14 (.A0(comb_d6[11]), .B0(comb6[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[12]), .B1(comb6[12]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15173), .COUT(n15174), .S0(comb7_71__N_1523[11]), 
          .S1(comb7_71__N_1523[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_12 (.A0(comb_d6[9]), .B0(comb6[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[10]), .B1(comb6[10]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15172), .COUT(n15173), .S0(comb7_71__N_1523[9]), 
          .S1(comb7_71__N_1523[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_10 (.A0(comb_d6[7]), .B0(comb6[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[8]), .B1(comb6[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15171), .COUT(n15172), .S0(comb7_71__N_1523[7]), 
          .S1(comb7_71__N_1523[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_8 (.A0(comb_d6[5]), .B0(comb6[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[6]), .B1(comb6[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15170), .COUT(n15171), .S0(comb7_71__N_1523[5]), 
          .S1(comb7_71__N_1523[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_6 (.A0(comb_d6[3]), .B0(comb6[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[4]), .B1(comb6[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15169), .COUT(n15170), .S0(comb7_71__N_1523[3]), 
          .S1(comb7_71__N_1523[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_4 (.A0(comb_d6[1]), .B0(comb6[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[2]), .B1(comb6[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15168), .COUT(n15169), .S0(comb7_71__N_1523[1]), 
          .S1(comb7_71__N_1523[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1118_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1118_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6[0]), .B1(comb6[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15168), .S1(comb7_71__N_1523[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1118_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1118_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1118_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1118_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_38 (.A0(comb_d7[35]), .B0(comb7[35]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15167), .S0(comb8_71__N_1595[35]), .S1(cout_adj_4986));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1121_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_36 (.A0(comb_d7[33]), .B0(comb7[33]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[34]), .B1(comb7[34]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15166), .COUT(n15167), .S0(comb8_71__N_1595[33]), 
          .S1(comb8_71__N_1595[34]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_34 (.A0(comb_d7[31]), .B0(comb7[31]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[32]), .B1(comb7[32]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15165), .COUT(n15166), .S0(comb8_71__N_1595[31]), 
          .S1(comb8_71__N_1595[32]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_32 (.A0(comb_d7[29]), .B0(comb7[29]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[30]), .B1(comb7[30]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15164), .COUT(n15165), .S0(comb8_71__N_1595[29]), 
          .S1(comb8_71__N_1595[30]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_30 (.A0(comb_d7[27]), .B0(comb7[27]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[28]), .B1(comb7[28]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15163), .COUT(n15164), .S0(comb8_71__N_1595[27]), 
          .S1(comb8_71__N_1595[28]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_28 (.A0(comb_d7[25]), .B0(comb7[25]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[26]), .B1(comb7[26]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15162), .COUT(n15163), .S0(comb8_71__N_1595[25]), 
          .S1(comb8_71__N_1595[26]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_26 (.A0(comb_d7[23]), .B0(comb7[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[24]), .B1(comb7[24]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15161), .COUT(n15162), .S0(comb8_71__N_1595[23]), 
          .S1(comb8_71__N_1595[24]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_24 (.A0(comb_d7[21]), .B0(comb7[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[22]), .B1(comb7[22]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15160), .COUT(n15161), .S0(comb8_71__N_1595[21]), 
          .S1(comb8_71__N_1595[22]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_22 (.A0(comb_d7[19]), .B0(comb7[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[20]), .B1(comb7[20]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15159), .COUT(n15160), .S0(comb8_71__N_1595[19]), 
          .S1(comb8_71__N_1595[20]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_20 (.A0(comb_d7[17]), .B0(comb7[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[18]), .B1(comb7[18]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15158), .COUT(n15159), .S0(comb8_71__N_1595[17]), 
          .S1(comb8_71__N_1595[18]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_18 (.A0(comb_d7[15]), .B0(comb7[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[16]), .B1(comb7[16]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15157), .COUT(n15158), .S0(comb8_71__N_1595[15]), 
          .S1(comb8_71__N_1595[16]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_16 (.A0(comb_d7[13]), .B0(comb7[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[14]), .B1(comb7[14]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15156), .COUT(n15157), .S0(comb8_71__N_1595[13]), 
          .S1(comb8_71__N_1595[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_14 (.A0(comb_d7[11]), .B0(comb7[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[12]), .B1(comb7[12]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15155), .COUT(n15156), .S0(comb8_71__N_1595[11]), 
          .S1(comb8_71__N_1595[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_12 (.A0(comb_d7[9]), .B0(comb7[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[10]), .B1(comb7[10]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15154), .COUT(n15155), .S0(comb8_71__N_1595[9]), 
          .S1(comb8_71__N_1595[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_10 (.A0(comb_d7[7]), .B0(comb7[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[8]), .B1(comb7[8]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15153), .COUT(n15154), .S0(comb8_71__N_1595[7]), 
          .S1(comb8_71__N_1595[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_8 (.A0(comb_d7[5]), .B0(comb7[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[6]), .B1(comb7[6]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15152), .COUT(n15153), .S0(comb8_71__N_1595[5]), 
          .S1(comb8_71__N_1595[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_6 (.A0(comb_d7[3]), .B0(comb7[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[4]), .B1(comb7[4]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15151), .COUT(n15152), .S0(comb8_71__N_1595[3]), 
          .S1(comb8_71__N_1595[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_4 (.A0(comb_d7[1]), .B0(comb7[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[2]), .B1(comb7[2]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15150), .COUT(n15151), .S0(comb8_71__N_1595[1]), 
          .S1(comb8_71__N_1595[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1121_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1121_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7[0]), .B1(comb7[0]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15150), .S1(comb8_71__N_1595[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1121_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1121_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1121_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1121_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1253_add_4_16 (.A0(amdemod_d_11__N_1871[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15149), .S0(n34_adj_4983));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1253_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1253_add_4_16.INIT1 = 16'h0000;
    defparam _add_1_1253_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1253_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1253_add_4_14 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1871[9]), .D0(VCC_net), .A1(amdemod_d_11__N_1871[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n15148), .COUT(n15149), 
          .S0(n40));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1253_add_4_14.INIT0 = 16'he1e1;
    defparam _add_1_1253_add_4_14.INIT1 = 16'h555f;
    defparam _add_1_1253_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1253_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1253_add_4_12 (.A0(n17134), .B0(amdemod_d_11__N_1871[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(n17137), .B1(amdemod_d_11__N_1871[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15147), .COUT(n15148), .S0(n46), 
          .S1(n43));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1253_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1253_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1253_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1253_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1253_add_4_10 (.A0(n17132), .B0(amdemod_d_11__N_1871[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1871[6]), .B1(amdemod_d_11__N_1841[11]), 
          .C1(n17134), .D1(amdemod_d_11__N_1840[11]), .CIN(n15146), .COUT(n15147), 
          .S0(n52), .S1(n49));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1253_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1253_add_4_10.INIT1 = 16'h656a;
    defparam _add_1_1253_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1253_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1253_add_4_8 (.A0(n17130), .B0(amdemod_d_11__N_1871[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1871[4]), .B1(amdemod_d_11__N_1851[13]), 
          .C1(n17132), .D1(amdemod_d_11__N_1850[13]), .CIN(n15145), .COUT(n15146), 
          .S0(n58_adj_4765), .S1(n55));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1253_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1253_add_4_8.INIT1 = 16'h656a;
    defparam _add_1_1253_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1253_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1253_add_4_6 (.A0(n17128), .B0(amdemod_d_11__N_1871[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1871[2]), .B1(amdemod_d_11__N_1861[13]), 
          .C1(n17130), .D1(amdemod_d_11__N_1860[13]), .CIN(n15144), .COUT(n15145), 
          .S0(n64_adj_4762), .S1(n61_adj_4764));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1253_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1253_add_4_6.INIT1 = 16'h656a;
    defparam _add_1_1253_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1253_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1253_add_4_4 (.A0(n17127), .B0(square_sum[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(amdemod_d_11__N_1871[0]), .B1(amdemod_d_11__N_1871[13]), 
          .C1(n17128), .D1(amdemod_d_11__N_1870[13]), .CIN(n15143), .COUT(n15144), 
          .S0(n70_adj_4759), .S1(n67_adj_4760));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1253_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1253_add_4_4.INIT1 = 16'h656a;
    defparam _add_1_1253_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1253_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1253_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15143), .S1(n73_adj_4751));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1253_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1253_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_1253_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1253_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_38 (.A0(integrator1_adj_6020[71]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15142), .S0(n78_adj_4987));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1124_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_36 (.A0(integrator1_adj_6020[69]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[70]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15141), .COUT(n15142), .S0(n84_adj_4989), 
          .S1(n81_adj_4988));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_34 (.A0(integrator1_adj_6020[67]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[68]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15140), .COUT(n15141), .S0(n90_adj_4991), 
          .S1(n87_adj_4990));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_32 (.A0(integrator1_adj_6020[65]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[66]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15139), .COUT(n15140), .S0(n96_adj_4993), 
          .S1(n93_adj_4992));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_30 (.A0(integrator1_adj_6020[63]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[64]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15138), .COUT(n15139), .S0(n102_adj_4995), 
          .S1(n99_adj_4994));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_28 (.A0(integrator1_adj_6020[61]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[62]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15137), .COUT(n15138), .S0(n108_adj_4997), 
          .S1(n105_adj_4996));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_26 (.A0(integrator1_adj_6020[59]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[60]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15136), .COUT(n15137), .S0(n114_adj_4999), 
          .S1(n111_adj_4998));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_24 (.A0(integrator1_adj_6020[57]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[58]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15135), .COUT(n15136), .S0(n120_adj_5001), 
          .S1(n117_adj_5000));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_22 (.A0(integrator1_adj_6020[55]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[56]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15134), .COUT(n15135), .S0(n126_adj_5003), 
          .S1(n123_adj_5002));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_20 (.A0(integrator1_adj_6020[53]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[54]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15133), .COUT(n15134), .S0(n132_adj_5005), 
          .S1(n129_adj_5004));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_18 (.A0(integrator1_adj_6020[51]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[52]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15132), .COUT(n15133), .S0(n138_adj_5007), 
          .S1(n135_adj_5006));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_16 (.A0(integrator1_adj_6020[49]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[50]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15131), .COUT(n15132), .S0(n144_adj_5009), 
          .S1(n141_adj_5008));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_14 (.A0(integrator1_adj_6020[47]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[48]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15130), .COUT(n15131), .S0(n150_adj_5011), 
          .S1(n147_adj_5010));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_12 (.A0(integrator1_adj_6020[45]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[46]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15129), .COUT(n15130), .S0(n156_adj_5013), 
          .S1(n153_adj_5012));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_10 (.A0(integrator1_adj_6020[43]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[44]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15128), .COUT(n15129), .S0(n162_adj_5015), 
          .S1(n159_adj_5014));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_8 (.A0(integrator1_adj_6020[41]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[42]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15127), .COUT(n15128), .S0(n168_adj_5017), 
          .S1(n165_adj_5016));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_6 (.A0(integrator1_adj_6020[39]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[40]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15126), .COUT(n15127), .S0(n174_adj_5019), 
          .S1(n171_adj_5018));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_4 (.A0(integrator1_adj_6020[37]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[38]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15125), .COUT(n15126), .S0(n180_adj_5021), 
          .S1(n177_adj_5020));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1124_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1124_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator1_adj_6020[36]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15125), .S1(n183_adj_5022));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_1124_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1124_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1124_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1124_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_38 (.A0(integrator2_adj_6021[71]), .B0(integrator1_adj_6020[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15124), .S0(n78_adj_5023));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_38.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1127_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_36 (.A0(integrator2_adj_6021[69]), .B0(integrator1_adj_6020[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[70]), .B1(integrator1_adj_6020[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15123), .COUT(n15124), .S0(n84_adj_5025), 
          .S1(n81_adj_5024));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_34 (.A0(integrator2_adj_6021[67]), .B0(integrator1_adj_6020[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[68]), .B1(integrator1_adj_6020[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15122), .COUT(n15123), .S0(n90_adj_5027), 
          .S1(n87_adj_5026));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_32 (.A0(integrator2_adj_6021[65]), .B0(integrator1_adj_6020[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[66]), .B1(integrator1_adj_6020[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15121), .COUT(n15122), .S0(n96_adj_5029), 
          .S1(n93_adj_5028));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_30 (.A0(integrator2_adj_6021[63]), .B0(integrator1_adj_6020[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[64]), .B1(integrator1_adj_6020[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15120), .COUT(n15121), .S0(n102_adj_5031), 
          .S1(n99_adj_5030));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_28 (.A0(integrator2_adj_6021[61]), .B0(integrator1_adj_6020[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[62]), .B1(integrator1_adj_6020[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15119), .COUT(n15120), .S0(n108_adj_5033), 
          .S1(n105_adj_5032));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_26 (.A0(integrator2_adj_6021[59]), .B0(integrator1_adj_6020[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[60]), .B1(integrator1_adj_6020[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15118), .COUT(n15119), .S0(n114_adj_5035), 
          .S1(n111_adj_5034));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_24 (.A0(integrator2_adj_6021[57]), .B0(integrator1_adj_6020[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[58]), .B1(integrator1_adj_6020[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15117), .COUT(n15118), .S0(n120_adj_5037), 
          .S1(n117_adj_5036));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_22 (.A0(integrator2_adj_6021[55]), .B0(integrator1_adj_6020[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[56]), .B1(integrator1_adj_6020[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15116), .COUT(n15117), .S0(n126_adj_5039), 
          .S1(n123_adj_5038));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_20 (.A0(integrator2_adj_6021[53]), .B0(integrator1_adj_6020[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[54]), .B1(integrator1_adj_6020[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15115), .COUT(n15116), .S0(n132_adj_5041), 
          .S1(n129_adj_5040));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_18 (.A0(integrator2_adj_6021[51]), .B0(integrator1_adj_6020[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[52]), .B1(integrator1_adj_6020[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15114), .COUT(n15115), .S0(n138_adj_5043), 
          .S1(n135_adj_5042));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_16 (.A0(integrator2_adj_6021[49]), .B0(integrator1_adj_6020[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[50]), .B1(integrator1_adj_6020[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15113), .COUT(n15114), .S0(n144_adj_5045), 
          .S1(n141_adj_5044));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_14 (.A0(integrator2_adj_6021[47]), .B0(integrator1_adj_6020[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[48]), .B1(integrator1_adj_6020[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15112), .COUT(n15113), .S0(n150_adj_5047), 
          .S1(n147_adj_5046));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_12 (.A0(integrator2_adj_6021[45]), .B0(integrator1_adj_6020[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[46]), .B1(integrator1_adj_6020[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15111), .COUT(n15112), .S0(n156_adj_5049), 
          .S1(n153_adj_5048));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_10 (.A0(integrator2_adj_6021[43]), .B0(integrator1_adj_6020[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[44]), .B1(integrator1_adj_6020[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15110), .COUT(n15111), .S0(n162_adj_5051), 
          .S1(n159_adj_5050));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_8 (.A0(integrator2_adj_6021[41]), .B0(integrator1_adj_6020[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[42]), .B1(integrator1_adj_6020[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15109), .COUT(n15110), .S0(n168_adj_5053), 
          .S1(n165_adj_5052));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_6 (.A0(integrator2_adj_6021[39]), .B0(integrator1_adj_6020[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[40]), .B1(integrator1_adj_6020[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15108), .COUT(n15109), .S0(n174_adj_5055), 
          .S1(n171_adj_5054));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_4 (.A0(integrator2_adj_6021[37]), .B0(integrator1_adj_6020[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2_adj_6021[38]), .B1(integrator1_adj_6020[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15107), .COUT(n15108), .S0(n180_adj_5057), 
          .S1(n177_adj_5056));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1127_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1127_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator2_adj_6021[36]), .B1(integrator1_adj_6020[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15107), .S1(n183_adj_5058));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_1127_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1127_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1127_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1127_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1256_add_4_15 (.A0(amdemod_d_11__N_1841[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15106), .S0(n32_adj_4742));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1256_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1256_add_4_15.INIT1 = 16'h0000;
    defparam _add_1_1256_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1256_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1256_add_4_13 (.A0(amdemod_d_11__N_1841[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1841[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15105), .COUT(n15106), .S0(n38_adj_4741));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1256_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1256_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1256_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1256_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1256_add_4_11 (.A0(amdemod_d_11__N_1841[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1841[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15104), .COUT(n15105), .S0(n44_adj_4739), 
          .S1(n41_adj_4740));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1256_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1256_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1256_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1256_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1256_add_4_9 (.A0(amdemod_d_11__N_1841[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1841[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15103), .COUT(n15104), .S0(n50_adj_4737), 
          .S1(n47_adj_4738));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1256_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1256_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1256_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1256_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1256_add_4_7 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1841[3]), .D0(VCC_net), .A1(amdemod_d_11__N_1841[4]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n15102), .COUT(n15103), 
          .S0(n56_adj_4735), .S1(n53_adj_4736));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1256_add_4_7.INIT0 = 16'h1e1e;
    defparam _add_1_1256_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1256_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1256_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1256_add_4_5 (.A0(n17134), .B0(amdemod_d_11__N_1841[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1841[2]), .B1(n17162), 
          .C1(n17279), .D1(n17146), .CIN(n15101), .COUT(n15102), .S0(n62_adj_4733), 
          .S1(n59_adj_4734));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1256_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1256_add_4_5.INIT1 = 16'h596a;
    defparam _add_1_1256_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1256_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1256_add_4_3 (.A0(square_sum[15]), .B0(amdemod_d_11__N_1841[11]), 
          .C0(n17134), .D0(amdemod_d_11__N_1840[11]), .A1(n17133), .B1(amdemod_d_11__N_1841[0]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15100), .COUT(n15101), .S0(n68_adj_4731), 
          .S1(n65_adj_4732));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1256_add_4_3.INIT0 = 16'h656a;
    defparam _add_1_1256_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1256_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1256_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1256_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15100), .S1(n71_adj_4730));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1256_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1256_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1256_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1256_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_37 (.A0(comb7_adj_6027[70]), .B0(cout_adj_5309), 
          .C0(n81_adj_5728), .D0(n3_adj_4911), .A1(comb7_adj_6027[71]), 
          .B1(cout_adj_5309), .C1(n78_adj_5727), .D1(n2_adj_4910), .CIN(n15098), 
          .S0(comb8_71__N_1595_adj_6054[70]), .S1(comb8_71__N_1595_adj_6054[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_35 (.A0(comb7_adj_6027[68]), .B0(cout_adj_5309), 
          .C0(n87_adj_5730), .D0(n5_adj_4913), .A1(comb7_adj_6027[69]), 
          .B1(cout_adj_5309), .C1(n84_adj_5729), .D1(n4_adj_4912), .CIN(n15097), 
          .COUT(n15098), .S0(comb8_71__N_1595_adj_6054[68]), .S1(comb8_71__N_1595_adj_6054[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_33 (.A0(comb7_adj_6027[66]), .B0(cout_adj_5309), 
          .C0(n93_adj_5732), .D0(n7_adj_4915), .A1(comb7_adj_6027[67]), 
          .B1(cout_adj_5309), .C1(n90_adj_5731), .D1(n6_adj_4914), .CIN(n15096), 
          .COUT(n15097), .S0(comb8_71__N_1595_adj_6054[66]), .S1(comb8_71__N_1595_adj_6054[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_31 (.A0(comb7_adj_6027[64]), .B0(cout_adj_5309), 
          .C0(n99_adj_5734), .D0(n9_adj_4917), .A1(comb7_adj_6027[65]), 
          .B1(cout_adj_5309), .C1(n96_adj_5733), .D1(n8_adj_4916), .CIN(n15095), 
          .COUT(n15096), .S0(comb8_71__N_1595_adj_6054[64]), .S1(comb8_71__N_1595_adj_6054[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_29 (.A0(comb7_adj_6027[62]), .B0(cout_adj_5309), 
          .C0(n105_adj_5736), .D0(n11_adj_4919), .A1(comb7_adj_6027[63]), 
          .B1(cout_adj_5309), .C1(n102_adj_5735), .D1(n10_adj_4918), .CIN(n15094), 
          .COUT(n15095), .S0(comb8_71__N_1595_adj_6054[62]), .S1(comb8_71__N_1595_adj_6054[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_27 (.A0(comb7_adj_6027[60]), .B0(cout_adj_5309), 
          .C0(n111_adj_5738), .D0(n13_adj_4921), .A1(comb7_adj_6027[61]), 
          .B1(cout_adj_5309), .C1(n108_adj_5737), .D1(n12_adj_4920), .CIN(n15093), 
          .COUT(n15094), .S0(comb8_71__N_1595_adj_6054[60]), .S1(comb8_71__N_1595_adj_6054[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_25 (.A0(comb7_adj_6027[58]), .B0(cout_adj_5309), 
          .C0(n117_adj_5740), .D0(n15_adj_4923), .A1(comb7_adj_6027[59]), 
          .B1(cout_adj_5309), .C1(n114_adj_5739), .D1(n14_adj_4922), .CIN(n15092), 
          .COUT(n15093), .S0(comb8_71__N_1595_adj_6054[58]), .S1(comb8_71__N_1595_adj_6054[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_23 (.A0(comb7_adj_6027[56]), .B0(cout_adj_5309), 
          .C0(n123_adj_5742), .D0(n17_adj_4925), .A1(comb7_adj_6027[57]), 
          .B1(cout_adj_5309), .C1(n120_adj_5741), .D1(n16_adj_4924), .CIN(n15091), 
          .COUT(n15092), .S0(comb8_71__N_1595_adj_6054[56]), .S1(comb8_71__N_1595_adj_6054[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_21 (.A0(comb7_adj_6027[54]), .B0(cout_adj_5309), 
          .C0(n129_adj_5744), .D0(n19_adj_4927), .A1(comb7_adj_6027[55]), 
          .B1(cout_adj_5309), .C1(n126_adj_5743), .D1(n18_adj_4926), .CIN(n15090), 
          .COUT(n15091), .S0(comb8_71__N_1595_adj_6054[54]), .S1(comb8_71__N_1595_adj_6054[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_19 (.A0(comb7_adj_6027[52]), .B0(cout_adj_5309), 
          .C0(n135_adj_5746), .D0(n21_adj_4929), .A1(comb7_adj_6027[53]), 
          .B1(cout_adj_5309), .C1(n132_adj_5745), .D1(n20_adj_4928), .CIN(n15089), 
          .COUT(n15090), .S0(comb8_71__N_1595_adj_6054[52]), .S1(comb8_71__N_1595_adj_6054[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_17 (.A0(comb7_adj_6027[50]), .B0(cout_adj_5309), 
          .C0(n141_adj_5748), .D0(n23_adj_4931), .A1(comb7_adj_6027[51]), 
          .B1(cout_adj_5309), .C1(n138_adj_5747), .D1(n22_adj_4930), .CIN(n15088), 
          .COUT(n15089), .S0(comb8_71__N_1595_adj_6054[50]), .S1(comb8_71__N_1595_adj_6054[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_15 (.A0(comb7_adj_6027[48]), .B0(cout_adj_5309), 
          .C0(n147_adj_5750), .D0(n25_adj_4933), .A1(comb7_adj_6027[49]), 
          .B1(cout_adj_5309), .C1(n144_adj_5749), .D1(n24_adj_4932), .CIN(n15087), 
          .COUT(n15088), .S0(comb8_71__N_1595_adj_6054[48]), .S1(comb8_71__N_1595_adj_6054[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_13 (.A0(comb7_adj_6027[46]), .B0(cout_adj_5309), 
          .C0(n153_adj_5752), .D0(n27_adj_4935), .A1(comb7_adj_6027[47]), 
          .B1(cout_adj_5309), .C1(n150_adj_5751), .D1(n26_adj_4934), .CIN(n15086), 
          .COUT(n15087), .S0(comb8_71__N_1595_adj_6054[46]), .S1(comb8_71__N_1595_adj_6054[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_11 (.A0(comb7_adj_6027[44]), .B0(cout_adj_5309), 
          .C0(n159_adj_5754), .D0(n29_adj_4937), .A1(comb7_adj_6027[45]), 
          .B1(cout_adj_5309), .C1(n156_adj_5753), .D1(n28_adj_4936), .CIN(n15085), 
          .COUT(n15086), .S0(comb8_71__N_1595_adj_6054[44]), .S1(comb8_71__N_1595_adj_6054[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_9 (.A0(comb7_adj_6027[42]), .B0(cout_adj_5309), 
          .C0(n165_adj_5756), .D0(n31_adj_4939), .A1(comb7_adj_6027[43]), 
          .B1(cout_adj_5309), .C1(n162_adj_5755), .D1(n30_adj_4938), .CIN(n15084), 
          .COUT(n15085), .S0(comb8_71__N_1595_adj_6054[42]), .S1(comb8_71__N_1595_adj_6054[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_7 (.A0(comb7_adj_6027[40]), .B0(cout_adj_5309), 
          .C0(n171_adj_5758), .D0(n33_adj_4941), .A1(comb7_adj_6027[41]), 
          .B1(cout_adj_5309), .C1(n168_adj_5757), .D1(n32_adj_4940), .CIN(n15083), 
          .COUT(n15084), .S0(comb8_71__N_1595_adj_6054[40]), .S1(comb8_71__N_1595_adj_6054[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_5 (.A0(comb7_adj_6027[38]), .B0(cout_adj_5309), 
          .C0(n177_adj_5760), .D0(n35_adj_4943), .A1(comb7_adj_6027[39]), 
          .B1(cout_adj_5309), .C1(n174_adj_5759), .D1(n34_adj_4942), .CIN(n15082), 
          .COUT(n15083), .S0(comb8_71__N_1595_adj_6054[38]), .S1(comb8_71__N_1595_adj_6054[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_3 (.A0(comb7_adj_6027[36]), .B0(cout_adj_5309), 
          .C0(n183_adj_5762), .D0(n37_adj_4945), .A1(comb7_adj_6027[37]), 
          .B1(cout_adj_5309), .C1(n180_adj_5761), .D1(n36_adj_4944), .CIN(n15081), 
          .COUT(n15082), .S0(comb8_71__N_1595_adj_6054[36]), .S1(comb8_71__N_1595_adj_6054[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1085_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1085_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1085_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_5309), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15081));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1085_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1085_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1085_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1085_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1028_add_4_15 (.A0(amdemod_d_11__N_2209), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15077), .S0(amdemod_d_11__N_1871[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1028_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1028_add_4_15.INIT1 = 16'h0000;
    defparam _add_1_1028_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1028_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1028_add_4_13 (.A0(amdemod_d_11__N_2215), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2212), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15076), .COUT(n15077), .S0(amdemod_d_11__N_1871[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1028_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1028_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1028_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1028_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1028_add_4_11 (.A0(amdemod_d_11__N_2221), .B0(n17162), 
          .C0(n17279), .D0(n17146), .A1(square_sum[23]), .B1(square_sum[22]), 
          .C1(amdemod_d_11__N_2218), .D1(VCC_net), .CIN(n15075), .COUT(n15076), 
          .S0(amdemod_d_11__N_1871[9]), .S1(amdemod_d_11__N_1871[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1028_add_4_11.INIT0 = 16'h596a;
    defparam _add_1_1028_add_4_11.INIT1 = 16'h1e1e;
    defparam _add_1_1028_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1028_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1028_add_4_9 (.A0(n17133), .B0(amdemod_d_11__N_2227), .C0(GND_net), 
          .D0(VCC_net), .A1(n17134), .B1(amdemod_d_11__N_2224), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15074), .COUT(n15075), .S0(amdemod_d_11__N_1871[7]), 
          .S1(amdemod_d_11__N_1871[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1028_add_4_9.INIT0 = 16'h9995;
    defparam _add_1_1028_add_4_9.INIT1 = 16'h9995;
    defparam _add_1_1028_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1028_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1028_add_4_7 (.A0(n17131), .B0(amdemod_d_11__N_2233), .C0(GND_net), 
          .D0(VCC_net), .A1(n17132), .B1(amdemod_d_11__N_2230), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15073), .COUT(n15074), .S0(amdemod_d_11__N_1871[5]), 
          .S1(amdemod_d_11__N_1871[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1028_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1028_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1028_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1028_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1028_add_4_5 (.A0(n17129), .B0(amdemod_d_11__N_2239), .C0(GND_net), 
          .D0(VCC_net), .A1(n17130), .B1(amdemod_d_11__N_2236), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15072), .COUT(n15073), .S0(amdemod_d_11__N_1871[3]), 
          .S1(amdemod_d_11__N_1871[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1028_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1028_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1028_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1028_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1028_add_4_3 (.A0(n17128), .B0(square_sum[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(n17128), .B1(amdemod_d_11__N_2242), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15071), .COUT(n15072), .S0(amdemod_d_11__N_1871[1]), 
          .S1(amdemod_d_11__N_1871[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1028_add_4_3.INIT0 = 16'h666a;
    defparam _add_1_1028_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1028_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1028_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1028_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15071), .S1(amdemod_d_11__N_1871[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1028_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1028_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1028_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1028_add_4_1.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_24 (.A0(n4_adj_5679), .B0(mult_result_i[22]), 
          .C0(GND_net), .D0(VCC_net), .A1(n2_adj_5678), .B1(mult_result_i[23]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15069), .S0(n55_adj_5703), 
          .S1(n52_adj_5702));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_add_4_24.INIT0 = 16'h666a;
    defparam square_sum_add_4_24.INIT1 = 16'h666a;
    defparam square_sum_add_4_24.INJECT1_0 = "NO";
    defparam square_sum_add_4_24.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_22 (.A0(n8_adj_5681), .B0(mult_result_i[20]), 
          .C0(GND_net), .D0(VCC_net), .A1(n6_adj_5680), .B1(mult_result_i[21]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15068), .COUT(n15069), .S0(n61_adj_5705), 
          .S1(n58_adj_5704));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_add_4_22.INIT0 = 16'h666a;
    defparam square_sum_add_4_22.INIT1 = 16'h666a;
    defparam square_sum_add_4_22.INJECT1_0 = "NO";
    defparam square_sum_add_4_22.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_20 (.A0(n12_adj_5683), .B0(mult_result_i[18]), 
          .C0(GND_net), .D0(VCC_net), .A1(n10_adj_5682), .B1(mult_result_i[19]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15067), .COUT(n15068), .S0(n67_adj_5707), 
          .S1(n64_adj_5706));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_add_4_20.INIT0 = 16'h666a;
    defparam square_sum_add_4_20.INIT1 = 16'h666a;
    defparam square_sum_add_4_20.INJECT1_0 = "NO";
    defparam square_sum_add_4_20.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_18 (.A0(n16_adj_5685), .B0(mult_result_i[16]), 
          .C0(GND_net), .D0(VCC_net), .A1(n14_adj_5684), .B1(mult_result_i[17]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15066), .COUT(n15067), .S0(n73_adj_5709), 
          .S1(n70_adj_5708));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_add_4_18.INIT0 = 16'h666a;
    defparam square_sum_add_4_18.INIT1 = 16'h666a;
    defparam square_sum_add_4_18.INJECT1_0 = "NO";
    defparam square_sum_add_4_18.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_16 (.A0(n20_adj_5687), .B0(mult_result_i[14]), 
          .C0(GND_net), .D0(VCC_net), .A1(n18_adj_5686), .B1(mult_result_i[15]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15065), .COUT(n15066), .S0(n79_adj_5711), 
          .S1(n76_adj_5710));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_add_4_16.INIT0 = 16'h666a;
    defparam square_sum_add_4_16.INIT1 = 16'h666a;
    defparam square_sum_add_4_16.INJECT1_0 = "NO";
    defparam square_sum_add_4_16.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_14 (.A0(n24_adj_5689), .B0(mult_result_i[12]), 
          .C0(GND_net), .D0(VCC_net), .A1(n22_adj_5688), .B1(mult_result_i[13]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15064), .COUT(n15065), .S0(n85_adj_5713), 
          .S1(n82_adj_5712));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_add_4_14.INIT0 = 16'h666a;
    defparam square_sum_add_4_14.INIT1 = 16'h666a;
    defparam square_sum_add_4_14.INJECT1_0 = "NO";
    defparam square_sum_add_4_14.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_12 (.A0(n28_adj_5691), .B0(mult_result_i[10]), 
          .C0(GND_net), .D0(VCC_net), .A1(n26_adj_5690), .B1(mult_result_i[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15063), .COUT(n15064), .S0(n91_adj_5715), 
          .S1(n88_adj_5714));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_add_4_12.INIT0 = 16'h666a;
    defparam square_sum_add_4_12.INIT1 = 16'h666a;
    defparam square_sum_add_4_12.INJECT1_0 = "NO";
    defparam square_sum_add_4_12.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_10 (.A0(n32_adj_5693), .B0(mult_result_i[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(n30_adj_5692), .B1(mult_result_i[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15062), .COUT(n15063), .S0(n97_adj_5717), 
          .S1(n94_adj_5716));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_add_4_10.INIT0 = 16'h666a;
    defparam square_sum_add_4_10.INIT1 = 16'h666a;
    defparam square_sum_add_4_10.INJECT1_0 = "NO";
    defparam square_sum_add_4_10.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_8 (.A0(n36_adj_5695), .B0(mult_result_i[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(n34_adj_5694), .B1(mult_result_i[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15061), .COUT(n15062), .S0(n103_adj_5719), 
          .S1(n100_adj_5718));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_add_4_8.INIT0 = 16'h666a;
    defparam square_sum_add_4_8.INIT1 = 16'h666a;
    defparam square_sum_add_4_8.INJECT1_0 = "NO";
    defparam square_sum_add_4_8.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_6 (.A0(n40_adj_5697), .B0(mult_result_i[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(n38_adj_5696), .B1(mult_result_i[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15060), .COUT(n15061), .S0(n109_adj_5721), 
          .S1(n106_adj_5720));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_add_4_6.INIT0 = 16'h666a;
    defparam square_sum_add_4_6.INIT1 = 16'h666a;
    defparam square_sum_add_4_6.INJECT1_0 = "NO";
    defparam square_sum_add_4_6.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_4 (.A0(n44_adj_5699), .B0(mult_result_i[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(n42_adj_5698), .B1(mult_result_i[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15059), .COUT(n15060), .S0(n115_adj_5723), 
          .S1(n112_adj_5722));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_add_4_4.INIT0 = 16'h666a;
    defparam square_sum_add_4_4.INIT1 = 16'h666a;
    defparam square_sum_add_4_4.INJECT1_0 = "NO";
    defparam square_sum_add_4_4.INJECT1_1 = "NO";
    CCU2C square_sum_add_4_2 (.A0(n48_adj_5701), .B0(mult_result_i[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(n46_adj_5700), .B1(mult_result_i[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15059), .S1(n118_adj_5724));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(90[22:51])
    defparam square_sum_add_4_2.INIT0 = 16'h0008;
    defparam square_sum_add_4_2.INIT1 = 16'h666a;
    defparam square_sum_add_4_2.INJECT1_0 = "NO";
    defparam square_sum_add_4_2.INJECT1_1 = "NO";
    LUT4 i2505_2_lut_2_lut (.A(n17289), .B(n292), .Z(n2102)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i2505_2_lut_2_lut.init = 16'hdddd;
    CCU2C _add_1_1034_add_4_13 (.A0(lo_sinewave[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15057), .S0(sinewave_out_11__N_236[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(48[23:35])
    defparam _add_1_1034_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_1034_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_1034_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_11 (.A0(lo_sinewave[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_sinewave[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15056), .COUT(n15057), .S0(sinewave_out_11__N_236[9]), 
          .S1(sinewave_out_11__N_236[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(48[23:35])
    defparam _add_1_1034_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_1034_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_1034_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_9 (.A0(lo_sinewave[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_sinewave[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15055), .COUT(n15056), .S0(sinewave_out_11__N_236[7]), 
          .S1(sinewave_out_11__N_236[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(48[23:35])
    defparam _add_1_1034_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_1034_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_1034_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_7 (.A0(lo_sinewave[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_sinewave[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15054), .COUT(n15055), .S0(sinewave_out_11__N_236[5]), 
          .S1(sinewave_out_11__N_236[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(48[23:35])
    defparam _add_1_1034_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_1034_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_1034_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_5 (.A0(lo_sinewave[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_sinewave[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15053), .COUT(n15054), .S0(sinewave_out_11__N_236[3]), 
          .S1(sinewave_out_11__N_236[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(48[23:35])
    defparam _add_1_1034_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_1034_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_1034_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_3 (.A0(lo_sinewave[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_sinewave[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15052), .COUT(n15053), .S0(sinewave_out_11__N_236[1]), 
          .S1(sinewave_out_11__N_236[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(48[23:35])
    defparam _add_1_1034_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_1034_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_1034_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1034_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_sinewave[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15052), .S1(sinewave_out_11__N_236[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(48[23:35])
    defparam _add_1_1034_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1034_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_1034_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1034_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_38 (.A0(comb_d7_adj_6028[71]), .B0(comb7_adj_6027[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15051), .S0(n78_adj_5727));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1145_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_36 (.A0(comb_d7_adj_6028[69]), .B0(comb7_adj_6027[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[70]), .B1(comb7_adj_6027[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15050), .COUT(n15051), .S0(n84_adj_5729), 
          .S1(n81_adj_5728));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_34 (.A0(comb_d7_adj_6028[67]), .B0(comb7_adj_6027[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[68]), .B1(comb7_adj_6027[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15049), .COUT(n15050), .S0(n90_adj_5731), 
          .S1(n87_adj_5730));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_32 (.A0(comb_d7_adj_6028[65]), .B0(comb7_adj_6027[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[66]), .B1(comb7_adj_6027[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15048), .COUT(n15049), .S0(n96_adj_5733), 
          .S1(n93_adj_5732));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_30 (.A0(comb_d7_adj_6028[63]), .B0(comb7_adj_6027[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[64]), .B1(comb7_adj_6027[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15047), .COUT(n15048), .S0(n102_adj_5735), 
          .S1(n99_adj_5734));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_28 (.A0(comb_d7_adj_6028[61]), .B0(comb7_adj_6027[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[62]), .B1(comb7_adj_6027[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15046), .COUT(n15047), .S0(n108_adj_5737), 
          .S1(n105_adj_5736));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_26 (.A0(comb_d7_adj_6028[59]), .B0(comb7_adj_6027[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[60]), .B1(comb7_adj_6027[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15045), .COUT(n15046), .S0(n114_adj_5739), 
          .S1(n111_adj_5738));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_24 (.A0(comb_d7_adj_6028[57]), .B0(comb7_adj_6027[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[58]), .B1(comb7_adj_6027[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15044), .COUT(n15045), .S0(n120_adj_5741), 
          .S1(n117_adj_5740));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_22 (.A0(comb_d7_adj_6028[55]), .B0(comb7_adj_6027[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[56]), .B1(comb7_adj_6027[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15043), .COUT(n15044), .S0(n126_adj_5743), 
          .S1(n123_adj_5742));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_20 (.A0(comb_d7_adj_6028[53]), .B0(comb7_adj_6027[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[54]), .B1(comb7_adj_6027[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15042), .COUT(n15043), .S0(n132_adj_5745), 
          .S1(n129_adj_5744));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_18 (.A0(comb_d7_adj_6028[51]), .B0(comb7_adj_6027[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[52]), .B1(comb7_adj_6027[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15041), .COUT(n15042), .S0(n138_adj_5747), 
          .S1(n135_adj_5746));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_16 (.A0(comb_d7_adj_6028[49]), .B0(comb7_adj_6027[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[50]), .B1(comb7_adj_6027[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15040), .COUT(n15041), .S0(n144_adj_5749), 
          .S1(n141_adj_5748));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_14 (.A0(comb_d7_adj_6028[47]), .B0(comb7_adj_6027[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[48]), .B1(comb7_adj_6027[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15039), .COUT(n15040), .S0(n150_adj_5751), 
          .S1(n147_adj_5750));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_12 (.A0(comb_d7_adj_6028[45]), .B0(comb7_adj_6027[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[46]), .B1(comb7_adj_6027[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15038), .COUT(n15039), .S0(n156_adj_5753), 
          .S1(n153_adj_5752));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_10 (.A0(comb_d7_adj_6028[43]), .B0(comb7_adj_6027[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[44]), .B1(comb7_adj_6027[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15037), .COUT(n15038), .S0(n162_adj_5755), 
          .S1(n159_adj_5754));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_8 (.A0(comb_d7_adj_6028[41]), .B0(comb7_adj_6027[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[42]), .B1(comb7_adj_6027[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15036), .COUT(n15037), .S0(n168_adj_5757), 
          .S1(n165_adj_5756));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_6 (.A0(comb_d7_adj_6028[39]), .B0(comb7_adj_6027[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[40]), .B1(comb7_adj_6027[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15035), .COUT(n15036), .S0(n174_adj_5759), 
          .S1(n171_adj_5758));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_4 (.A0(comb_d7_adj_6028[37]), .B0(comb7_adj_6027[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d7_adj_6028[38]), .B1(comb7_adj_6027[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15034), .COUT(n15035), .S0(n180_adj_5761), 
          .S1(n177_adj_5760));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1145_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1145_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d7_adj_6028[36]), .B1(comb7_adj_6027[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15034), .S1(n183_adj_5762));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1145_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1145_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1145_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1145_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1037_add_4_13 (.A0(lo_cosinewave[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15033), .S0(cosinewave_out_11__N_250[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(49[25:39])
    defparam _add_1_1037_add_4_13.INIT0 = 16'h5555;
    defparam _add_1_1037_add_4_13.INIT1 = 16'h0000;
    defparam _add_1_1037_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1037_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1037_add_4_11 (.A0(lo_cosinewave[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_cosinewave[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15032), .COUT(n15033), .S0(cosinewave_out_11__N_250[9]), 
          .S1(cosinewave_out_11__N_250[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(49[25:39])
    defparam _add_1_1037_add_4_11.INIT0 = 16'h5555;
    defparam _add_1_1037_add_4_11.INIT1 = 16'h5555;
    defparam _add_1_1037_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1037_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1037_add_4_9 (.A0(lo_cosinewave[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_cosinewave[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15031), .COUT(n15032), .S0(cosinewave_out_11__N_250[7]), 
          .S1(cosinewave_out_11__N_250[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(49[25:39])
    defparam _add_1_1037_add_4_9.INIT0 = 16'h5555;
    defparam _add_1_1037_add_4_9.INIT1 = 16'h5555;
    defparam _add_1_1037_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1037_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1037_add_4_7 (.A0(lo_cosinewave[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_cosinewave[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15030), .COUT(n15031), .S0(cosinewave_out_11__N_250[5]), 
          .S1(cosinewave_out_11__N_250[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(49[25:39])
    defparam _add_1_1037_add_4_7.INIT0 = 16'h5555;
    defparam _add_1_1037_add_4_7.INIT1 = 16'h5555;
    defparam _add_1_1037_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1037_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1037_add_4_5 (.A0(lo_cosinewave[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_cosinewave[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15029), .COUT(n15030), .S0(cosinewave_out_11__N_250[3]), 
          .S1(cosinewave_out_11__N_250[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(49[25:39])
    defparam _add_1_1037_add_4_5.INIT0 = 16'h5555;
    defparam _add_1_1037_add_4_5.INIT1 = 16'h5555;
    defparam _add_1_1037_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1037_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1037_add_4_3 (.A0(lo_cosinewave[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_cosinewave[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15028), .COUT(n15029), .S0(cosinewave_out_11__N_250[1]), 
          .S1(cosinewave_out_11__N_250[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(49[25:39])
    defparam _add_1_1037_add_4_3.INIT0 = 16'h5555;
    defparam _add_1_1037_add_4_3.INIT1 = 16'h5555;
    defparam _add_1_1037_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1037_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1037_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(lo_cosinewave[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15028), .S1(cosinewave_out_11__N_250[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(49[25:39])
    defparam _add_1_1037_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1037_add_4_1.INIT1 = 16'haaa5;
    defparam _add_1_1037_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1037_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_38 (.A0(comb_d6_adj_6026[71]), .B0(comb6_adj_6025[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15027), .S0(n78_adj_5763));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1148_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_36 (.A0(comb_d6_adj_6026[69]), .B0(comb6_adj_6025[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[70]), .B1(comb6_adj_6025[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15026), .COUT(n15027), .S0(n84_adj_5765), 
          .S1(n81_adj_5764));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_34 (.A0(comb_d6_adj_6026[67]), .B0(comb6_adj_6025[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[68]), .B1(comb6_adj_6025[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15025), .COUT(n15026), .S0(n90_adj_5767), 
          .S1(n87_adj_5766));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_32 (.A0(comb_d6_adj_6026[65]), .B0(comb6_adj_6025[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[66]), .B1(comb6_adj_6025[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15024), .COUT(n15025), .S0(n96_adj_5769), 
          .S1(n93_adj_5768));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_30 (.A0(comb_d6_adj_6026[63]), .B0(comb6_adj_6025[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[64]), .B1(comb6_adj_6025[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15023), .COUT(n15024), .S0(n102_adj_5771), 
          .S1(n99_adj_5770));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_28 (.A0(comb_d6_adj_6026[61]), .B0(comb6_adj_6025[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[62]), .B1(comb6_adj_6025[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15022), .COUT(n15023), .S0(n108_adj_5773), 
          .S1(n105_adj_5772));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_26 (.A0(comb_d6_adj_6026[59]), .B0(comb6_adj_6025[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[60]), .B1(comb6_adj_6025[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15021), .COUT(n15022), .S0(n114_adj_5775), 
          .S1(n111_adj_5774));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_24 (.A0(comb_d6_adj_6026[57]), .B0(comb6_adj_6025[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[58]), .B1(comb6_adj_6025[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15020), .COUT(n15021), .S0(n120_adj_5777), 
          .S1(n117_adj_5776));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_22 (.A0(comb_d6_adj_6026[55]), .B0(comb6_adj_6025[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[56]), .B1(comb6_adj_6025[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15019), .COUT(n15020), .S0(n126_adj_5779), 
          .S1(n123_adj_5778));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_20 (.A0(comb_d6_adj_6026[53]), .B0(comb6_adj_6025[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[54]), .B1(comb6_adj_6025[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15018), .COUT(n15019), .S0(n132_adj_5781), 
          .S1(n129_adj_5780));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_18 (.A0(comb_d6_adj_6026[51]), .B0(comb6_adj_6025[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[52]), .B1(comb6_adj_6025[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15017), .COUT(n15018), .S0(n138_adj_5783), 
          .S1(n135_adj_5782));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_16 (.A0(comb_d6_adj_6026[49]), .B0(comb6_adj_6025[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[50]), .B1(comb6_adj_6025[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15016), .COUT(n15017), .S0(n144_adj_5785), 
          .S1(n141_adj_5784));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_14 (.A0(comb_d6_adj_6026[47]), .B0(comb6_adj_6025[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[48]), .B1(comb6_adj_6025[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15015), .COUT(n15016), .S0(n150_adj_5787), 
          .S1(n147_adj_5786));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_12 (.A0(comb_d6_adj_6026[45]), .B0(comb6_adj_6025[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[46]), .B1(comb6_adj_6025[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15014), .COUT(n15015), .S0(n156_adj_5789), 
          .S1(n153_adj_5788));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_10 (.A0(comb_d6_adj_6026[43]), .B0(comb6_adj_6025[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[44]), .B1(comb6_adj_6025[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15013), .COUT(n15014), .S0(n162_adj_5791), 
          .S1(n159_adj_5790));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_8 (.A0(comb_d6_adj_6026[41]), .B0(comb6_adj_6025[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[42]), .B1(comb6_adj_6025[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15012), .COUT(n15013), .S0(n168_adj_5793), 
          .S1(n165_adj_5792));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_6 (.A0(comb_d6_adj_6026[39]), .B0(comb6_adj_6025[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[40]), .B1(comb6_adj_6025[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15011), .COUT(n15012), .S0(n174_adj_5795), 
          .S1(n171_adj_5794));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_4 (.A0(comb_d6_adj_6026[37]), .B0(comb6_adj_6025[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d6_adj_6026[38]), .B1(comb6_adj_6025[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15010), .COUT(n15011), .S0(n180_adj_5797), 
          .S1(n177_adj_5796));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1148_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1148_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d6_adj_6026[36]), .B1(comb6_adj_6025[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15010), .S1(n183_adj_5798));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam _add_1_1148_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1148_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1148_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1148_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_37 (.A0(integrator3_adj_6022[70]), .B0(cout_adj_5165), 
          .C0(n81_adj_5499), .D0(integrator4_adj_6023[70]), .A1(integrator3_adj_6022[71]), 
          .B1(cout_adj_5165), .C1(n78_adj_5498), .D1(integrator4_adj_6023[71]), 
          .CIN(n15008), .S0(integrator4_71__N_634_adj_6039[70]), .S1(integrator4_71__N_634_adj_6039[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_35 (.A0(integrator3_adj_6022[68]), .B0(cout_adj_5165), 
          .C0(n87_adj_5501), .D0(integrator4_adj_6023[68]), .A1(integrator3_adj_6022[69]), 
          .B1(cout_adj_5165), .C1(n84_adj_5500), .D1(integrator4_adj_6023[69]), 
          .CIN(n15007), .COUT(n15008), .S0(integrator4_71__N_634_adj_6039[68]), 
          .S1(integrator4_71__N_634_adj_6039[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_33 (.A0(integrator3_adj_6022[66]), .B0(cout_adj_5165), 
          .C0(n93_adj_5503), .D0(integrator4_adj_6023[66]), .A1(integrator3_adj_6022[67]), 
          .B1(cout_adj_5165), .C1(n90_adj_5502), .D1(integrator4_adj_6023[67]), 
          .CIN(n15006), .COUT(n15007), .S0(integrator4_71__N_634_adj_6039[66]), 
          .S1(integrator4_71__N_634_adj_6039[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_31 (.A0(integrator3_adj_6022[64]), .B0(cout_adj_5165), 
          .C0(n99_adj_5505), .D0(integrator4_adj_6023[64]), .A1(integrator3_adj_6022[65]), 
          .B1(cout_adj_5165), .C1(n96_adj_5504), .D1(integrator4_adj_6023[65]), 
          .CIN(n15005), .COUT(n15006), .S0(integrator4_71__N_634_adj_6039[64]), 
          .S1(integrator4_71__N_634_adj_6039[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_29 (.A0(integrator3_adj_6022[62]), .B0(cout_adj_5165), 
          .C0(n105_adj_5507), .D0(integrator4_adj_6023[62]), .A1(integrator3_adj_6022[63]), 
          .B1(cout_adj_5165), .C1(n102_adj_5506), .D1(integrator4_adj_6023[63]), 
          .CIN(n15004), .COUT(n15005), .S0(integrator4_71__N_634_adj_6039[62]), 
          .S1(integrator4_71__N_634_adj_6039[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_27 (.A0(integrator3_adj_6022[60]), .B0(cout_adj_5165), 
          .C0(n111_adj_5509), .D0(integrator4_adj_6023[60]), .A1(integrator3_adj_6022[61]), 
          .B1(cout_adj_5165), .C1(n108_adj_5508), .D1(integrator4_adj_6023[61]), 
          .CIN(n15003), .COUT(n15004), .S0(integrator4_71__N_634_adj_6039[60]), 
          .S1(integrator4_71__N_634_adj_6039[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_25 (.A0(integrator3_adj_6022[58]), .B0(cout_adj_5165), 
          .C0(n117_adj_5511), .D0(integrator4_adj_6023[58]), .A1(integrator3_adj_6022[59]), 
          .B1(cout_adj_5165), .C1(n114_adj_5510), .D1(integrator4_adj_6023[59]), 
          .CIN(n15002), .COUT(n15003), .S0(integrator4_71__N_634_adj_6039[58]), 
          .S1(integrator4_71__N_634_adj_6039[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_23 (.A0(integrator3_adj_6022[56]), .B0(cout_adj_5165), 
          .C0(n123_adj_5513), .D0(integrator4_adj_6023[56]), .A1(integrator3_adj_6022[57]), 
          .B1(cout_adj_5165), .C1(n120_adj_5512), .D1(integrator4_adj_6023[57]), 
          .CIN(n15001), .COUT(n15002), .S0(integrator4_71__N_634_adj_6039[56]), 
          .S1(integrator4_71__N_634_adj_6039[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_21 (.A0(integrator3_adj_6022[54]), .B0(cout_adj_5165), 
          .C0(n129_adj_5515), .D0(integrator4_adj_6023[54]), .A1(integrator3_adj_6022[55]), 
          .B1(cout_adj_5165), .C1(n126_adj_5514), .D1(integrator4_adj_6023[55]), 
          .CIN(n15000), .COUT(n15001), .S0(integrator4_71__N_634_adj_6039[54]), 
          .S1(integrator4_71__N_634_adj_6039[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_19 (.A0(integrator3_adj_6022[52]), .B0(cout_adj_5165), 
          .C0(n135_adj_5517), .D0(integrator4_adj_6023[52]), .A1(integrator3_adj_6022[53]), 
          .B1(cout_adj_5165), .C1(n132_adj_5516), .D1(integrator4_adj_6023[53]), 
          .CIN(n14999), .COUT(n15000), .S0(integrator4_71__N_634_adj_6039[52]), 
          .S1(integrator4_71__N_634_adj_6039[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_17 (.A0(integrator3_adj_6022[50]), .B0(cout_adj_5165), 
          .C0(n141_adj_5519), .D0(integrator4_adj_6023[50]), .A1(integrator3_adj_6022[51]), 
          .B1(cout_adj_5165), .C1(n138_adj_5518), .D1(integrator4_adj_6023[51]), 
          .CIN(n14998), .COUT(n14999), .S0(integrator4_71__N_634_adj_6039[50]), 
          .S1(integrator4_71__N_634_adj_6039[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_15 (.A0(integrator3_adj_6022[48]), .B0(cout_adj_5165), 
          .C0(n147_adj_5521), .D0(integrator4_adj_6023[48]), .A1(integrator3_adj_6022[49]), 
          .B1(cout_adj_5165), .C1(n144_adj_5520), .D1(integrator4_adj_6023[49]), 
          .CIN(n14997), .COUT(n14998), .S0(integrator4_71__N_634_adj_6039[48]), 
          .S1(integrator4_71__N_634_adj_6039[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_13 (.A0(integrator3_adj_6022[46]), .B0(cout_adj_5165), 
          .C0(n153_adj_5523), .D0(integrator4_adj_6023[46]), .A1(integrator3_adj_6022[47]), 
          .B1(cout_adj_5165), .C1(n150_adj_5522), .D1(integrator4_adj_6023[47]), 
          .CIN(n14996), .COUT(n14997), .S0(integrator4_71__N_634_adj_6039[46]), 
          .S1(integrator4_71__N_634_adj_6039[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_11 (.A0(integrator3_adj_6022[44]), .B0(cout_adj_5165), 
          .C0(n159_adj_5525), .D0(integrator4_adj_6023[44]), .A1(integrator3_adj_6022[45]), 
          .B1(cout_adj_5165), .C1(n156_adj_5524), .D1(integrator4_adj_6023[45]), 
          .CIN(n14995), .COUT(n14996), .S0(integrator4_71__N_634_adj_6039[44]), 
          .S1(integrator4_71__N_634_adj_6039[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1097_add_4_9 (.A0(integrator3_adj_6022[42]), .B0(cout_adj_5165), 
          .C0(n165_adj_5527), .D0(integrator4_adj_6023[42]), .A1(integrator3_adj_6022[43]), 
          .B1(cout_adj_5165), .C1(n162_adj_5526), .D1(integrator4_adj_6023[43]), 
          .CIN(n14994), .COUT(n14995), .S0(integrator4_71__N_634_adj_6039[42]), 
          .S1(integrator4_71__N_634_adj_6039[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(69[20:45])
    defparam _add_1_1097_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1097_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1097_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1097_add_4_9.INJECT1_1 = "NO";
    LUT4 i1629_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(led_c_3), .D(n214), 
         .Z(n11351)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1629_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1605_3_lut_4_lut (.A(n17288), .B(n17150), .C(led_c_3), .D(n253), 
         .Z(n11327)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1605_3_lut_4_lut.init = 16'hf707;
    LUT4 mux_251_i25_4_lut (.A(n11333), .B(n247_adj_5943), .C(n17136), 
         .D(n2244), .Z(n2020)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i25_4_lut.init = 16'hc0ca;
    LUT4 i4701_2_lut (.A(integrator1_adj_6020[0]), .B(mix_cosinewave[0]), 
         .Z(integrator1_71__N_418_adj_6036[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4701_2_lut.init = 16'h6666;
    LUT4 i4694_2_lut (.A(n48_adj_5701), .B(mult_result_i[0]), .Z(n121)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4694_2_lut.init = 16'h6666;
    VLO i1 (.Z(GND_net));
    LUT4 i1595_3_lut_4_lut (.A(n17288), .B(n17150), .C(n17289), .D(n271), 
         .Z(n11317)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1595_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_251_i26_4_lut (.A(n11335), .B(n244_adj_5942), .C(n17136), 
         .D(n2244), .Z(n2019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i26_4_lut.init = 16'hcfca;
    LUT4 i26_4_lut_adj_200 (.A(n2244), .B(n253_adj_5945), .C(n17136), 
         .D(n13_adj_4747), .Z(n11_adj_4729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i26_4_lut_adj_200.init = 16'hcacf;
    LUT4 mux_251_i24_4_lut (.A(n11331), .B(n250_adj_5944), .C(n17136), 
         .D(n2244), .Z(n2021)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i24_4_lut.init = 16'hcfca;
    LUT4 mux_251_i21_4_lut (.A(n11327), .B(n259_adj_5947), .C(n17136), 
         .D(n2244), .Z(n2024)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i21_4_lut.init = 16'hcfca;
    LUT4 i1585_3_lut_4_lut (.A(n17288), .B(n17150), .C(led_c_3), .D(n289), 
         .Z(n11307)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1585_3_lut_4_lut.init = 16'hf808;
    LUT4 i4697_2_lut (.A(integrator2_adj_6021[0]), .B(integrator1_adj_6020[0]), 
         .Z(integrator2_71__N_490_adj_6037[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4697_2_lut.init = 16'h6666;
    LUT4 i1587_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(n17289), .D(n286), 
         .Z(n11309)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1587_3_lut_4_lut.init = 16'hf707;
    LUT4 i1581_3_lut_4_lut (.A(n17288), .B(n17150), .C(n17289), .D(n298), 
         .Z(n11303)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1581_3_lut_4_lut.init = 16'hf808;
    LUT4 i4727_4_lut (.A(n16451), .B(n17153), .C(n17049), .D(n16957), 
         .Z(clk_80mhz_enable_1507)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C))) */ ;
    defparam i4727_4_lut.init = 16'hc0c8;
    LUT4 i2424_rep_269_2_lut (.A(led_c_2), .B(led_c_1), .Z(n16957)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2424_rep_269_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_201 (.A(n17043), .B(n17149), .C(n11789), .D(n16245), 
         .Z(n16409)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_201.init = 16'ha080;
    LUT4 i2_2_lut_3_lut_3_lut (.A(led_c_3), .B(n17150), .C(led_c_2), .Z(n15867)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i2_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 i4689_2_lut (.A(integrator3_adj_6022[0]), .B(integrator2_adj_6021[0]), 
         .Z(integrator3_71__N_562_adj_6038[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4689_2_lut.init = 16'h6666;
    LUT4 i1878_4_lut (.A(n256_adj_5946), .B(n250), .C(led_c_3), .D(n17144), 
         .Z(n11612)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1878_4_lut.init = 16'hcac0;
    LUT4 i4688_2_lut (.A(integrator4_adj_6023[0]), .B(integrator3_adj_6022[0]), 
         .Z(integrator4_71__N_634_adj_6039[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4688_2_lut.init = 16'h6666;
    LUT4 mux_251_i19_4_lut (.A(n11323), .B(n265_adj_5949), .C(n17136), 
         .D(n2244), .Z(n2026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i19_4_lut.init = 16'hcfca;
    LUT4 i284_2_lut_3_lut_3_lut (.A(led_c_3), .B(n16220), .C(led_c_4), 
         .Z(n2244)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i284_2_lut_3_lut_3_lut.init = 16'h0404;
    LUT4 i1876_4_lut (.A(n262_adj_5948), .B(n256), .C(led_c_3), .D(n17144), 
         .Z(n11610)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1876_4_lut.init = 16'hcac0;
    LUT4 mux_251_i17_4_lut (.A(n11319), .B(n271_adj_5951), .C(n17136), 
         .D(n2244), .Z(n2028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i17_4_lut.init = 16'hcfca;
    LUT4 mux_251_i51_4_lut (.A(n2193), .B(n169_adj_5917), .C(n17136), 
         .D(n2244), .Z(n1994)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i51_4_lut.init = 16'hcfca;
    LUT4 i4687_2_lut (.A(integrator5_adj_6024[0]), .B(integrator4_adj_6023[0]), 
         .Z(integrator5_71__N_706_adj_6040[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4687_2_lut.init = 16'h6666;
    LUT4 i1_3_lut_4_lut_4_lut_adj_202 (.A(led_c_1), .B(led_c_2), .C(led_c_3), 
         .D(n17149), .Z(n16203)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_202.init = 16'hfff7;
    LUT4 i2543_2_lut (.A(n163), .B(n17289), .Z(n2193)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i2543_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_4_lut_4_lut_4_lut (.A(led_c_1), .B(led_c_0), .C(led_c_4), 
         .D(led_c_3), .Z(n16388)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_4_lut_4_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_342_3_lut_4_lut_4_lut (.A(led_c_1), .B(led_c_4), .C(n17155), 
         .D(led_c_6), .Z(n17139)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;
    defparam i1_2_lut_rep_342_3_lut_4_lut_4_lut.init = 16'hdfff;
    LUT4 i1675_3_lut_4_lut (.A(n17288), .B(n17150), .C(n17289), .D(n133), 
         .Z(n11397)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1675_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i4705_2_lut (.A(integrator2[0]), .B(integrator1[0]), .Z(integrator2_71__N_490[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4705_2_lut.init = 16'h6666;
    LUT4 mux_366_i22_3_lut (.A(led_c_2), .B(led_c_4), .C(n1827), .Z(n2559)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_366_i22_3_lut.init = 16'h3a3a;
    LUT4 mux_251_i52_4_lut (.A(n11381), .B(n166_adj_5916), .C(n17136), 
         .D(n2244), .Z(n1993)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i52_4_lut.init = 16'hcfca;
    LUT4 mux_251_i18_4_lut (.A(n2226), .B(n268_adj_5950), .C(n17136), 
         .D(n2244), .Z(n2027)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i18_4_lut.init = 16'hcfca;
    LUT4 i2532_2_lut (.A(n262), .B(n17289), .Z(n2226)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i2532_2_lut.init = 16'h8888;
    LUT4 mux_251_i15_4_lut (.A(n11317), .B(n277_adj_5953), .C(n17136), 
         .D(n2244), .Z(n2030)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i15_4_lut.init = 16'hcfca;
    LUT4 i1671_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(led_c_3), .D(n139), 
         .Z(n11393)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1671_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_251_i16_4_lut (.A(n2094), .B(n274_adj_5952), .C(n17136), 
         .D(n11259), .Z(n2029)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i16_4_lut.init = 16'hc0ca;
    LUT4 mux_251_i13_4_lut (.A(n2097), .B(n283_adj_5955), .C(n17136), 
         .D(n11259), .Z(n2032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i13_4_lut.init = 16'hcfca;
    LUT4 i2506_2_lut (.A(n277), .B(led_c_3), .Z(n2097)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i2506_2_lut.init = 16'h8888;
    Mixer mixer_inst (.mix_sinewave({mix_sinewave}), .clk_80mhz(clk_80mhz), 
          .diff_out_c(diff_out_c), .mix_cosinewave({mix_cosinewave}), .rf_in_c(rf_in_c), 
          .\lo_cosinewave[10] (lo_cosinewave[10]), .cosinewave_out_11__N_250({cosinewave_out_11__N_250}), 
          .\lo_sinewave[4] (lo_sinewave[4]), .sinewave_out_11__N_236({sinewave_out_11__N_236}), 
          .\lo_cosinewave[11] (lo_cosinewave[11]), .\lo_sinewave[5] (lo_sinewave[5]), 
          .\lo_sinewave[6] (lo_sinewave[6]), .\lo_cosinewave[1] (lo_cosinewave[1]), 
          .\lo_sinewave[7] (lo_sinewave[7]), .\lo_sinewave[8] (lo_sinewave[8]), 
          .\lo_sinewave[9] (lo_sinewave[9]), .\lo_sinewave[10] (lo_sinewave[10]), 
          .\lo_sinewave[11] (lo_sinewave[11]), .\lo_sinewave[12] (lo_sinewave[12]), 
          .\lo_cosinewave[2] (lo_cosinewave[2]), .\lo_cosinewave[3] (lo_cosinewave[3]), 
          .\lo_cosinewave[4] (lo_cosinewave[4]), .\lo_cosinewave[5] (lo_cosinewave[5]), 
          .\lo_cosinewave[6] (lo_cosinewave[6]), .\lo_cosinewave[12] (lo_cosinewave[12]), 
          .\lo_cosinewave[7] (lo_cosinewave[7]), .\lo_cosinewave[8] (lo_cosinewave[8]), 
          .\lo_sinewave[2] (lo_sinewave[2]), .\lo_sinewave[1] (lo_sinewave[1]), 
          .\lo_cosinewave[9] (lo_cosinewave[9]), .\lo_sinewave[3] (lo_sinewave[3])) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(137[7] 145[6])
    LUT4 mux_251_i14_4_lut (.A(n2230), .B(n280_adj_5954), .C(n17136), 
         .D(n2244), .Z(n2031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i14_4_lut.init = 16'hcfca;
    LUT4 i1615_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(n17289), .D(n235), 
         .Z(n11337)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1615_3_lut_4_lut.init = 16'hf808;
    LUT4 i2528_2_lut (.A(n274), .B(n17289), .Z(n2230)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i2528_2_lut.init = 16'h8888;
    LUT4 pwm_out_I_0_1_lut (.A(pwm_out_p4_c), .Z(pwm_out_n4_c)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(229[25:33])
    defparam pwm_out_I_0_1_lut.init = 16'h5555;
    LUT4 i1673_3_lut_4_lut (.A(n17288), .B(n17150), .C(n17289), .D(n136), 
         .Z(n11395)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1673_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_251_i27_4_lut (.A(n11337), .B(n241_adj_5941), .C(n17136), 
         .D(n2244), .Z(n2018)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i27_4_lut.init = 16'hc0ca;
    LUT4 mux_251_i49_4_lut (.A(n11377), .B(n175_adj_5919), .C(n17136), 
         .D(n2244), .Z(n1996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i49_4_lut.init = 16'hcfca;
    LUT4 mux_251_i11_4_lut (.A(n11311), .B(n289_adj_5957), .C(n17136), 
         .D(n2244), .Z(n2034)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i11_4_lut.init = 16'hc0ca;
    LUT4 i1665_3_lut_4_lut (.A(n17288), .B(n17150), .C(led_c_3), .D(n151), 
         .Z(n11387)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1665_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1617_3_lut_4_lut (.A(n17288), .B(n17150), .C(led_c_3), .D(n232), 
         .Z(n11339)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1617_3_lut_4_lut.init = 16'hf707;
    LUT4 mux_251_i50_4_lut (.A(n2060), .B(n172_adj_5918), .C(n17136), 
         .D(n11259), .Z(n1995)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i50_4_lut.init = 16'hcfca;
    LUT4 i1653_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(led_c_3), .D(n172), 
         .Z(n11375)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1653_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1647_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(n17289), .D(n184), 
         .Z(n11369)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1647_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i2511_2_lut (.A(n166), .B(led_c_3), .Z(n2060)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i2511_2_lut.init = 16'h8888;
    LUT4 mux_251_i28_4_lut (.A(n11339), .B(n238_adj_5940), .C(n17136), 
         .D(n2244), .Z(n2017)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i28_4_lut.init = 16'hc0ca;
    LUT4 i1613_3_lut_4_lut (.A(n17288), .B(n17150), .C(n17289), .D(n238), 
         .Z(n11335)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1613_3_lut_4_lut.init = 16'hf808;
    LUT4 i1627_3_lut_4_lut (.A(n17288), .B(n17150), .C(n17289), .D(n217), 
         .Z(n11349)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1627_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_251_i10_4_lut (.A(n11309), .B(n292_adj_5958), .C(n17136), 
         .D(n2244), .Z(n2035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i10_4_lut.init = 16'hcfca;
    LUT4 mux_251_i7_4_lut (.A(n2237), .B(n301_adj_5961), .C(n17136), .D(n2244), 
         .Z(n2038)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i7_4_lut.init = 16'hc0ca;
    LUT4 mux_251_i8_4_lut (.A(n2102), .B(n298_adj_5960), .C(n17136), .D(n11259), 
         .Z(n2037)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i8_4_lut.init = 16'hc0ca;
    LUT4 i1611_3_lut_4_lut (.A(led_c_2), .B(n17150), .C(led_c_3), .D(n241), 
         .Z(n11333)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1611_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_251_i5_4_lut (.A(n11301), .B(n307), .C(n17136), .D(n2244), 
         .Z(n2040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i5_4_lut.init = 16'hcfca;
    LUT4 mux_251_i6_4_lut (.A(n11303), .B(n304), .C(n17136), .D(n2244), 
         .Z(n2039)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam mux_251_i6_4_lut.init = 16'hc0ca;
    LUT4 i1601_3_lut_4_lut (.A(n17288), .B(n17150), .C(led_c_3), .D(n259), 
         .Z(n11323)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(239[9] 259[12])
    defparam i1601_3_lut_4_lut.init = 16'hfb0b;
    FD1P3AX phase_inc_gen_i0_i2 (.D(n317), .SP(clk_80mhz_enable_1447), .CK(clk_80mhz), 
            .Q(phase_inc_gen[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i2.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i3 (.D(n314), .SP(clk_80mhz_enable_1447), .CK(clk_80mhz), 
            .Q(phase_inc_gen[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i3.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i4 (.D(n311), .SP(clk_80mhz_enable_1497), .CK(clk_80mhz), 
            .Q(phase_inc_gen[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i4.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i5 (.D(n308), .SP(clk_80mhz_enable_1497), .CK(clk_80mhz), 
            .Q(phase_inc_gen[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i5.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i6 (.D(n305), .SP(clk_80mhz_enable_1497), .CK(clk_80mhz), 
            .Q(phase_inc_gen[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i6.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i7 (.D(n302), .SP(clk_80mhz_enable_1497), .CK(clk_80mhz), 
            .Q(phase_inc_gen[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i7.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i8 (.D(n299), .SP(clk_80mhz_enable_1497), .CK(clk_80mhz), 
            .Q(phase_inc_gen[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i8.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i9 (.D(n296), .SP(clk_80mhz_enable_1497), .CK(clk_80mhz), 
            .Q(phase_inc_gen[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i9.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i10 (.D(n293), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i10.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i11 (.D(n290), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i11.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i12 (.D(n287), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i12.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i13 (.D(n284), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i13.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i14 (.D(n281), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i14.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i15 (.D(n278), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i15.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i16 (.D(n275), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[16]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i16.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i17 (.D(n272), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[17]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i17.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i18 (.D(n269), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[18]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i18.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i19 (.D(n266), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[19]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i19.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i20 (.D(n263), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[20]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i20.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i21 (.D(n260), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i21.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i22 (.D(n257), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[22]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i22.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i23 (.D(n254), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i23.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i24 (.D(n251), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[24]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i24.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i25 (.D(n248), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i25.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i26 (.D(n245), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[26]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i26.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i27 (.D(n242), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i27.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i28 (.D(n239), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[28]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i28.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i29 (.D(n236), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i29.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i30 (.D(n233), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[30]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i30.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i31 (.D(n230), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i31.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i32 (.D(n227), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[32]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i32.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i33 (.D(n224), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i33.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i34 (.D(n221), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[34]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i34.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i35 (.D(n218), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i35.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i36 (.D(n215), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[36]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i36.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i37 (.D(n212), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i37.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i38 (.D(n209), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[38]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i38.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i39 (.D(n206), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i39.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i40 (.D(n203), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[40]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i40.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i41 (.D(n200), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i41.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i42 (.D(n197), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[42]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i42.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i43 (.D(n194), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i43.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i44 (.D(n191), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[44]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i44.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i45 (.D(n188), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i45.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i46 (.D(n185), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[46]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i46.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i47 (.D(n182), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i47.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i48 (.D(n179), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[48]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i48.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i49 (.D(n176), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i49.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i50 (.D(n173), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[50]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i50.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i51 (.D(n170), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i51.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i52 (.D(n167), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[52]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i52.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i53 (.D(n164), .SP(clk_80mhz_enable_1497), 
            .CK(clk_80mhz), .Q(phase_inc_gen[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i53.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i54 (.D(n161), .SP(clk_80mhz_enable_1507), 
            .CK(clk_80mhz), .Q(phase_inc_gen[54]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i54.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i55 (.D(n158), .SP(clk_80mhz_enable_1507), 
            .CK(clk_80mhz), .Q(phase_inc_gen[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i55.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i56 (.D(n155), .SP(clk_80mhz_enable_1507), 
            .CK(clk_80mhz), .Q(phase_inc_gen[56]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i56.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i57 (.D(n152), .SP(clk_80mhz_enable_1507), 
            .CK(clk_80mhz), .Q(phase_inc_gen[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i57.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i58 (.D(n149), .SP(clk_80mhz_enable_1507), 
            .CK(clk_80mhz), .Q(phase_inc_gen[58]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i58.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i59 (.D(n146), .SP(clk_80mhz_enable_1507), 
            .CK(clk_80mhz), .Q(phase_inc_gen[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i59.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i60 (.D(n143), .SP(clk_80mhz_enable_1507), 
            .CK(clk_80mhz), .Q(phase_inc_gen[60]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i60.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i61 (.D(n140), .SP(clk_80mhz_enable_1507), 
            .CK(clk_80mhz), .Q(phase_inc_gen[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i61.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i62 (.D(n137), .SP(clk_80mhz_enable_1507), 
            .CK(clk_80mhz), .Q(phase_inc_gen[62]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i62.GSR = "ENABLED";
    FD1P3AX phase_inc_gen_i0_i63 (.D(n134), .SP(clk_80mhz_enable_1507), 
            .CK(clk_80mhz), .Q(phase_inc_gen[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam phase_inc_gen_i0_i63.GSR = "ENABLED";
    CCU2C _add_1_993_add_4_6 (.A0(integrator1_adj_6020[4]), .B0(mix_cosinewave[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[5]), .B1(mix_cosinewave[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15321), .COUT(n15322), .S0(integrator1_71__N_418_adj_6036[4]), 
          .S1(integrator1_71__N_418_adj_6036[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_61 (.A0(phase_inc_gen[63]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15675), .S0(n124));
    defparam _add_1_1241_add_4_61.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_61.INIT1 = 16'h0000;
    defparam _add_1_1241_add_4_61.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_61.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_59 (.A0(phase_inc_gen[61]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[62]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15674), .COUT(n15675), .S0(n130), .S1(n127));
    defparam _add_1_1241_add_4_59.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_59.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_59.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_59.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_347 (.A(led_c_4), .B(n16220), .Z(n17144)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam i1_2_lut_rep_347.init = 16'h8888;
    CCU2C _add_1_1241_add_4_57 (.A0(phase_inc_gen[59]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[60]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15673), .COUT(n15674), .S0(n136), .S1(n133));
    defparam _add_1_1241_add_4_57.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_57.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_57.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_57.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_55 (.A0(phase_inc_gen[57]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[58]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15672), .COUT(n15673), .S0(n142), .S1(n139));
    defparam _add_1_1241_add_4_55.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_55.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_55.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_55.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_53 (.A0(phase_inc_gen[55]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[56]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15671), .COUT(n15672), .S0(n148), .S1(n145));
    defparam _add_1_1241_add_4_53.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_53.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_53.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_53.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_18 (.A0(integrator_d_tmp[15]), .B0(integrator_tmp[15]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[16]), .B1(integrator_tmp[16]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15352), .COUT(n15353), .S0(comb6_71__N_1451[15]), 
          .S1(comb6_71__N_1451[16]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_10 (.A0(integrator3[43]), .B0(integrator2[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[44]), .B1(integrator2[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15552), .COUT(n15553), .S0(n162_adj_5339), 
          .S1(n159_adj_5338));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_14 (.A0(integrator_d_tmp[11]), .B0(integrator_tmp[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[12]), .B1(integrator_tmp[12]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15350), .COUT(n15351), .S0(comb6_71__N_1451[11]), 
          .S1(comb6_71__N_1451[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_51 (.A0(phase_inc_gen[53]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[54]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15670), .COUT(n15671), .S0(n154), .S1(n151));
    defparam _add_1_1241_add_4_51.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_51.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_51.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_51.INJECT1_1 = "NO";
    LUT4 i2538_3_lut (.A(led_c_0), .B(n11789), .C(n16203), .Z(n12278)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i2538_3_lut.init = 16'hc8c8;
    \CIC(REGISTER_WIDTH=72,DECIMATION_RATIO=4096)  cic_sine_inst (.integrator_d_tmp({integrator_d_tmp}), 
            .clk_80mhz(clk_80mhz), .integrator_tmp({integrator_tmp}), .n30(n30_adj_2970), 
            .integrator5({integrator5}), .integrator2({integrator2}), .integrator2_71__N_490({integrator2_71__N_490}), 
            .n33(n33_adj_2967), .integrator3({integrator3}), .integrator3_71__N_562({integrator3_71__N_562}), 
            .integrator4({integrator4}), .integrator4_71__N_634({integrator4_71__N_634}), 
            .integrator5_71__N_706({integrator5_71__N_706}), .comb6({comb6}), 
            .comb6_71__N_1451({comb6_71__N_1451}), .cic_sine_clk(cic_sine_clk), 
            .comb_d6({comb_d6}), .comb7({comb7}), .comb7_71__N_1523({comb7_71__N_1523}), 
            .comb_d7({comb_d7}), .comb8({comb8}), .comb8_71__N_1595({comb8_71__N_1595}), 
            .comb_d8({comb_d8}), .comb9({comb9}), .comb9_71__N_1667({comb9_71__N_1667}), 
            .comb_d9({comb_d9}), .mult_i_b({mult_i_b}), .integrator1({integrator1}), 
            .integrator1_71__N_418({integrator1_71__N_418}), .count({count}), 
            .n32(n32_adj_2968), .n35(n35_adj_2965), .n34(n34_adj_2966), 
            .n37(n37_adj_2963), .n36(n36_adj_2964), .n67({n28_adj_5077, 
            n31_adj_5078, n34_adj_5079, n37_adj_5080, n40_adj_5081, 
            n43_adj_5082, n46_adj_5083, n49_adj_5084, n52_adj_5085, 
            n55_adj_5086, n58_adj_5087, n61_adj_5088}), .\cic_gain[0] (cic_gain[0]), 
            .\comb10[66] (comb10_adj_6033[66]), .\comb10[67] (comb10_adj_6033[67]), 
            .\comb10[69] (comb10_adj_6033[69]), .\comb10[68] (comb10_adj_6033[68]), 
            .\comb10[65] (comb10_adj_6033[65]), .\cic_gain[1] (cic_gain[1]), 
            .\comb10[70] (comb10_adj_6033[70]), .\comb10[71] (comb10_adj_6033[71]), 
            .n63(n63), .\data_out_11__N_1811[2] (data_out_11__N_1811_adj_6058[2]), 
            .n64(n64), .\data_out_11__N_1811[3] (data_out_11__N_1811_adj_6058[3]), 
            .n65(n65_adj_4746), .\data_out_11__N_1811[4] (data_out_11__N_1811_adj_6058[4]), 
            .n66(n66), .\data_out_11__N_1811[5] (data_out_11__N_1811_adj_6058[5]), 
            .\data_out_11__N_1811[6] (data_out_11__N_1811_adj_6058[6]), .\data_out_11__N_1811[7] (data_out_11__N_1811_adj_6058[7]), 
            .n118(n118_adj_5862), .n120(n120_adj_5903), .cout(cout_adj_5306), 
            .n115(n115_adj_5861), .n117(n117_adj_5902), .n112(n112_adj_5860), 
            .n114(n114_adj_5901), .n109(n109_adj_5859), .n111(n111_adj_5900), 
            .n106(n106_adj_5858), .n108(n108_adj_5899), .n103(n103_adj_5857), 
            .n105(n105_adj_5898), .n100(n100_adj_5856), .n102(n102_adj_5897), 
            .\comb10[64] (comb10_adj_6033[64]), .\comb10[62] (comb10_adj_6033[62]), 
            .\comb10[63] (comb10_adj_6033[63]), .n97(n97_adj_5855), .n99(n99_adj_5896), 
            .\comb10[61] (comb10_adj_6033[61]), .n94(n94_adj_5854), .n96(n96_adj_5895), 
            .n91(n91_adj_5853), .n93(n93_adj_5894), .n16607(n16607), .\comb10[59] (comb10_adj_6033[59]), 
            .n62(n62_adj_4745), .\comb10[60] (comb10_adj_6033[60]), .n88(n88_adj_5852), 
            .n90(n90_adj_5893), .n85(n85_adj_5851), .n87(n87_adj_5892), 
            .n82(n82_adj_5850), .n84(n84_adj_5891), .n79(n79_adj_5849), 
            .n81(n81_adj_5890), .n76(n76_adj_5848), .n78(n78_adj_5889), 
            .n3(n3_adj_4767), .n2(n2_adj_4766), .n5(n5_adj_4769), .n4(n4_adj_4768), 
            .n7(n7_adj_4771), .n6(n6_adj_4770), .n9(n9_adj_4773), .n8(n8_adj_4772), 
            .n11(n11_adj_4775), .n10(n10_adj_4774), .n13(n13_adj_4777), 
            .n12(n12_adj_4776), .n15(n15_adj_4779), .n14(n14_adj_4778), 
            .n17(n17_adj_4781), .n16(n16_adj_4780), .n19(n19_adj_4783), 
            .n18(n18_adj_4782), .n21(n21_adj_4785), .n20(n20_adj_4784), 
            .n23(n23_adj_4787), .n22(n22_adj_4786), .n25(n25_adj_4789), 
            .n24(n24_adj_4788), .n27(n27_adj_4791), .n26(n26_adj_4790), 
            .n29(n29_adj_4793), .n28_adj_115(n28_adj_4792), .n31_adj_116(n31_adj_4795), 
            .n30_adj_117(n30_adj_4794), .n33_adj_118(n33_adj_4797), .n32_adj_119(n32_adj_4796), 
            .n35_adj_120(n35_adj_4799), .n34_adj_121(n34_adj_4798), .n37_adj_122(n37_adj_4801), 
            .n36_adj_123(n36_adj_4800), .n3_adj_124(n3), .n2_adj_125(n2), 
            .n5_adj_126(n5), .n4_adj_127(n4), .n3_adj_128(n3_adj_4803), 
            .n2_adj_129(n2_adj_4802), .n5_adj_130(n5_adj_4805), .n4_adj_131(n4_adj_4804), 
            .n7_adj_132(n7_adj_4807), .n6_adj_133(n6_adj_4806), .n9_adj_134(n9_adj_4809), 
            .n8_adj_135(n8_adj_4808), .n11_adj_136(n11_adj_4811), .n10_adj_137(n10_adj_4810), 
            .n13_adj_138(n13_adj_4813), .n12_adj_139(n12_adj_4812), .n15_adj_140(n15_adj_4815), 
            .n14_adj_141(n14_adj_4814), .n17_adj_142(n17_adj_4817), .n16_adj_143(n16_adj_4816), 
            .n19_adj_144(n19_adj_4819), .n18_adj_145(n18_adj_4818), .n21_adj_146(n21_adj_4821), 
            .n20_adj_147(n20_adj_4820), .n7_adj_148(n7), .n6_adj_149(n6), 
            .n9_adj_150(n9), .n8_adj_151(n8), .n11_adj_152(n11), .n10_adj_153(n10), 
            .n13_adj_154(n13), .n12_adj_155(n12), .n15_adj_156(n15), .n14_adj_157(n14), 
            .n17_adj_158(n17), .n16_adj_159(n16_adj_2947), .n19_adj_160(n19), 
            .\data_out_11__N_1811[10] (data_out_11__N_1811_adj_6058[10]), 
            .n18_adj_161(n18), .n21_adj_162(n21), .n20_adj_163(n20), .n23_adj_164(n23), 
            .n22_adj_165(n22), .n23_adj_166(n23_adj_4823), .n22_adj_167(n22_adj_4822), 
            .n25_adj_168(n25_adj_4825), .n24_adj_169(n24_adj_4824), .n27_adj_170(n27_adj_4827), 
            .\data_out_11__N_1811[11] (data_out_11__N_1811_adj_6058[11]), 
            .n26_adj_171(n26_adj_4826), .n29_adj_172(n29_adj_4829), .n28_adj_173(n28_adj_4828), 
            .n31_adj_174(n31_adj_4831), .n30_adj_175(n30_adj_4830), .n25_adj_176(n25), 
            .n24_adj_177(n24), .n33_adj_178(n33_adj_4833), .n32_adj_179(n32_adj_4832), 
            .n35_adj_180(n35_adj_4835), .n34_adj_181(n34_adj_4834), .n37_adj_182(n37_adj_4837), 
            .n36_adj_183(n36_adj_4836), .n27_adj_184(n27_adj_2946), .n26_adj_185(n26), 
            .n29_adj_186(n29), .n28_adj_187(n28), .n31_adj_188(n31), .n30_adj_189(n30), 
            .n33_adj_190(n33), .n32_adj_191(n32), .n35_adj_192(n35), .n34_adj_193(n34), 
            .n37_adj_194(n37), .n36_adj_195(n36), .\data_out_11__N_1811[8] (data_out_11__N_1811_adj_6058[8]), 
            .n3_adj_196(n3_adj_2961), .n2_adj_197(n2_adj_2962), .n5_adj_198(n5_adj_2959), 
            .n4_adj_199(n4_adj_2960), .n7_adj_200(n7_adj_2957), .\data_out_11__N_1811[9] (data_out_11__N_1811_adj_6058[9]), 
            .n6_adj_201(n6_adj_2958), .n9_adj_202(n9_adj_2955), .n8_adj_203(n8_adj_2956), 
            .n11_adj_204(n11_adj_2953), .n10_adj_205(n10_adj_2954), .n13_adj_206(n13_adj_2951), 
            .n12_adj_207(n12_adj_2952), .n15_adj_208(n15_adj_2949), .n14_adj_209(n14_adj_2950), 
            .n17_adj_210(n17_adj_4763), .n16_adj_211(n16), .n19_adj_212(n19_adj_4748), 
            .n18_adj_213(n18_adj_4761), .n21_adj_214(n21_adj_4743), .n20_adj_215(n20_adj_4744), 
            .n23_adj_216(n23_adj_4727), .n22_adj_217(n22_adj_4728), .n25_adj_218(n25_adj_2974), 
            .n24_adj_219(n24_adj_4716), .n27_adj_220(n27), .n26_adj_221(n26_adj_2973), 
            .n29_adj_222(n29_adj_2971), .n28_adj_223(n28_adj_2972), .n31_adj_224(n31_adj_2969)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(155[7] 161[6])
    FD1S3AX rx_byte_i4_rep_372 (.D(rx_byte1[3]), .CK(clk_80mhz), .Q(n17289));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(234[12] 260[8])
    defparam rx_byte_i4_rep_372.GSR = "ENABLED";
    CCU2C _add_1_1181_add_4_8 (.A0(integrator3[41]), .B0(integrator2[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[42]), .B1(integrator2[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15551), .COUT(n15552), .S0(n168_adj_5341), 
          .S1(n165_adj_5340));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_49 (.A0(phase_inc_gen[51]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[52]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15669), .COUT(n15670), .S0(n160), .S1(n157));
    defparam _add_1_1241_add_4_49.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_49.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_49.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_49.INJECT1_1 = "NO";
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 i5756_4_lut (.A(n17335), .B(led_c_3), .C(n17278), .D(n17144), 
         .Z(clk_80mhz_enable_1444)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))) */ ;
    defparam i5756_4_lut.init = 16'ha0a2;
    CCU2C _add_1_1181_add_4_6 (.A0(integrator3[39]), .B0(integrator2[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[40]), .B1(integrator2[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15550), .COUT(n15551), .S0(n174_adj_5343), 
          .S1(n171_adj_5342));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_4 (.A0(integrator3[37]), .B0(integrator2[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator3[38]), .B1(integrator2[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15549), .COUT(n15550), .S0(n180_adj_5345), 
          .S1(n177_adj_5344));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_1181_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1181_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator3[36]), .B1(integrator2[36]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15549), .S1(n183_adj_5346));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(68[20:45])
    defparam _add_1_1181_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1181_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_1181_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1181_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_38 (.A0(comb_d8_adj_6030[71]), .B0(comb8_adj_6029[71]), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15548), .S0(n78_adj_5624));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_38.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_38.INIT1 = 16'h0000;
    defparam _add_1_1142_add_4_38.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_38.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_36 (.A0(comb_d8_adj_6030[69]), .B0(comb8_adj_6029[69]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[70]), .B1(comb8_adj_6029[70]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15547), .COUT(n15548), .S0(n84_adj_5626), 
          .S1(n81_adj_5625));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_36.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_36.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_34 (.A0(comb_d8_adj_6030[67]), .B0(comb8_adj_6029[67]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[68]), .B1(comb8_adj_6029[68]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15546), .COUT(n15547), .S0(n90_adj_5628), 
          .S1(n87_adj_5627));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_34.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_32 (.A0(comb_d8_adj_6030[65]), .B0(comb8_adj_6029[65]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[66]), .B1(comb8_adj_6029[66]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15545), .COUT(n15546), .S0(n96_adj_5630), 
          .S1(n93_adj_5629));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_30 (.A0(comb_d8_adj_6030[63]), .B0(comb8_adj_6029[63]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[64]), .B1(comb8_adj_6029[64]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15544), .COUT(n15545), .S0(n102_adj_5632), 
          .S1(n99_adj_5631));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_28 (.A0(comb_d8_adj_6030[61]), .B0(comb8_adj_6029[61]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[62]), .B1(comb8_adj_6029[62]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15543), .COUT(n15544), .S0(n108_adj_5634), 
          .S1(n105_adj_5633));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_32 (.A0(integrator1_adj_6020[30]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[31]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15334), .COUT(n15335), .S0(integrator1_71__N_418_adj_6036[30]), 
          .S1(integrator1_71__N_418_adj_6036[31]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_32.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_32.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_32.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_26 (.A0(comb_d8_adj_6030[59]), .B0(comb8_adj_6029[59]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[60]), .B1(comb8_adj_6029[60]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15542), .COUT(n15543), .S0(n114_adj_5636), 
          .S1(n111_adj_5635));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_24 (.A0(integrator1_adj_6020[22]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[23]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15330), .COUT(n15331), .S0(integrator1_71__N_418_adj_6036[22]), 
          .S1(integrator1_71__N_418_adj_6036[23]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_24.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_24 (.A0(comb_d8_adj_6030[57]), .B0(comb8_adj_6029[57]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[58]), .B1(comb8_adj_6029[58]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15541), .COUT(n15542), .S0(n120_adj_5638), 
          .S1(n117_adj_5637));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_22 (.A0(comb_d8_adj_6030[55]), .B0(comb8_adj_6029[55]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[56]), .B1(comb8_adj_6029[56]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15540), .COUT(n15541), .S0(n126_adj_5640), 
          .S1(n123_adj_5639));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_20 (.A0(comb_d8_adj_6030[53]), .B0(comb8_adj_6029[53]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[54]), .B1(comb8_adj_6029[54]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15539), .COUT(n15540), .S0(n132_adj_5642), 
          .S1(n129_adj_5641));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_20.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_8 (.A0(phase_inc_gen1[6]), .B0(phase_accum[6]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[7]), .B1(phase_accum[7]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15472), .COUT(n15473), .S0(n303), 
          .S1(n300));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_8.INIT0 = 16'h666a;
    defparam phase_accum_add_4_8.INIT1 = 16'h666a;
    defparam phase_accum_add_4_8.INJECT1_0 = "NO";
    defparam phase_accum_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_18 (.A0(comb_d8_adj_6030[51]), .B0(comb8_adj_6029[51]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[52]), .B1(comb8_adj_6029[52]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15538), .COUT(n15539), .S0(n138_adj_5644), 
          .S1(n135_adj_5643));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_16 (.A0(comb_d8_adj_6030[49]), .B0(comb8_adj_6029[49]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[50]), .B1(comb8_adj_6029[50]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15537), .COUT(n15538), .S0(n144_adj_5646), 
          .S1(n141_adj_5645));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_16.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_6 (.A0(phase_inc_gen1[4]), .B0(phase_accum[4]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[5]), .B1(phase_accum[5]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15471), .COUT(n15472), .S0(n309), 
          .S1(n306));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_6.INIT0 = 16'h666a;
    defparam phase_accum_add_4_6.INIT1 = 16'h666a;
    defparam phase_accum_add_4_6.INJECT1_0 = "NO";
    defparam phase_accum_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_14 (.A0(comb_d8_adj_6030[47]), .B0(comb8_adj_6029[47]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[48]), .B1(comb8_adj_6029[48]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15536), .COUT(n15537), .S0(n150_adj_5648), 
          .S1(n147_adj_5647));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_12 (.A0(comb_d8_adj_6030[45]), .B0(comb8_adj_6029[45]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[46]), .B1(comb8_adj_6029[46]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15535), .COUT(n15536), .S0(n156_adj_5650), 
          .S1(n153_adj_5649));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_8 (.A0(integrator_d_tmp[5]), .B0(integrator_tmp[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[6]), .B1(integrator_tmp[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15347), .COUT(n15348), .S0(comb6_71__N_1451[5]), 
          .S1(comb6_71__N_1451[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_10 (.A0(comb_d8_adj_6030[43]), .B0(comb8_adj_6029[43]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[44]), .B1(comb8_adj_6029[44]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15534), .COUT(n15535), .S0(n162_adj_5652), 
          .S1(n159_adj_5651));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_47 (.A0(phase_inc_gen[49]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[50]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15668), .COUT(n15669), .S0(n166), .S1(n163));
    defparam _add_1_1241_add_4_47.INIT0 = 16'haaa0;
    defparam _add_1_1241_add_4_47.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_47.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_47.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_8 (.A0(comb_d8_adj_6030[41]), .B0(comb8_adj_6029[41]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[42]), .B1(comb8_adj_6029[42]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15533), .COUT(n15534), .S0(n168_adj_5654), 
          .S1(n165_adj_5653));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_6 (.A0(comb_d8_adj_6030[39]), .B0(comb8_adj_6029[39]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[40]), .B1(comb8_adj_6029[40]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15532), .COUT(n15533), .S0(n174_adj_5656), 
          .S1(n171_adj_5655));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_10 (.A0(integrator_d_tmp[7]), .B0(integrator_tmp[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[8]), .B1(integrator_tmp[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15348), .COUT(n15349), .S0(comb6_71__N_1451[7]), 
          .S1(comb6_71__N_1451[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_4 (.A0(comb_d8_adj_6030[37]), .B0(comb8_adj_6029[37]), 
          .C0(GND_net), .D0(VCC_net), .A1(comb_d8_adj_6030[38]), .B1(comb8_adj_6029[38]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15531), .COUT(n15532), .S0(n180_adj_5658), 
          .S1(n177_adj_5657));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1142_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1190_add_4_4 (.A0(n17132), .B0(square_sum[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(n17132), .B1(amdemod_d_11__N_2098), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15338), .COUT(n15339), .S0(amdemod_d_11__N_1850[1]), 
          .S1(amdemod_d_11__N_1850[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1190_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1190_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_1190_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1190_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1142_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(comb_d8_adj_6030[36]), .B1(comb8_adj_6029[36]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15531), .S1(n183_adj_5659));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam _add_1_1142_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1142_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1142_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1142_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1190_add_4_6 (.A0(amdemod_d_11__N_2095), .B0(amdemod_d_11__N_1841[11]), 
          .C0(n17134), .D0(amdemod_d_11__N_1840[11]), .A1(n17134), .B1(amdemod_d_11__N_2092), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15339), .COUT(n15340), .S0(amdemod_d_11__N_1850[3]), 
          .S1(amdemod_d_11__N_1850[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1190_add_4_6.INIT0 = 16'h656a;
    defparam _add_1_1190_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_1190_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1190_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_45 (.A0(phase_inc_gen[47]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[48]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15667), .COUT(n15668), .S0(n172), .S1(n169));
    defparam _add_1_1241_add_4_45.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_45.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_45.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_45.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_37 (.A0(comb7[70]), .B0(cout_adj_4986), .C0(n81_adj_5270), 
          .D0(n3_adj_4767), .A1(comb7[71]), .B1(cout_adj_4986), .C1(n78_adj_5269), 
          .D1(n2_adj_4766), .CIN(n15529), .S0(comb8_71__N_1595[70]), .S1(comb8_71__N_1595[71]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_37.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_37.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_35 (.A0(comb7[68]), .B0(cout_adj_4986), .C0(n87_adj_5272), 
          .D0(n5_adj_4769), .A1(comb7[69]), .B1(cout_adj_4986), .C1(n84_adj_5271), 
          .D1(n4_adj_4768), .CIN(n15528), .COUT(n15529), .S0(comb8_71__N_1595[68]), 
          .S1(comb8_71__N_1595[69]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_35.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_35.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_43 (.A0(phase_inc_gen[45]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[46]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15666), .COUT(n15667), .S0(n178), .S1(n175));
    defparam _add_1_1241_add_4_43.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_43.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_43.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_43.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_6 (.A0(integrator_d_tmp[3]), .B0(integrator_tmp[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[4]), .B1(integrator_tmp[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15346), .COUT(n15347), .S0(comb6_71__N_1451[3]), 
          .S1(comb6_71__N_1451[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_33 (.A0(comb7[66]), .B0(cout_adj_4986), .C0(n93_adj_5274), 
          .D0(n7_adj_4771), .A1(comb7[67]), .B1(cout_adj_4986), .C1(n90_adj_5273), 
          .D1(n6_adj_4770), .CIN(n15527), .COUT(n15528), .S0(comb8_71__N_1595[66]), 
          .S1(comb8_71__N_1595[67]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_33.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_33.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_33.INJECT1_1 = "NO";
    CCU2C _add_1_1190_add_4_8 (.A0(n17137), .B0(amdemod_d_11__N_2089), .C0(GND_net), 
          .D0(VCC_net), .A1(square_sum[23]), .B1(square_sum[22]), .C1(amdemod_d_11__N_2086), 
          .D1(VCC_net), .CIN(n15340), .COUT(n15341), .S0(amdemod_d_11__N_1850[5]), 
          .S1(amdemod_d_11__N_1850[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1190_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_1190_add_4_8.INIT1 = 16'he1e1;
    defparam _add_1_1190_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_1190_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_31 (.A0(comb7[64]), .B0(cout_adj_4986), .C0(n99_adj_5276), 
          .D0(n9_adj_4773), .A1(comb7[65]), .B1(cout_adj_4986), .C1(n96_adj_5275), 
          .D1(n8_adj_4772), .CIN(n15526), .COUT(n15527), .S0(comb8_71__N_1595[64]), 
          .S1(comb8_71__N_1595[65]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_31.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_31.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_41 (.A0(phase_inc_gen[43]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[44]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15665), .COUT(n15666), .S0(n184), .S1(n181));
    defparam _add_1_1241_add_4_41.INIT0 = 16'haaa0;
    defparam _add_1_1241_add_4_41.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_41.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_41.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_29 (.A0(comb7[62]), .B0(cout_adj_4986), .C0(n105_adj_5278), 
          .D0(n11_adj_4775), .A1(comb7[63]), .B1(cout_adj_4986), .C1(n102_adj_5277), 
          .D1(n10_adj_4774), .CIN(n15525), .COUT(n15526), .S0(comb8_71__N_1595[62]), 
          .S1(comb8_71__N_1595[63]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_29.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_29.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_27 (.A0(comb7[60]), .B0(cout_adj_4986), .C0(n111_adj_5280), 
          .D0(n13_adj_4777), .A1(comb7[61]), .B1(cout_adj_4986), .C1(n108_adj_5279), 
          .D1(n12_adj_4776), .CIN(n15524), .COUT(n15525), .S0(comb8_71__N_1595[60]), 
          .S1(comb8_71__N_1595[61]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_27.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_27.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_34 (.A0(integrator1_adj_6020[32]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[33]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15335), .COUT(n15336), .S0(integrator1_71__N_418_adj_6036[32]), 
          .S1(integrator1_71__N_418_adj_6036[33]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_34.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_34.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_34.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_25 (.A0(comb7[58]), .B0(cout_adj_4986), .C0(n117_adj_5282), 
          .D0(n15_adj_4779), .A1(comb7[59]), .B1(cout_adj_4986), .C1(n114_adj_5281), 
          .D1(n14_adj_4778), .CIN(n15523), .COUT(n15524), .S0(comb8_71__N_1595[58]), 
          .S1(comb8_71__N_1595[59]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_25.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_25.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_36 (.A0(integrator1_adj_6020[34]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[35]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15336), .COUT(n15337), .S0(integrator1_71__N_418_adj_6036[34]), 
          .S1(integrator1_71__N_418_adj_6036[35]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_36.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_36.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_36.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_36.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_23 (.A0(comb7[56]), .B0(cout_adj_4986), .C0(n123_adj_5284), 
          .D0(n17_adj_4781), .A1(comb7[57]), .B1(cout_adj_4986), .C1(n120_adj_5283), 
          .D1(n16_adj_4780), .CIN(n15522), .COUT(n15523), .S0(comb8_71__N_1595[56]), 
          .S1(comb8_71__N_1595[57]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_23.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_23.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_21 (.A0(comb7[54]), .B0(cout_adj_4986), .C0(n129_adj_5286), 
          .D0(n19_adj_4783), .A1(comb7[55]), .B1(cout_adj_4986), .C1(n126_adj_5285), 
          .D1(n18_adj_4782), .CIN(n15521), .COUT(n15522), .S0(comb8_71__N_1595[54]), 
          .S1(comb8_71__N_1595[55]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_21.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_21.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15337), .S0(cout_adj_5076));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_993_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_993_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_26 (.A0(integrator1_adj_6020[24]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[25]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15331), .COUT(n15332), .S0(integrator1_71__N_418_adj_6036[24]), 
          .S1(integrator1_71__N_418_adj_6036[25]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_26.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_26.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_19 (.A0(comb7[52]), .B0(cout_adj_4986), .C0(n135_adj_5288), 
          .D0(n21_adj_4785), .A1(comb7[53]), .B1(cout_adj_4986), .C1(n132_adj_5287), 
          .D1(n20_adj_4784), .CIN(n15520), .COUT(n15521), .S0(comb8_71__N_1595[52]), 
          .S1(comb8_71__N_1595[53]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_19.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_19.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_28 (.A0(integrator1_adj_6020[26]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[27]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15332), .COUT(n15333), .S0(integrator1_71__N_418_adj_6036[26]), 
          .S1(integrator1_71__N_418_adj_6036[27]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_28.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_28.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_17 (.A0(comb7[50]), .B0(cout_adj_4986), .C0(n141_adj_5290), 
          .D0(n23_adj_4787), .A1(comb7[51]), .B1(cout_adj_4986), .C1(n138_adj_5289), 
          .D1(n22_adj_4786), .CIN(n15519), .COUT(n15520), .S0(comb8_71__N_1595[50]), 
          .S1(comb8_71__N_1595[51]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_17.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_17.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_39 (.A0(phase_inc_gen[41]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[42]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15664), .COUT(n15665), .S0(n190), .S1(n187));
    defparam _add_1_1241_add_4_39.INIT0 = 16'haaa0;
    defparam _add_1_1241_add_4_39.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_39.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_39.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_4 (.A0(phase_inc_gen1[2]), .B0(phase_accum[2]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[3]), .B1(phase_accum[3]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15470), .COUT(n15471), .S0(n315), 
          .S1(n312));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_4.INIT0 = 16'h666a;
    defparam phase_accum_add_4_4.INIT1 = 16'h666a;
    defparam phase_accum_add_4_4.INJECT1_0 = "NO";
    defparam phase_accum_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_15 (.A0(comb7[48]), .B0(cout_adj_4986), .C0(n147_adj_5292), 
          .D0(n25_adj_4789), .A1(comb7[49]), .B1(cout_adj_4986), .C1(n144_adj_5291), 
          .D1(n24_adj_4788), .CIN(n15518), .COUT(n15519), .S0(comb8_71__N_1595[48]), 
          .S1(comb8_71__N_1595[49]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_15.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_15.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_13 (.A0(comb7[46]), .B0(cout_adj_4986), .C0(n153_adj_5294), 
          .D0(n27_adj_4791), .A1(comb7[47]), .B1(cout_adj_4986), .C1(n150_adj_5293), 
          .D1(n26_adj_4790), .CIN(n15517), .COUT(n15518), .S0(comb8_71__N_1595[46]), 
          .S1(comb8_71__N_1595[47]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_13.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_13.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1250_add_4_9 (.A0(square_sum[23]), .B0(square_sum[22]), 
          .C0(amdemod_d_11__N_1850[5]), .D0(VCC_net), .A1(amdemod_d_11__N_1850[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n15465), .COUT(n15466), 
          .S0(n50), .S1(n47));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1250_add_4_9.INIT0 = 16'h1e1e;
    defparam _add_1_1250_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1250_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1250_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_37 (.A0(phase_inc_gen[39]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[40]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15663), .COUT(n15664), .S0(n196), .S1(n193));
    defparam _add_1_1241_add_4_37.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_37.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_37.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_37.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_30 (.A0(integrator1_adj_6020[28]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[29]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15333), .COUT(n15334), .S0(integrator1_71__N_418_adj_6036[28]), 
          .S1(integrator1_71__N_418_adj_6036[29]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_30.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_30.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_11 (.A0(comb7[44]), .B0(cout_adj_4986), .C0(n159_adj_5296), 
          .D0(n29_adj_4793), .A1(comb7[45]), .B1(cout_adj_4986), .C1(n156_adj_5295), 
          .D1(n28_adj_4792), .CIN(n15516), .COUT(n15517), .S0(comb8_71__N_1595[44]), 
          .S1(comb8_71__N_1595[45]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_11.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_11.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_9 (.A0(comb7[42]), .B0(cout_adj_4986), .C0(n165_adj_5298), 
          .D0(n31_adj_4795), .A1(comb7[43]), .B1(cout_adj_4986), .C1(n162_adj_5297), 
          .D1(n30_adj_4794), .CIN(n15515), .COUT(n15516), .S0(comb8_71__N_1595[42]), 
          .S1(comb8_71__N_1595[43]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_9.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_9.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_993_add_4_22 (.A0(integrator1_adj_6020[20]), .B0(mix_cosinewave[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator1_adj_6020[21]), .B1(mix_cosinewave[11]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15329), .COUT(n15330), .S0(integrator1_71__N_418_adj_6036[20]), 
          .S1(integrator1_71__N_418_adj_6036[21]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(66[20:45])
    defparam _add_1_993_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_993_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_993_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_993_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_7 (.A0(comb7[40]), .B0(cout_adj_4986), .C0(n171_adj_5300), 
          .D0(n33_adj_4797), .A1(comb7[41]), .B1(cout_adj_4986), .C1(n168_adj_5299), 
          .D1(n32_adj_4796), .CIN(n15514), .COUT(n15515), .S0(comb8_71__N_1595[40]), 
          .S1(comb8_71__N_1595[41]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_7.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_7.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_5 (.A0(comb7[38]), .B0(cout_adj_4986), .C0(n177_adj_5302), 
          .D0(n35_adj_4799), .A1(comb7[39]), .B1(cout_adj_4986), .C1(n174_adj_5301), 
          .D1(n34_adj_4798), .CIN(n15513), .COUT(n15514), .S0(comb8_71__N_1595[38]), 
          .S1(comb8_71__N_1595[39]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_5.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_5.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(integrator_d_tmp[0]), .B1(integrator_tmp[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15345), .S1(comb6_71__N_1451[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_1115_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_3 (.A0(comb7[36]), .B0(cout_adj_4986), .C0(n183_adj_5304), 
          .D0(n37_adj_4801), .A1(comb7[37]), .B1(cout_adj_4986), .C1(n180_adj_5303), 
          .D1(n36_adj_4800), .CIN(n15512), .COUT(n15513), .S0(comb8_71__N_1595[36]), 
          .S1(comb8_71__N_1595[37]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_1070_add_4_3.INIT1 = 16'hd1e2;
    defparam _add_1_1070_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1250_add_4_7 (.A0(n17134), .B0(amdemod_d_11__N_1850[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1850[4]), .B1(n17162), 
          .C1(n17279), .D1(n17146), .CIN(n15464), .COUT(n15465), .S0(n56), 
          .S1(n53));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1250_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1250_add_4_7.INIT1 = 16'h596a;
    defparam _add_1_1250_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1250_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1070_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cout_adj_4986), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15512));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam _add_1_1070_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1070_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_1070_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1070_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_15 (.A0(amdemod_d_11__N_2137), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15508), .S0(amdemod_d_11__N_1861[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1023_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1023_add_4_15.INIT1 = 16'h0000;
    defparam _add_1_1023_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1190_add_4_16 (.A0(amdemod_d_11__N_2065), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15344), .S0(amdemod_d_11__N_1850[13]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam _add_1_1190_add_4_16.INIT0 = 16'h555f;
    defparam _add_1_1190_add_4_16.INIT1 = 16'h0000;
    defparam _add_1_1190_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_1190_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_35 (.A0(phase_inc_gen[37]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[38]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15662), .COUT(n15663), .S0(n202), .S1(n199));
    defparam _add_1_1241_add_4_35.INIT0 = 16'haaa0;
    defparam _add_1_1241_add_4_35.INIT1 = 16'h555f;
    defparam _add_1_1241_add_4_35.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_35.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_13 (.A0(amdemod_d_11__N_2143), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2140), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15507), .COUT(n15508), .S0(amdemod_d_11__N_1861[11]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1023_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1023_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1023_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_11 (.A0(amdemod_d_11__N_2149), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_2146), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15506), .COUT(n15507), .S0(amdemod_d_11__N_1861[9]), 
          .S1(amdemod_d_11__N_1861[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1023_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1023_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1023_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1115_add_4_4 (.A0(integrator_d_tmp[1]), .B0(integrator_tmp[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator_d_tmp[2]), .B1(integrator_tmp[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15345), .COUT(n15346), .S0(comb6_71__N_1451[1]), 
          .S1(comb6_71__N_1451[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam _add_1_1115_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_1115_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_1115_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_1115_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_9 (.A0(amdemod_d_11__N_2155), .B0(n17162), .C0(n17279), 
          .D0(n17146), .A1(square_sum[23]), .B1(square_sum[22]), .C1(amdemod_d_11__N_2152), 
          .D1(VCC_net), .CIN(n15505), .COUT(n15506), .S0(amdemod_d_11__N_1861[7]), 
          .S1(amdemod_d_11__N_1861[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1023_add_4_9.INIT0 = 16'h596a;
    defparam _add_1_1023_add_4_9.INIT1 = 16'h1e1e;
    defparam _add_1_1023_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_9.INJECT1_1 = "NO";
    PFUMX i5820 (.BLUT(n17176), .ALUT(n17177), .C0(n16220), .Z(n17178));
    CCU2C _add_1_1023_add_4_7 (.A0(n17133), .B0(amdemod_d_11__N_2161), .C0(GND_net), 
          .D0(VCC_net), .A1(n17134), .B1(amdemod_d_11__N_2158), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15504), .COUT(n15505), .S0(amdemod_d_11__N_1861[5]), 
          .S1(amdemod_d_11__N_1861[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1023_add_4_7.INIT0 = 16'h9995;
    defparam _add_1_1023_add_4_7.INIT1 = 16'h9995;
    defparam _add_1_1023_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_5 (.A0(n17131), .B0(amdemod_d_11__N_2167), .C0(GND_net), 
          .D0(VCC_net), .A1(n17132), .B1(amdemod_d_11__N_2164), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15503), .COUT(n15504), .S0(amdemod_d_11__N_1861[3]), 
          .S1(amdemod_d_11__N_1861[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1023_add_4_5.INIT0 = 16'h9995;
    defparam _add_1_1023_add_4_5.INIT1 = 16'h9995;
    defparam _add_1_1023_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_33 (.A0(phase_inc_gen[35]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[36]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15661), .COUT(n15662), .S0(n208), .S1(n205));
    defparam _add_1_1241_add_4_33.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_33.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_33.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_2 (.A0(phase_inc_gen1[0]), .B0(phase_accum[0]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[1]), .B1(phase_accum[1]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n15470), .S1(n318));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_2.INIT0 = 16'h0008;
    defparam phase_accum_add_4_2.INIT1 = 16'h666a;
    defparam phase_accum_add_4_2.INJECT1_0 = "NO";
    defparam phase_accum_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_3 (.A0(n17130), .B0(square_sum[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(n17130), .B1(amdemod_d_11__N_2170), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15502), .COUT(n15503), .S0(amdemod_d_11__N_1861[1]), 
          .S1(amdemod_d_11__N_1861[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1023_add_4_3.INIT0 = 16'h666a;
    defparam _add_1_1023_add_4_3.INIT1 = 16'h9995;
    defparam _add_1_1023_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1023_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(square_sum[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n15502), .S1(amdemod_d_11__N_1861[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1023_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1023_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1023_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1023_add_4_1.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_64 (.A0(phase_inc_gen1[62]), .B0(phase_acc[62]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[63]), .B1(phase_acc[63]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15500), .S0(n135_adj_5661), 
          .S1(n132_adj_5660));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_64.INIT0 = 16'h666a;
    defparam phase_accum_add_4_64.INIT1 = 16'h666a;
    defparam phase_accum_add_4_64.INJECT1_0 = "NO";
    defparam phase_accum_add_4_64.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_62 (.A0(phase_inc_gen1[60]), .B0(phase_acc[60]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[61]), .B1(phase_acc[61]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15499), .COUT(n15500), .S0(n141_adj_5663), 
          .S1(n138_adj_5662));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_62.INIT0 = 16'h666a;
    defparam phase_accum_add_4_62.INIT1 = 16'h666a;
    defparam phase_accum_add_4_62.INJECT1_0 = "NO";
    defparam phase_accum_add_4_62.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_31 (.A0(phase_inc_gen[33]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[34]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15660), .COUT(n15661), .S0(n214), .S1(n211));
    defparam _add_1_1241_add_4_31.INIT0 = 16'haaa0;
    defparam _add_1_1241_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_31.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_60 (.A0(phase_inc_gen1[58]), .B0(phase_acc[58]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[59]), .B1(phase_acc[59]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15498), .COUT(n15499), .S0(n147_adj_5665), 
          .S1(n144_adj_5664));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_60.INIT0 = 16'h666a;
    defparam phase_accum_add_4_60.INIT1 = 16'h666a;
    defparam phase_accum_add_4_60.INJECT1_0 = "NO";
    defparam phase_accum_add_4_60.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_58 (.A0(phase_inc_gen1[56]), .B0(phase_acc[56]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[57]), .B1(phase_acc[57]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15497), .COUT(n15498), .S0(n153_adj_5667), 
          .S1(n150_adj_5666));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_58.INIT0 = 16'h666a;
    defparam phase_accum_add_4_58.INIT1 = 16'h666a;
    defparam phase_accum_add_4_58.INJECT1_0 = "NO";
    defparam phase_accum_add_4_58.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_56 (.A0(phase_inc_gen1[54]), .B0(phase_accum[54]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[55]), .B1(phase_accum[55]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15496), .COUT(n15497), .S0(n159_adj_5669), 
          .S1(n156_adj_5668));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_56.INIT0 = 16'h666a;
    defparam phase_accum_add_4_56.INIT1 = 16'h666a;
    defparam phase_accum_add_4_56.INJECT1_0 = "NO";
    defparam phase_accum_add_4_56.INJECT1_1 = "NO";
    CCU2C _add_1_1241_add_4_29 (.A0(phase_inc_gen[31]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(phase_inc_gen[32]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n15659), .COUT(n15660), .S0(n220), .S1(n217));
    defparam _add_1_1241_add_4_29.INIT0 = 16'h555f;
    defparam _add_1_1241_add_4_29.INIT1 = 16'haaa0;
    defparam _add_1_1241_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1241_add_4_29.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_54 (.A0(phase_inc_gen1[52]), .B0(phase_accum[52]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[53]), .B1(phase_accum[53]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15495), .COUT(n15496), .S0(n165_adj_5671), 
          .S1(n162_adj_5670));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_54.INIT0 = 16'h666a;
    defparam phase_accum_add_4_54.INIT1 = 16'h666a;
    defparam phase_accum_add_4_54.INJECT1_0 = "NO";
    defparam phase_accum_add_4_54.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_52 (.A0(phase_inc_gen1[50]), .B0(phase_accum[50]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[51]), .B1(phase_accum[51]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15494), .COUT(n15495), .S0(n171_adj_5673), 
          .S1(n168_adj_5672));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_52.INIT0 = 16'h666a;
    defparam phase_accum_add_4_52.INIT1 = 16'h666a;
    defparam phase_accum_add_4_52.INJECT1_0 = "NO";
    defparam phase_accum_add_4_52.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_50 (.A0(phase_inc_gen1[48]), .B0(phase_accum[48]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[49]), .B1(phase_accum[49]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15493), .COUT(n15494), .S0(n177_adj_5675), 
          .S1(n174_adj_5674));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_50.INIT0 = 16'h666a;
    defparam phase_accum_add_4_50.INIT1 = 16'h666a;
    defparam phase_accum_add_4_50.INJECT1_0 = "NO";
    defparam phase_accum_add_4_50.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_48 (.A0(phase_inc_gen1[46]), .B0(phase_accum[46]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[47]), .B1(phase_accum[47]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15492), .COUT(n15493), .S0(n183_adj_5677), 
          .S1(n180_adj_5676));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_48.INIT0 = 16'h666a;
    defparam phase_accum_add_4_48.INIT1 = 16'h666a;
    defparam phase_accum_add_4_48.INJECT1_0 = "NO";
    defparam phase_accum_add_4_48.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_46 (.A0(phase_inc_gen1[44]), .B0(phase_accum[44]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[45]), .B1(phase_accum[45]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15491), .COUT(n15492), .S0(n189), 
          .S1(n186));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_46.INIT0 = 16'h666a;
    defparam phase_accum_add_4_46.INIT1 = 16'h666a;
    defparam phase_accum_add_4_46.INJECT1_0 = "NO";
    defparam phase_accum_add_4_46.INJECT1_1 = "NO";
    CCU2C _add_1_981_add_4_10 (.A0(integrator2[8]), .B0(integrator1[8]), 
          .C0(GND_net), .D0(VCC_net), .A1(integrator2[9]), .B1(integrator1[9]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15429), .COUT(n15430), .S0(integrator2_71__N_490[8]), 
          .S1(integrator2_71__N_490[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(67[20:45])
    defparam _add_1_981_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_981_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_981_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_981_add_4_10.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_44 (.A0(phase_inc_gen1[42]), .B0(phase_accum[42]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[43]), .B1(phase_accum[43]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15490), .COUT(n15491), .S0(n195), 
          .S1(n192));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_44.INIT0 = 16'h666a;
    defparam phase_accum_add_4_44.INIT1 = 16'h666a;
    defparam phase_accum_add_4_44.INJECT1_0 = "NO";
    defparam phase_accum_add_4_44.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_42 (.A0(phase_inc_gen1[40]), .B0(phase_accum[40]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[41]), .B1(phase_accum[41]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15489), .COUT(n15490), .S0(n201), 
          .S1(n198));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_42.INIT0 = 16'h666a;
    defparam phase_accum_add_4_42.INIT1 = 16'h666a;
    defparam phase_accum_add_4_42.INJECT1_0 = "NO";
    defparam phase_accum_add_4_42.INJECT1_1 = "NO";
    CCU2C _add_1_1250_add_4_15 (.A0(amdemod_d_11__N_1850[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15468), .S0(n32_adj_4715));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1250_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1250_add_4_15.INIT1 = 16'h0000;
    defparam _add_1_1250_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1250_add_4_15.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_40 (.A0(phase_inc_gen1[38]), .B0(phase_accum[38]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[39]), .B1(phase_accum[39]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15488), .COUT(n15489), .S0(n207), 
          .S1(n204));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_40.INIT0 = 16'h666a;
    defparam phase_accum_add_4_40.INIT1 = 16'h666a;
    defparam phase_accum_add_4_40.INJECT1_0 = "NO";
    defparam phase_accum_add_4_40.INJECT1_1 = "NO";
    CCU2C _add_1_1250_add_4_13 (.A0(amdemod_d_11__N_1850[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(amdemod_d_11__N_1850[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15467), .COUT(n15468), .S0(n38));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam _add_1_1250_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1250_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1250_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1250_add_4_13.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_38 (.A0(phase_inc_gen1[36]), .B0(phase_accum[36]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[37]), .B1(phase_accum[37]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15487), .COUT(n15488), .S0(n213), 
          .S1(n210));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_38.INIT0 = 16'h666a;
    defparam phase_accum_add_4_38.INIT1 = 16'h666a;
    defparam phase_accum_add_4_38.INJECT1_0 = "NO";
    defparam phase_accum_add_4_38.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_36 (.A0(phase_inc_gen1[34]), .B0(phase_accum[34]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[35]), .B1(phase_accum[35]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15486), .COUT(n15487), .S0(n219), 
          .S1(n216));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_36.INIT0 = 16'h666a;
    defparam phase_accum_add_4_36.INIT1 = 16'h666a;
    defparam phase_accum_add_4_36.INJECT1_0 = "NO";
    defparam phase_accum_add_4_36.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_34 (.A0(phase_inc_gen1[32]), .B0(phase_accum[32]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[33]), .B1(phase_accum[33]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15485), .COUT(n15486), .S0(n225), 
          .S1(n222));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_34.INIT0 = 16'h666a;
    defparam phase_accum_add_4_34.INIT1 = 16'h666a;
    defparam phase_accum_add_4_34.INJECT1_0 = "NO";
    defparam phase_accum_add_4_34.INJECT1_1 = "NO";
    PWM pwm_inst (.\data_in_reg[0] (data_in_reg[0]), .clk_80mhz(clk_80mhz), 
        .\data_in_reg_11__N_2339[0] (data_in_reg_11__N_2339[0]), .count({count_adj_6105}), 
        .\data_in_reg[1] (data_in_reg[1]), .\data_in_reg_11__N_2339[1] (data_in_reg_11__N_2339[1]), 
        .\data_in_reg[2] (data_in_reg[2]), .\data_in_reg_11__N_2339[2] (data_in_reg_11__N_2339[2]), 
        .\data_in_reg[3] (data_in_reg[3]), .\data_in_reg_11__N_2339[3] (data_in_reg_11__N_2339[3]), 
        .\data_in_reg[4] (data_in_reg[4]), .\data_in_reg_11__N_2339[4] (data_in_reg_11__N_2339[4]), 
        .\data_in_reg[5] (data_in_reg[5]), .\data_in_reg_11__N_2339[5] (data_in_reg_11__N_2339[5]), 
        .\data_in_reg[6] (data_in_reg[6]), .\data_in_reg_11__N_2339[6] (data_in_reg_11__N_2339[6]), 
        .\data_in_reg[7] (data_in_reg[7]), .\data_in_reg_11__N_2339[7] (data_in_reg_11__N_2339[7]), 
        .\data_in_reg[8] (data_in_reg[8]), .\data_in_reg_11__N_2339[8] (data_in_reg_11__N_2339[8]), 
        .\data_in_reg[9] (data_in_reg[9]), .GND_net(GND_net), .VCC_net(VCC_net), 
        .\amdemod_out[9] (amdemod_out[9])) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(198[7] 202[6])
    PFUMX i5818 (.BLUT(n17172), .ALUT(n17173), .C0(n316), .Z(n17174));
    SinCos SinCos_inst (.clk_80mhz(clk_80mhz), .VCC_net(VCC_net), .GND_net(GND_net), 
           .\phase_acc[57] (phase_acc[57]), .\phase_acc[58] (phase_acc[58]), 
           .\phase_acc[59] (phase_acc[59]), .\phase_acc[60] (phase_acc[60]), 
           .\phase_acc[61] (phase_acc[61]), .\phase_acc[62] (phase_acc[62]), 
           .\phase_acc[63] (phase_acc[63]), .\lo_sinewave[1] (lo_sinewave[1]), 
           .\lo_sinewave[2] (lo_sinewave[2]), .\lo_sinewave[3] (lo_sinewave[3]), 
           .\lo_sinewave[4] (lo_sinewave[4]), .\lo_sinewave[5] (lo_sinewave[5]), 
           .\lo_sinewave[6] (lo_sinewave[6]), .\lo_sinewave[7] (lo_sinewave[7]), 
           .\lo_sinewave[8] (lo_sinewave[8]), .\lo_sinewave[9] (lo_sinewave[9]), 
           .\lo_sinewave[10] (lo_sinewave[10]), .\lo_sinewave[11] (lo_sinewave[11]), 
           .\lo_sinewave[12] (lo_sinewave[12]), .\lo_cosinewave[1] (lo_cosinewave[1]), 
           .\lo_cosinewave[2] (lo_cosinewave[2]), .\lo_cosinewave[3] (lo_cosinewave[3]), 
           .\lo_cosinewave[4] (lo_cosinewave[4]), .\lo_cosinewave[5] (lo_cosinewave[5]), 
           .\lo_cosinewave[6] (lo_cosinewave[6]), .\lo_cosinewave[7] (lo_cosinewave[7]), 
           .\lo_cosinewave[8] (lo_cosinewave[8]), .\lo_cosinewave[9] (lo_cosinewave[9]), 
           .\lo_cosinewave[10] (lo_cosinewave[10]), .\lo_cosinewave[11] (lo_cosinewave[11]), 
           .\lo_cosinewave[12] (lo_cosinewave[12]), .\phase_acc[56] (phase_acc[56])) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    CCU2C phase_accum_add_4_32 (.A0(phase_inc_gen1[30]), .B0(phase_accum[30]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[31]), .B1(phase_accum[31]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15484), .COUT(n15485), .S0(n231), 
          .S1(n228));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_32.INIT0 = 16'h666a;
    defparam phase_accum_add_4_32.INIT1 = 16'h666a;
    defparam phase_accum_add_4_32.INJECT1_0 = "NO";
    defparam phase_accum_add_4_32.INJECT1_1 = "NO";
    CCU2C phase_accum_add_4_30 (.A0(phase_inc_gen1[28]), .B0(phase_accum[28]), 
          .C0(GND_net), .D0(VCC_net), .A1(phase_inc_gen1[29]), .B1(phase_accum[29]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n15483), .COUT(n15484), .S0(n237), 
          .S1(n234));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/NCO.v(39[20:48])
    defparam phase_accum_add_4_30.INIT0 = 16'h666a;
    defparam phase_accum_add_4_30.INIT1 = 16'h666a;
    defparam phase_accum_add_4_30.INJECT1_0 = "NO";
    defparam phase_accum_add_4_30.INJECT1_1 = "NO";
    \CIC(REGISTER_WIDTH=72,DECIMATION_RATIO=4096)_U0  cic_cosine_inst (.comb_d6({comb_d6_adj_6026}), 
            .n21(n21_adj_4893), .n20(n20_adj_4892), .integrator_tmp({integrator_tmp_adj_6018}), 
            .clk_80mhz(clk_80mhz), .integrator5({integrator5_adj_6024}), 
            .integrator_d_tmp({integrator_d_tmp_adj_6019}), .integrator2({integrator2_adj_6021}), 
            .integrator2_71__N_490({integrator2_71__N_490_adj_6037}), .integrator3({integrator3_adj_6022}), 
            .integrator3_71__N_562({integrator3_71__N_562_adj_6038}), .integrator4({integrator4_adj_6023}), 
            .integrator4_71__N_634({integrator4_71__N_634_adj_6039}), .integrator5_71__N_706({integrator5_71__N_706_adj_6040}), 
            .comb6({comb6_adj_6025}), .comb6_71__N_1451({comb6_71__N_1451_adj_6052}), 
            .comb7({comb7_adj_6027}), .comb7_71__N_1523({comb7_71__N_1523_adj_6053}), 
            .comb_d7({comb_d7_adj_6028}), .comb8({comb8_adj_6029}), .comb8_71__N_1595({comb8_71__N_1595_adj_6054}), 
            .comb_d8({comb_d8_adj_6030}), .comb9({comb9_adj_6031}), .comb9_71__N_1667({comb9_71__N_1667_adj_6055}), 
            .comb_d9({comb_d9_adj_6032}), .n23(n23_adj_4895), .cic_cosine_out({cic_cosine_out}), 
            .integrator1({integrator1_adj_6020}), .integrator1_71__N_418({integrator1_71__N_418_adj_6036}), 
            .n22(n22_adj_4894), .n25(n25_adj_4897), .n3(n3_adj_4839), 
            .n2(n2_adj_4838), .n5(n5_adj_4841), .n24(n24_adj_4896), .n4(n4_adj_4840), 
            .n27(n27_adj_4899), .n26(n26_adj_4898), .n7(n7_adj_4843), 
            .n6(n6_adj_4842), .n9(n9_adj_4845), .n29(n29_adj_4901), .n8(n8_adj_4844), 
            .n28(n28_adj_4900), .n31(n31_adj_4903), .n30(n30_adj_4902), 
            .n11(n11_adj_4847), .count({count_adj_6035}), .n67({n28_adj_5167, 
            n31_adj_5168, n34_adj_5169, n37_adj_5170, n40_adj_5171, 
            n43_adj_5172, n46_adj_5173, n49_adj_5174, n52_adj_5175, 
            n55_adj_5176, n58_adj_5177, n61_adj_5178}), .n33(n33_adj_4905), 
            .n10(n10_adj_4846), .n13(n13_adj_4849), .n12(n12_adj_4848), 
            .n15(n15_adj_4851), .n32(n32_adj_4904), .n14(n14_adj_4850), 
            .n17(n17_adj_4853), .n16(n16_adj_4852), .n19(n19_adj_4855), 
            .n18(n18_adj_4854), .n35(n35_adj_4907), .n21_adj_3(n21_adj_4857), 
            .n20_adj_4(n20_adj_4856), .n23_adj_5(n23_adj_4859), .n34_adj_6(n34_adj_4906), 
            .n37_adj_7(n37_adj_4909), .n22_adj_8(n22_adj_4858), .n36(n36_adj_4908), 
            .n25_adj_9(n25_adj_4861), .n3_adj_10(n3_adj_4911), .n24_adj_11(n24_adj_4860), 
            .n27_adj_12(n27_adj_4863), .\cic_gain[1] (cic_gain[1]), .\comb10[59] (comb10_adj_6033[59]), 
            .n16607(n16607), .n2_adj_13(n2_adj_4910), .n5_adj_14(n5_adj_4913), 
            .n3_adj_15(n3_adj_4947), .\comb10[60] (comb10_adj_6033[60]), 
            .n62(n62_adj_4745), .n2_adj_16(n2_adj_4946), .n5_adj_17(n5_adj_4949), 
            .n26_adj_18(n26_adj_4862), .n29_adj_19(n29_adj_4865), .n4_adj_20(n4_adj_4912), 
            .n28_adj_21(n28_adj_4864), .n4_adj_22(n4_adj_4948), .n7_adj_23(n7_adj_4915), 
            .n7_adj_24(n7_adj_4951), .n6_adj_25(n6_adj_4950), .n9_adj_26(n9_adj_4953), 
            .n8_adj_27(n8_adj_4952), .n6_adj_28(n6_adj_4914), .n9_adj_29(n9_adj_4917), 
            .n8_adj_30(n8_adj_4916), .n11_adj_31(n11_adj_4919), .n10_adj_32(n10_adj_4918), 
            .n13_adj_33(n13_adj_4921), .n12_adj_34(n12_adj_4920), .n15_adj_35(n15_adj_4923), 
            .n14_adj_36(n14_adj_4922), .n17_adj_37(n17_adj_4925), .n16_adj_38(n16_adj_4924), 
            .n19_adj_39(n19_adj_4927), .n18_adj_40(n18_adj_4926), .n31_adj_41(n31_adj_4867), 
            .n21_adj_42(n21_adj_4929), .n20_adj_43(n20_adj_4928), .n23_adj_44(n23_adj_4931), 
            .n22_adj_45(n22_adj_4930), .n30_adj_46(n30_adj_4866), .n33_adj_47(n33_adj_4869), 
            .n32_adj_48(n32_adj_4868), .n35_adj_49(n35_adj_4871), .n34_adj_50(n34_adj_4870), 
            .n37_adj_51(n37_adj_4873), .n36_adj_52(n36_adj_4872), .n25_adj_53(n25_adj_4933), 
            .n3_adj_54(n3_adj_4875), .n24_adj_55(n24_adj_4932), .n27_adj_56(n27_adj_4935), 
            .n2_adj_57(n2_adj_4874), .n26_adj_58(n26_adj_4934), .n29_adj_59(n29_adj_4937), 
            .n5_adj_60(n5_adj_4877), .n28_adj_61(n28_adj_4936), .n4_adj_62(n4_adj_4876), 
            .n7_adj_63(n7_adj_4879), .n6_adj_64(n6_adj_4878), .n9_adj_65(n9_adj_4881), 
            .n8_adj_66(n8_adj_4880), .n11_adj_67(n11_adj_4883), .n10_adj_68(n10_adj_4882), 
            .n13_adj_69(n13_adj_4885), .n12_adj_70(n12_adj_4884), .n15_adj_71(n15_adj_4887), 
            .n14_adj_72(n14_adj_4886), .n17_adj_73(n17_adj_4889), .n16_adj_74(n16_adj_4888), 
            .n19_adj_75(n19_adj_4891), .n18_adj_76(n18_adj_4890), .n31_adj_77(n31_adj_4939), 
            .n11_adj_78(n11_adj_4955), .n10_adj_79(n10_adj_4954), .n13_adj_80(n13_adj_4957), 
            .n12_adj_81(n12_adj_4956), .n15_adj_82(n15_adj_4959), .n14_adj_83(n14_adj_4958), 
            .n30_adj_84(n30_adj_4938), .\comb10[61] (comb10_adj_6033[61]), 
            .\comb10[62] (comb10_adj_6033[62]), .\comb10[63] (comb10_adj_6033[63]), 
            .\comb10[64] (comb10_adj_6033[64]), .\comb10[65] (comb10_adj_6033[65]), 
            .\comb10[66] (comb10_adj_6033[66]), .\comb10[67] (comb10_adj_6033[67]), 
            .\comb10[68] (comb10_adj_6033[68]), .\comb10[69] (comb10_adj_6033[69]), 
            .\comb10[70] (comb10_adj_6033[70]), .\comb10[71] (comb10_adj_6033[71]), 
            .\data_out_11__N_1811[2] (data_out_11__N_1811_adj_6058[2]), .\data_out_11__N_1811[3] (data_out_11__N_1811_adj_6058[3]), 
            .\data_out_11__N_1811[4] (data_out_11__N_1811_adj_6058[4]), .\data_out_11__N_1811[5] (data_out_11__N_1811_adj_6058[5]), 
            .\data_out_11__N_1811[6] (data_out_11__N_1811_adj_6058[6]), .\data_out_11__N_1811[7] (data_out_11__N_1811_adj_6058[7]), 
            .\data_out_11__N_1811[8] (data_out_11__N_1811_adj_6058[8]), .\data_out_11__N_1811[9] (data_out_11__N_1811_adj_6058[9]), 
            .\data_out_11__N_1811[10] (data_out_11__N_1811_adj_6058[10]), 
            .\data_out_11__N_1811[11] (data_out_11__N_1811_adj_6058[11]), 
            .n33_adj_85(n33_adj_4941), .n32_adj_86(n32_adj_4940), .n35_adj_87(n35_adj_4943), 
            .n34_adj_88(n34_adj_4942), .n37_adj_89(n37_adj_4945), .n36_adj_90(n36_adj_4944), 
            .n118(n118), .n120(n120_adj_5597), .cout(cout_adj_5125), .n115(n115), 
            .n117(n117_adj_5596), .n112(n112), .n114(n114_adj_5595), .n109(n109), 
            .n111(n111_adj_5594), .n106(n106), .n108(n108_adj_5593), .n103(n103), 
            .n105(n105_adj_5592), .n100(n100), .n102(n102_adj_5591), .n97(n97), 
            .n99(n99_adj_5590), .n94(n94), .n96(n96_adj_5589), .n91(n91), 
            .n93(n93_adj_5588), .n88(n88), .n90(n90_adj_5587), .n85(n85), 
            .n87(n87_adj_5586), .n82(n82), .n84(n84_adj_5585), .n79(n79_adj_5497), 
            .n81(n81_adj_5584), .n76(n76_adj_5496), .n78(n78_adj_5583), 
            .\cic_gain[0] (cic_gain[0]), .n63(n63), .n64(n64), .n65(n65_adj_4746), 
            .n66(n66), .n17_adj_91(n17_adj_4961), .n16_adj_92(n16_adj_4960), 
            .n19_adj_93(n19_adj_4963), .n18_adj_94(n18_adj_4962), .n21_adj_95(n21_adj_4965), 
            .n20_adj_96(n20_adj_4964), .n23_adj_97(n23_adj_4967), .n22_adj_98(n22_adj_4966), 
            .n25_adj_99(n25_adj_4969), .n24_adj_100(n24_adj_4968), .n27_adj_101(n27_adj_4971), 
            .n26_adj_102(n26_adj_4970), .n29_adj_103(n29_adj_4973), .n28_adj_104(n28_adj_4972), 
            .n31_adj_105(n31_adj_4975), .n30_adj_106(n30_adj_4974), .n33_adj_107(n33_adj_4977), 
            .n32_adj_108(n32_adj_4976), .n35_adj_109(n35_adj_4979), .n34_adj_110(n34_adj_4978), 
            .n37_adj_111(n37_adj_4981), .n36_adj_112(n36_adj_4980)) /* synthesis syn_module_defined=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(171[7] 177[6])
    
endmodule
//
// Verilog Description of module \uart_rx(CLKS_PER_BIT=87) 
//

module \uart_rx(CLKS_PER_BIT=87)  (clk_80mhz, rx_serial_c, rx_byte1, rx_data_valid1, 
            GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input clk_80mhz;
    input rx_serial_c;
    output [7:0]rx_byte1;
    output rx_data_valid1;
    input GND_net;
    input VCC_net;
    
    wire [7:0]UartClk /* synthesis SET_AS_NETWORK=\uart_rx_inst/UartClk[2], is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(37[14:21])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(64[10:19])
    wire [15:0]r_Clock_Count;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(39[18:31])
    
    wire UartClk_2_enable_36, n11936;
    wire [15:0]n69;
    wire [2:0]r_SM_Main;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(43[17:26])
    
    wire n17033, r_Rx_DV_last, r_Rx_DV, r_Rx_Data_R, r_Rx_Data, UartClk_2_enable_27;
    wire [7:0]r_Rx_Byte;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(41[17:26])
    wire [2:0]r_Bit_Index;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(40[17:28])
    
    wire UartClk_2_enable_8, n16350;
    wire [2:0]n30;
    wire [2:0]n17;
    
    wire n16352, n16329, UartClk_2_enable_9, UartClk_2_enable_10, UartClk_2_enable_11, 
        UartClk_2_enable_12, UartClk_2_enable_13, n17161, n15925, n17032, 
        n17138, UartClk_2_enable_14, n12346, n16212, n17151, n12318, 
        n17031, n17156, n17140, r_Rx_DV_N_2466, UartClk_2_enable_15, 
        UartClk_2_enable_29, n16234, UartClk_2_enable_33, n24, n16463, 
        n12320, n16437, n16315, n16433, n17166, n11933, r_Rx_DV_last_N_2465, 
        n14844, n14843, n14842, n14841, n14840, n14839, n14838, 
        n14837, n14514, n17145, n16455;
    wire [2:0]n132;
    
    wire n26, n17165, n17164, n16459;
    
    FD1P3IX r_Clock_Count_505__i4 (.D(n69[4]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i4.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i0 (.D(n17033), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i0.GSR = "ENABLED";
    FD1S3AX r_Rx_DV_last_60 (.D(r_Rx_DV), .CK(clk_80mhz), .Q(r_Rx_DV_last)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(47[11] 52[8])
    defparam r_Rx_DV_last_60.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_R_61 (.D(rx_serial_c), .CK(UartClk[2]), .Q(r_Rx_Data_R)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(57[11] 62[8])
    defparam r_Rx_Data_R_61.GSR = "ENABLED";
    FD1S3AY r_Rx_Data_62 (.D(r_Rx_Data_R), .CK(UartClk[2]), .Q(r_Rx_Data)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(57[11] 62[8])
    defparam r_Rx_Data_62.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i3 (.D(n69[3]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i3.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i2 (.D(n69[2]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i2.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i0 (.D(r_Rx_Byte[0]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(rx_byte1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i0.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i0 (.D(n16350), .SP(UartClk_2_enable_8), .CK(UartClk[2]), 
            .Q(r_Bit_Index[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i0.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i1 (.D(n69[1]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i1.GSR = "ENABLED";
    FD1S3AX UartClk_503_541__i0 (.D(n17[0]), .CK(clk_80mhz), .Q(n30[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_503_541__i0.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i2 (.D(n16352), .SP(UartClk_2_enable_8), .CK(UartClk[2]), 
            .Q(r_Bit_Index[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i2.GSR = "ENABLED";
    FD1P3AX r_Bit_Index_i1 (.D(n16329), .SP(UartClk_2_enable_8), .CK(UartClk[2]), 
            .Q(r_Bit_Index[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Bit_Index_i1.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i7 (.D(r_Rx_Data), .SP(UartClk_2_enable_9), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i7.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i6 (.D(r_Rx_Data), .SP(UartClk_2_enable_10), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i5 (.D(r_Rx_Data), .SP(UartClk_2_enable_11), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i4 (.D(r_Rx_Data), .SP(UartClk_2_enable_12), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i3 (.D(r_Rx_Data), .SP(UartClk_2_enable_13), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i3.GSR = "ENABLED";
    LUT4 r_SM_Main_2__N_2400_2__bdd_3_lut_4_lut (.A(n17161), .B(n15925), 
         .C(r_SM_Main[0]), .D(r_Rx_Data), .Z(n17032)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D))) */ ;
    defparam r_SM_Main_2__N_2400_2__bdd_3_lut_4_lut.init = 16'hd0df;
    LUT4 i5737_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n17138), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_14)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(114[17:39])
    defparam i5737_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_354 (.A(n12346), .B(n16212), .Z(n17151)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_354.init = 16'heeee;
    LUT4 r_SM_Main_2__N_2400_2__bdd_3_lut_5773_4_lut (.A(n12346), .B(n16212), 
         .C(r_SM_Main[0]), .D(n12318), .Z(n17031)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam r_SM_Main_2__N_2400_2__bdd_3_lut_5773_4_lut.init = 16'h1e10;
    LUT4 i1_2_lut_rep_341_3_lut_4_lut (.A(n12346), .B(n16212), .C(r_SM_Main[0]), 
         .D(n17156), .Z(n17138)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;
    defparam i1_2_lut_rep_341_3_lut_4_lut.init = 16'hfff1;
    LUT4 i5719_2_lut_3_lut_4_lut (.A(n12346), .B(n16212), .C(r_SM_Main[0]), 
         .D(n17156), .Z(UartClk_2_enable_27)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i5719_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i5739_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n17138), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_13)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(114[17:39])
    defparam i5739_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1724_2_lut_rep_343_3_lut (.A(n12346), .B(n16212), .C(r_SM_Main[0]), 
         .Z(n17140)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;
    defparam i1724_2_lut_rep_343_3_lut.init = 16'hf1f1;
    LUT4 i5759_2_lut_3_lut_4_lut (.A(n12346), .B(n16212), .C(n17156), 
         .D(r_SM_Main[0]), .Z(r_Rx_DV_N_2466)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i5759_2_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 i5734_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n17138), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_15)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(114[17:39])
    defparam i5734_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i5715_2_lut_3_lut_4_lut (.A(r_Bit_Index[2]), .B(n17138), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_29)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(114[17:39])
    defparam i5715_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_rep_359 (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .Z(n17156)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_359.init = 16'hbbbb;
    LUT4 i5747_2_lut_4_lut (.A(r_Bit_Index[2]), .B(n17138), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_10)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(114[17:39])
    defparam i5747_2_lut_4_lut.init = 16'h0200;
    LUT4 i5732_2_lut_3_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .Z(n16234)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(69[7] 161[14])
    defparam i5732_2_lut_3_lut.init = 16'hdfdf;
    LUT4 i21_4_lut_4_lut (.A(r_SM_Main[1]), .B(r_SM_Main[2]), .C(r_SM_Main[0]), 
         .D(n17151), .Z(UartClk_2_enable_33)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(69[7] 161[14])
    defparam i21_4_lut_4_lut.init = 16'h2505;
    LUT4 i5742_2_lut_4_lut (.A(r_Bit_Index[2]), .B(n17138), .C(r_Bit_Index[0]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_12)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(114[17:39])
    defparam i5742_2_lut_4_lut.init = 16'h0002;
    LUT4 i5762_3_lut_4_lut (.A(n17151), .B(r_SM_Main[0]), .C(r_Bit_Index[0]), 
         .D(r_SM_Main[1]), .Z(n16350)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(69[7] 161[14])
    defparam i5762_3_lut_4_lut.init = 16'h0200;
    FD1P3AX r_Rx_Byte_i2 (.D(r_Rx_Data), .SP(UartClk_2_enable_14), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX r_Rx_Byte_i1 (.D(r_Rx_Data), .SP(UartClk_2_enable_15), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i1.GSR = "ENABLED";
    LUT4 i5745_2_lut_4_lut (.A(r_Bit_Index[0]), .B(n17138), .C(r_Bit_Index[2]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_11)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i5745_2_lut_4_lut.init = 16'h0020;
    LUT4 i1_4_lut (.A(r_SM_Main[2]), .B(n24), .C(n17151), .D(r_SM_Main[1]), 
         .Z(n11936)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i1_4_lut.init = 16'h5044;
    LUT4 i1_4_lut_adj_189 (.A(r_Rx_Data), .B(r_SM_Main[0]), .C(n15925), 
         .D(n17161), .Z(n24)) /* synthesis lut_function=(!(A (B)+!A (B (C+!(D))))) */ ;
    defparam i1_4_lut_adj_189.init = 16'h3733;
    LUT4 i1_4_lut_adj_190 (.A(r_Clock_Count[1]), .B(n16212), .C(n16463), 
         .D(r_Clock_Count[6]), .Z(n15925)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(85[17:52])
    defparam i1_4_lut_adj_190.init = 16'hfffd;
    LUT4 i5749_2_lut_4_lut (.A(r_Bit_Index[0]), .B(n17138), .C(r_Bit_Index[2]), 
         .D(r_Bit_Index[1]), .Z(UartClk_2_enable_9)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i5749_2_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut (.A(r_Clock_Count[2]), .B(r_Clock_Count[4]), .Z(n16463)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(85[17:52])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2604_4_lut (.A(n12320), .B(r_Clock_Count[6]), .C(r_Clock_Count[5]), 
         .D(r_Clock_Count[4]), .Z(n12346)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i2604_4_lut.init = 16'hc8c0;
    LUT4 i2580_3_lut (.A(r_Clock_Count[1]), .B(r_Clock_Count[3]), .C(r_Clock_Count[2]), 
         .Z(n12320)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2580_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_191 (.A(n16437), .B(n16315), .C(n16433), .D(r_Clock_Count[11]), 
         .Z(n16212)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(85[17:52])
    defparam i1_4_lut_adj_191.init = 16'hfffe;
    FD1S3IX r_SM_Main_i2 (.D(n17151), .CK(UartClk[2]), .CD(n16234), .Q(r_SM_Main[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_192 (.A(r_Clock_Count[12]), .B(r_Clock_Count[10]), 
         .Z(n16437)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_192.init = 16'heeee;
    LUT4 i1_4_lut_adj_193 (.A(r_Clock_Count[9]), .B(r_Clock_Count[7]), .C(r_Clock_Count[14]), 
         .D(r_Clock_Count[15]), .Z(n16315)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(85[17:52])
    defparam i1_4_lut_adj_193.init = 16'hfffe;
    LUT4 i1_2_lut_adj_194 (.A(r_Clock_Count[8]), .B(r_Clock_Count[13]), 
         .Z(n16433)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(85[17:52])
    defparam i1_2_lut_adj_194.init = 16'heeee;
    FD1P3IX r_Clock_Count_505__i15 (.D(n69[15]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[15])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i15.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i14 (.D(n69[14]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[14])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i14.GSR = "ENABLED";
    FD1S3IX r_SM_Main_i1 (.D(n17166), .CK(UartClk[2]), .CD(r_SM_Main[2]), 
            .Q(r_SM_Main[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_SM_Main_i1.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i1 (.D(r_Rx_Byte[1]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(rx_byte1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i1.GSR = "ENABLED";
    FD1S3IX o_Rx_DV_59 (.D(r_Rx_DV_last_N_2465), .CK(clk_80mhz), .CD(n11933), 
            .Q(rx_data_valid1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(47[11] 52[8])
    defparam o_Rx_DV_59.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i13 (.D(n69[13]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[13])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i13.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i12 (.D(n69[12]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[12])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i12.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i11 (.D(n69[11]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[11])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i11.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i2 (.D(r_Rx_Byte[2]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(rx_byte1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i2.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i3 (.D(r_Rx_Byte[3]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(rx_byte1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i3.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i4 (.D(r_Rx_Byte[4]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(rx_byte1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i4.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i5 (.D(r_Rx_Byte[5]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(rx_byte1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i5.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i6 (.D(r_Rx_Byte[6]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(rx_byte1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i6.GSR = "ENABLED";
    FD1P3AX o_Rx_Byte_i7 (.D(r_Rx_Byte[7]), .SP(UartClk_2_enable_27), .CK(UartClk[2]), 
            .Q(rx_byte1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam o_Rx_Byte_i7.GSR = "ENABLED";
    FD1S3AX UartClk_503_541__i1 (.D(n17[1]), .CK(clk_80mhz), .Q(n30[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_503_541__i1.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i10 (.D(n69[10]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[10])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i10.GSR = "ENABLED";
    FD1S3AX UartClk_503_541__i2 (.D(n17[2]), .CK(clk_80mhz), .Q(UartClk[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_503_541__i2.GSR = "ENABLED";
    CCU2C r_Clock_Count_505_add_4_17 (.A0(r_Clock_Count[15]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n14844), .S0(n69[15]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505_add_4_17.INIT0 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_17.INIT1 = 16'h0000;
    defparam r_Clock_Count_505_add_4_17.INJECT1_0 = "NO";
    defparam r_Clock_Count_505_add_4_17.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_505_add_4_15 (.A0(r_Clock_Count[13]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[14]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14843), .COUT(n14844), .S0(n69[13]), 
          .S1(n69[14]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505_add_4_15.INIT0 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_15.INIT1 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_15.INJECT1_0 = "NO";
    defparam r_Clock_Count_505_add_4_15.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_505_add_4_13 (.A0(r_Clock_Count[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14842), .COUT(n14843), .S0(n69[11]), 
          .S1(n69[12]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505_add_4_13.INIT0 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_13.INIT1 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_13.INJECT1_0 = "NO";
    defparam r_Clock_Count_505_add_4_13.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_505_add_4_11 (.A0(r_Clock_Count[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14841), .COUT(n14842), .S0(n69[9]), 
          .S1(n69[10]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505_add_4_11.INIT0 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_11.INIT1 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_11.INJECT1_0 = "NO";
    defparam r_Clock_Count_505_add_4_11.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_505_add_4_9 (.A0(r_Clock_Count[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14840), .COUT(n14841), .S0(n69[7]), 
          .S1(n69[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505_add_4_9.INIT0 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_9.INIT1 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_9.INJECT1_0 = "NO";
    defparam r_Clock_Count_505_add_4_9.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_505_add_4_7 (.A0(r_Clock_Count[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14839), .COUT(n14840), .S0(n69[5]), 
          .S1(n69[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505_add_4_7.INIT0 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_7.INIT1 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_7.INJECT1_0 = "NO";
    defparam r_Clock_Count_505_add_4_7.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_505_add_4_5 (.A0(r_Clock_Count[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14838), .COUT(n14839), .S0(n69[3]), 
          .S1(n69[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505_add_4_5.INIT0 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_5.INIT1 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_5.INJECT1_0 = "NO";
    defparam r_Clock_Count_505_add_4_5.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_505_add_4_3 (.A0(r_Clock_Count[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(r_Clock_Count[2]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n14837), .COUT(n14838), .S0(n69[1]), 
          .S1(n69[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505_add_4_3.INIT0 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_3.INIT1 = 16'haaa0;
    defparam r_Clock_Count_505_add_4_3.INJECT1_0 = "NO";
    defparam r_Clock_Count_505_add_4_3.INJECT1_1 = "NO";
    CCU2C r_Clock_Count_505_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(r_Clock_Count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n14837), .S1(n69[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505_add_4_1.INIT0 = 16'h0000;
    defparam r_Clock_Count_505_add_4_1.INIT1 = 16'h555f;
    defparam r_Clock_Count_505_add_4_1.INJECT1_0 = "NO";
    defparam r_Clock_Count_505_add_4_1.INJECT1_1 = "NO";
    FD1P3AX r_Rx_Byte_i0 (.D(r_Rx_Data), .SP(UartClk_2_enable_29), .CK(UartClk[2]), 
            .Q(r_Rx_Byte[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_Byte_i0.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i9 (.D(n69[9]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i9.GSR = "ENABLED";
    CCU2C UartClk_503_541_add_4_3 (.A0(n30[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(UartClk[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n14514), .S0(n17[1]), .S1(n17[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_503_541_add_4_3.INIT0 = 16'haaa0;
    defparam UartClk_503_541_add_4_3.INIT1 = 16'haaa0;
    defparam UartClk_503_541_add_4_3.INJECT1_0 = "NO";
    defparam UartClk_503_541_add_4_3.INJECT1_1 = "NO";
    CCU2C UartClk_503_541_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n14514), .S1(n17[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(49[15:29])
    defparam UartClk_503_541_add_4_1.INIT0 = 16'h0000;
    defparam UartClk_503_541_add_4_1.INIT1 = 16'h555f;
    defparam UartClk_503_541_add_4_1.INJECT1_0 = "NO";
    defparam UartClk_503_541_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_348_4_lut (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), 
         .C(r_Clock_Count[0]), .D(n15925), .Z(n17145)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_348_4_lut.init = 16'hff7f;
    LUT4 i5710_4_lut (.A(n16455), .B(n16212), .C(n12346), .D(r_SM_Main[1]), 
         .Z(UartClk_2_enable_8)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;
    defparam i5710_4_lut.init = 16'h5455;
    LUT4 i1_2_lut_adj_195 (.A(r_SM_Main[0]), .B(r_SM_Main[2]), .Z(n16455)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_195.init = 16'heeee;
    LUT4 i1_4_lut_adj_196 (.A(n132[2]), .B(n17140), .C(n12318), .D(r_SM_Main[1]), 
         .Z(n16352)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_196.init = 16'h0200;
    LUT4 i745_3_lut (.A(r_Bit_Index[2]), .B(r_Bit_Index[1]), .C(r_Bit_Index[0]), 
         .Z(n132[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(119[36:54])
    defparam i745_3_lut.init = 16'h6a6a;
    LUT4 i1_3_lut (.A(r_Bit_Index[1]), .B(r_Bit_Index[0]), .C(r_Bit_Index[2]), 
         .Z(n12318)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i39_2_lut (.A(r_Bit_Index[0]), .B(r_Bit_Index[1]), .Z(n26)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i39_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_197 (.A(n26), .B(n17151), .C(r_SM_Main[0]), .D(r_SM_Main[1]), 
         .Z(n16329)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_197.init = 16'h0800;
    LUT4 i5444_3_lut_rep_364 (.A(r_Clock_Count[3]), .B(r_Clock_Count[5]), 
         .C(r_Clock_Count[0]), .Z(n17161)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5444_3_lut_rep_364.init = 16'h8080;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut (.A(r_SM_Main[0]), 
         .B(n16212), .C(n12346), .Z(n17165)) /* synthesis lut_function=(!(A (B+(C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(69[7] 161[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_then_3_lut.init = 16'h5757;
    LUT4 r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut (.A(r_SM_Main[0]), 
         .B(n17145), .C(r_Rx_Data), .Z(n17164)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(69[7] 161[14])
    defparam r_SM_Main_2__I_0_69_Mux_1_i3_4_lut_else_3_lut.init = 16'h0202;
    LUT4 i5722_4_lut (.A(r_SM_Main[2]), .B(r_SM_Main[1]), .C(n17145), 
         .D(n16459), .Z(UartClk_2_enable_36)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(69[7] 161[14])
    defparam i5722_4_lut.init = 16'h5455;
    LUT4 i1_2_lut_adj_198 (.A(r_Rx_Data), .B(r_SM_Main[0]), .Z(n16459)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_198.init = 16'h8888;
    LUT4 i2193_1_lut (.A(r_Rx_DV), .Z(n11933)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam i2193_1_lut.init = 16'h5555;
    LUT4 r_Rx_DV_last_I_0_1_lut (.A(r_Rx_DV_last), .Z(r_Rx_DV_last_N_2465)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(50[30:43])
    defparam r_Rx_DV_last_I_0_1_lut.init = 16'h5555;
    PFUMX i5774 (.BLUT(n17032), .ALUT(n17031), .C0(r_SM_Main[1]), .Z(n17033));
    FD1P3IX r_Clock_Count_505__i8 (.D(n69[8]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i8.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i7 (.D(n69[7]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i7.GSR = "ENABLED";
    FD1P3AX r_Rx_DV_64 (.D(r_Rx_DV_N_2466), .SP(UartClk_2_enable_33), .CK(UartClk[2]), 
            .Q(r_Rx_DV)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=209, LSE_RLINE=214 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(66[10] 162[8])
    defparam r_Rx_DV_64.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i0 (.D(n69[0]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i0.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i6 (.D(n69[6]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i6.GSR = "ENABLED";
    FD1P3IX r_Clock_Count_505__i5 (.D(n69[5]), .SP(UartClk_2_enable_36), 
            .CD(n11936), .CK(UartClk[2]), .Q(r_Clock_Count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/UartRX.v(137[34:54])
    defparam r_Clock_Count_505__i5.GSR = "ENABLED";
    PFUMX i5813 (.BLUT(n17164), .ALUT(n17165), .C0(r_SM_Main[1]), .Z(n17166));
    
endmodule
//
// Verilog Description of module AMDemodulator
//

module AMDemodulator (cic_sine_clk, cic_cosine_out, \data_in_reg_11__N_2339[0] , 
            \square_sum[22] , \square_sum[23] , n11179, amdemod_d_11__N_1874, 
            amdemod_d_11__N_2023, amdemod_d_11__N_2146, amdemod_d_11__N_2149, 
            amdemod_d_11__N_2020, amdemod_d_11__N_2281, amdemod_d_11__N_2284, 
            amdemod_d_11__N_2026, amdemod_d_11__N_2152, \square_sum[21] , 
            \square_sum[20] , n4, \amdemod_d_11__N_1870[13] , \amdemod_d_11__N_1871[13] , 
            n17128, n80, n79, n78, n77, n76, n75, n74, n73, 
            n72, n71, n70, n69, n68, n67, n66, n65, n64, n63, 
            n62, n61, n60, n59, n58, n57, VCC_net, GND_net, 
            n17146, n17157, n34, n34_adj_225, n17134, n32, n32_adj_226, 
            n71_adj_227, n71_adj_228, n73_adj_229, n73_adj_230, n68_adj_231, 
            n68_adj_232, n70_adj_233, n70_adj_234, n65_adj_235, n65_adj_236, 
            n67_adj_237, n67_adj_238, n62_adj_239, n62_adj_240, n64_adj_241, 
            n64_adj_242, n59_adj_243, n59_adj_244, n61_adj_245, n61_adj_246, 
            n53, n53_adj_247, n55, n55_adj_248, n46, n46_adj_249, 
            n17132, n56, n56_adj_250, n58_adj_251, n58_adj_252, n41, 
            n41_adj_253, n50, n50_adj_254, n52, n52_adj_255, mult_i_b, 
            mult_result_i, n43, n43_adj_256, n47, n47_adj_257, n49, 
            n49_adj_258, n38, n38_adj_259, n40, n40_adj_260, n44, 
            n44_adj_261, n46_adj_262, n46_adj_263, n71_adj_264, n71_adj_265, 
            n17130, n41_adj_266, n41_adj_267, n43_adj_268, n43_adj_269, 
            n73_adj_270, n73_adj_271, n68_adj_272, n68_adj_273, n70_adj_274, 
            n70_adj_275, n65_adj_276, n65_adj_277, n67_adj_278, n67_adj_279, 
            n62_adj_280, n62_adj_281, \amdemod_d_11__N_1850[13] , \amdemod_d_11__N_1851[13] , 
            n17131, n17129, n64_adj_282, n64_adj_283, n59_adj_284, 
            n59_adj_285, n38_adj_286, n38_adj_287, n61_adj_288, n61_adj_289, 
            n40_adj_290, n40_adj_291, \amdemod_d_11__N_1880[13] , \amdemod_d_11__N_1881[13] , 
            n56_adj_292, n56_adj_293, n71_adj_294, n71_adj_295, n73_adj_296, 
            n73_adj_297, n58_adj_298, n58_adj_299, n53_adj_300, n53_adj_301, 
            n55_adj_302, n55_adj_303, n50_adj_304, n50_adj_305, n34_adj_306, 
            n34_adj_307, amdemod_d_11__N_2155, \data_in_reg_11__N_2339[1] , 
            \data_in_reg_11__N_2339[2] , \data_in_reg_11__N_2339[3] , \data_in_reg_11__N_2339[4] , 
            \data_in_reg_11__N_2339[5] , \data_in_reg_11__N_2339[6] , \data_in_reg_11__N_2339[7] , 
            \data_in_reg_11__N_2339[8] , \amdemod_out[9] , \amdemod_d_11__N_1860[13] , 
            \amdemod_d_11__N_1861[13] , n17127, amdemod_d_11__N_2287, 
            \amdemod_d_11__N_1840[11] , \amdemod_d_11__N_1841[11] , n52_adj_308, 
            n52_adj_309, n17163, n17137, n47_adj_310, n47_adj_311, 
            n49_adj_312, n49_adj_313, n44_adj_314, n44_adj_315, n46_adj_316, 
            n46_adj_317, n41_adj_318, n41_adj_319, n43_adj_320, n43_adj_321, 
            n38_adj_322, n38_adj_323, n40_adj_324, n40_adj_325, n17133, 
            n71_adj_326, n71_adj_327, n73_adj_328, n73_adj_329, n65_adj_330, 
            n65_adj_331, n67_adj_332, n67_adj_333, n68_adj_334, n68_adj_335, 
            n70_adj_336, n70_adj_337, n65_adj_338, n65_adj_339, n67_adj_340, 
            n67_adj_341, n62_adj_342, n62_adj_343, n64_adj_344, n64_adj_345, 
            n59_adj_346, n59_adj_347, n61_adj_348, n61_adj_349, amdemod_d_11__N_2290, 
            amdemod_d_11__N_2293, amdemod_d_11__N_2158, amdemod_d_11__N_2296, 
            amdemod_d_11__N_2161, n56_adj_350, n56_adj_351, amdemod_d_11__N_2167, 
            amdemod_d_11__N_2299, n34_adj_352, n34_adj_353, n68_adj_354, 
            n68_adj_355, n17162, amdemod_d_11__N_2302, amdemod_d_11__N_2164, 
            n58_adj_356, n58_adj_357, n39, n39_adj_358, n52_adj_441, 
            n52_adj_442, n44_adj_372, n44_adj_373, n46_adj_374, n46_adj_375, 
            n32_adj_376, n32_adj_377, amdemod_d_11__N_2305, n70_adj_378, 
            n70_adj_379, \amdemod_d_11__N_1830[1] , n34_adj_380, n34_adj_381, 
            n32_adj_382, n32_adj_383, n48, n48_adj_384, n53_adj_385, 
            n53_adj_386, amdemod_d_11__N_2308, amdemod_d_11__N_2311, n41_adj_387, 
            n41_adj_388, n36, n36_adj_389, n42, n42_adj_390, amdemod_d_11__N_2314, 
            amdemod_d_11__N_2209, amdemod_d_11__N_2170, n24, n24_adj_391, 
            amdemod_d_11__N_2212, n45, n45_adj_392, n30, n30_adj_393, 
            n33, n33_adj_394, amdemod_d_11__N_2215, n27, n27_adj_395, 
            amdemod_d_11__N_2218, amdemod_d_11__N_2221, amdemod_d_11__N_2224, 
            n56_adj_396, n56_adj_397, amdemod_d_11__N_2227, amdemod_d_11__N_2230, 
            n6, amdemod_d_11__N_2065, amdemod_d_11__N_2233, n58_adj_398, 
            n58_adj_399, amdemod_d_11__N_2236, amdemod_d_11__N_2068, amdemod_d_11__N_2239, 
            n17279, amdemod_d_11__N_2242, n53_adj_400, n53_adj_401, 
            n4_adj_402, amdemod_d_11__N_2071, amdemod_d_11__N_2137, amdemod_d_11__N_2074, 
            n62_adj_403, n62_adj_404, n64_adj_405, n64_adj_406, amdemod_d_11__N_2140, 
            amdemod_d_11__N_2077, n43_adj_407, n43_adj_408, n55_adj_409, 
            n55_adj_410, n50_adj_411, n50_adj_412, amdemod_d_11__N_2143, 
            amdemod_d_11__N_2083, amdemod_d_11__N_2080, n55_adj_413, n55_adj_414, 
            amdemod_d_11__N_2086, n38_adj_415, n38_adj_416, n59_adj_417, 
            n59_adj_418, amdemod_d_11__N_2089, n40_adj_419, n40_adj_420, 
            amdemod_d_11__N_2092, n61_adj_421, n61_adj_422, amdemod_d_11__N_2095, 
            amdemod_d_11__N_2098, amdemod_d_11__N_2005, n50_adj_423, n50_adj_424, 
            n52_adj_425, n52_adj_426, n52_adj_427, n52_adj_428, n32_adj_429, 
            n32_adj_430, amdemod_d_11__N_2011, n47_adj_431, n47_adj_432, 
            n47_adj_433, n47_adj_434, n49_adj_435, n49_adj_436, n49_adj_437, 
            n49_adj_438, n44_adj_439, n44_adj_440, amdemod_d_11__N_2008, 
            amdemod_d_11__N_2017, amdemod_d_11__N_2014) /* synthesis syn_module_defined=1 */ ;
    input cic_sine_clk;
    input [11:0]cic_cosine_out;
    output \data_in_reg_11__N_2339[0] ;
    input \square_sum[22] ;
    input \square_sum[23] ;
    output n11179;
    output amdemod_d_11__N_1874;
    output amdemod_d_11__N_2023;
    output amdemod_d_11__N_2146;
    output amdemod_d_11__N_2149;
    output amdemod_d_11__N_2020;
    output amdemod_d_11__N_2281;
    output amdemod_d_11__N_2284;
    output amdemod_d_11__N_2026;
    output amdemod_d_11__N_2152;
    input \square_sum[21] ;
    input \square_sum[20] ;
    output n4;
    input \amdemod_d_11__N_1870[13] ;
    input \amdemod_d_11__N_1871[13] ;
    output n17128;
    output n80;
    output n79;
    output n78;
    output n77;
    output n76;
    output n75;
    output n74;
    output n73;
    output n72;
    output n71;
    output n70;
    output n69;
    output n68;
    output n67;
    output n66;
    output n65;
    output n64;
    output n63;
    output n62;
    output n61;
    output n60;
    output n59;
    output n58;
    output n57;
    input VCC_net;
    input GND_net;
    output n17146;
    output n17157;
    input n34;
    input n34_adj_225;
    output n17134;
    input n32;
    input n32_adj_226;
    input n71_adj_227;
    input n71_adj_228;
    input n73_adj_229;
    input n73_adj_230;
    input n68_adj_231;
    input n68_adj_232;
    input n70_adj_233;
    input n70_adj_234;
    input n65_adj_235;
    input n65_adj_236;
    input n67_adj_237;
    input n67_adj_238;
    input n62_adj_239;
    input n62_adj_240;
    input n64_adj_241;
    input n64_adj_242;
    input n59_adj_243;
    input n59_adj_244;
    input n61_adj_245;
    input n61_adj_246;
    input n53;
    input n53_adj_247;
    input n55;
    input n55_adj_248;
    input n46;
    input n46_adj_249;
    output n17132;
    input n56;
    input n56_adj_250;
    input n58_adj_251;
    input n58_adj_252;
    input n41;
    input n41_adj_253;
    input n50;
    input n50_adj_254;
    input n52;
    input n52_adj_255;
    input [11:0]mult_i_b;
    output [23:0]mult_result_i;
    input n43;
    input n43_adj_256;
    input n47;
    input n47_adj_257;
    input n49;
    input n49_adj_258;
    input n38;
    input n38_adj_259;
    input n40;
    input n40_adj_260;
    input n44;
    input n44_adj_261;
    input n46_adj_262;
    input n46_adj_263;
    input n71_adj_264;
    input n71_adj_265;
    output n17130;
    input n41_adj_266;
    input n41_adj_267;
    input n43_adj_268;
    input n43_adj_269;
    input n73_adj_270;
    input n73_adj_271;
    input n68_adj_272;
    input n68_adj_273;
    input n70_adj_274;
    input n70_adj_275;
    input n65_adj_276;
    input n65_adj_277;
    input n67_adj_278;
    input n67_adj_279;
    input n62_adj_280;
    input n62_adj_281;
    input \amdemod_d_11__N_1850[13] ;
    input \amdemod_d_11__N_1851[13] ;
    output n17131;
    output n17129;
    input n64_adj_282;
    input n64_adj_283;
    input n59_adj_284;
    input n59_adj_285;
    input n38_adj_286;
    input n38_adj_287;
    input n61_adj_288;
    input n61_adj_289;
    input n40_adj_290;
    input n40_adj_291;
    input \amdemod_d_11__N_1880[13] ;
    input \amdemod_d_11__N_1881[13] ;
    input n56_adj_292;
    input n56_adj_293;
    input n71_adj_294;
    input n71_adj_295;
    input n73_adj_296;
    input n73_adj_297;
    input n58_adj_298;
    input n58_adj_299;
    input n53_adj_300;
    input n53_adj_301;
    input n55_adj_302;
    input n55_adj_303;
    input n50_adj_304;
    input n50_adj_305;
    input n34_adj_306;
    input n34_adj_307;
    output amdemod_d_11__N_2155;
    output \data_in_reg_11__N_2339[1] ;
    output \data_in_reg_11__N_2339[2] ;
    output \data_in_reg_11__N_2339[3] ;
    output \data_in_reg_11__N_2339[4] ;
    output \data_in_reg_11__N_2339[5] ;
    output \data_in_reg_11__N_2339[6] ;
    output \data_in_reg_11__N_2339[7] ;
    output \data_in_reg_11__N_2339[8] ;
    output \amdemod_out[9] ;
    input \amdemod_d_11__N_1860[13] ;
    input \amdemod_d_11__N_1861[13] ;
    output n17127;
    output amdemod_d_11__N_2287;
    input \amdemod_d_11__N_1840[11] ;
    input \amdemod_d_11__N_1841[11] ;
    input n52_adj_308;
    input n52_adj_309;
    output n17163;
    output n17137;
    input n47_adj_310;
    input n47_adj_311;
    input n49_adj_312;
    input n49_adj_313;
    input n44_adj_314;
    input n44_adj_315;
    input n46_adj_316;
    input n46_adj_317;
    input n41_adj_318;
    input n41_adj_319;
    input n43_adj_320;
    input n43_adj_321;
    input n38_adj_322;
    input n38_adj_323;
    input n40_adj_324;
    input n40_adj_325;
    output n17133;
    input n71_adj_326;
    input n71_adj_327;
    input n73_adj_328;
    input n73_adj_329;
    input n65_adj_330;
    input n65_adj_331;
    input n67_adj_332;
    input n67_adj_333;
    input n68_adj_334;
    input n68_adj_335;
    input n70_adj_336;
    input n70_adj_337;
    input n65_adj_338;
    input n65_adj_339;
    input n67_adj_340;
    input n67_adj_341;
    input n62_adj_342;
    input n62_adj_343;
    input n64_adj_344;
    input n64_adj_345;
    input n59_adj_346;
    input n59_adj_347;
    input n61_adj_348;
    input n61_adj_349;
    output amdemod_d_11__N_2290;
    output amdemod_d_11__N_2293;
    output amdemod_d_11__N_2158;
    output amdemod_d_11__N_2296;
    output amdemod_d_11__N_2161;
    input n56_adj_350;
    input n56_adj_351;
    output amdemod_d_11__N_2167;
    output amdemod_d_11__N_2299;
    input n34_adj_352;
    input n34_adj_353;
    input n68_adj_354;
    input n68_adj_355;
    output n17162;
    output amdemod_d_11__N_2302;
    output amdemod_d_11__N_2164;
    input n58_adj_356;
    input n58_adj_357;
    input n39;
    input n39_adj_358;
    input [8:0]n52_adj_441;
    input [8:0]n52_adj_442;
    input n44_adj_372;
    input n44_adj_373;
    input n46_adj_374;
    input n46_adj_375;
    input n32_adj_376;
    input n32_adj_377;
    output amdemod_d_11__N_2305;
    input n70_adj_378;
    input n70_adj_379;
    output \amdemod_d_11__N_1830[1] ;
    input n34_adj_380;
    input n34_adj_381;
    input n32_adj_382;
    input n32_adj_383;
    input n48;
    input n48_adj_384;
    input n53_adj_385;
    input n53_adj_386;
    output amdemod_d_11__N_2308;
    output amdemod_d_11__N_2311;
    input n41_adj_387;
    input n41_adj_388;
    input n36;
    input n36_adj_389;
    input n42;
    input n42_adj_390;
    output amdemod_d_11__N_2314;
    output amdemod_d_11__N_2209;
    output amdemod_d_11__N_2170;
    input n24;
    input n24_adj_391;
    output amdemod_d_11__N_2212;
    input n45;
    input n45_adj_392;
    input n30;
    input n30_adj_393;
    input n33;
    input n33_adj_394;
    output amdemod_d_11__N_2215;
    input n27;
    input n27_adj_395;
    output amdemod_d_11__N_2218;
    output amdemod_d_11__N_2221;
    output amdemod_d_11__N_2224;
    input n56_adj_396;
    input n56_adj_397;
    output amdemod_d_11__N_2227;
    output amdemod_d_11__N_2230;
    output n6;
    output amdemod_d_11__N_2065;
    output amdemod_d_11__N_2233;
    input n58_adj_398;
    input n58_adj_399;
    output amdemod_d_11__N_2236;
    output amdemod_d_11__N_2068;
    output amdemod_d_11__N_2239;
    output n17279;
    output amdemod_d_11__N_2242;
    input n53_adj_400;
    input n53_adj_401;
    output n4_adj_402;
    output amdemod_d_11__N_2071;
    output amdemod_d_11__N_2137;
    output amdemod_d_11__N_2074;
    input n62_adj_403;
    input n62_adj_404;
    input n64_adj_405;
    input n64_adj_406;
    output amdemod_d_11__N_2140;
    output amdemod_d_11__N_2077;
    input n43_adj_407;
    input n43_adj_408;
    input n55_adj_409;
    input n55_adj_410;
    input n50_adj_411;
    input n50_adj_412;
    output amdemod_d_11__N_2143;
    output amdemod_d_11__N_2083;
    output amdemod_d_11__N_2080;
    input n55_adj_413;
    input n55_adj_414;
    output amdemod_d_11__N_2086;
    input n38_adj_415;
    input n38_adj_416;
    input n59_adj_417;
    input n59_adj_418;
    output amdemod_d_11__N_2089;
    input n40_adj_419;
    input n40_adj_420;
    output amdemod_d_11__N_2092;
    input n61_adj_421;
    input n61_adj_422;
    output amdemod_d_11__N_2095;
    output amdemod_d_11__N_2098;
    output amdemod_d_11__N_2005;
    input n50_adj_423;
    input n50_adj_424;
    input n52_adj_425;
    input n52_adj_426;
    input n52_adj_427;
    input n52_adj_428;
    input n32_adj_429;
    input n32_adj_430;
    output amdemod_d_11__N_2011;
    input n47_adj_431;
    input n47_adj_432;
    input n47_adj_433;
    input n47_adj_434;
    input n49_adj_435;
    input n49_adj_436;
    input n49_adj_437;
    input n49_adj_438;
    input n44_adj_439;
    input n44_adj_440;
    output amdemod_d_11__N_2008;
    output amdemod_d_11__N_2017;
    output amdemod_d_11__N_2014;
    
    wire cic_sine_clk /* synthesis SET_AS_NETWORK=cic_sine_clk, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(86[10:22])
    wire [12:0]n1;
    wire [12:0]amdemod_d;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(30[38:47])
    
    wire n16687, n16688, n16925, n16816, n16817, amdemod_d_11__N_1829, 
        n16744, n16745, n16927, n16747, n16748, n16819, n16820, 
        n16786, n16787, n16804, n16805, n16813, n16814, n16750, 
        n16751, amdemod_d_11__N_1873, n16923, n16771, n16772, amdemod_d_11__N_1879, 
        n16811, n16810, n16808, n16807, n16802, n16801, n16799, 
        n16798, n16796, n16795, n16769, n16768, n16741, n16793, 
        n16792, n16739, n16790, n16789, n16738, n16784, n16783, 
        n16736, n16735, n16781, n16780, n16724, n16778, n16777, 
        n16723, n16721, n16720, n16718, n16717, n16715, n16726, 
        n16727, n16714, n16712, amdemod_d_11__N_1863, n16775, n16711, 
        n16774, n16709, n16730, n16729, n16708, n16706, n16705, 
        n16703, n16753, n16754, n16926, n16924, n16928, n16657, 
        n16658, n16929, n16930, n16931, n16702, n17281, n16700, 
        n16699, n16697, amdemod_d_11__N_1848, n16696, n16694, n16693, 
        amdemod_d_11__N_1868, n16691, n16690, amdemod_d_11__N_1858, 
        n16685, amdemod_d_11__N_1853, amdemod_d_11__N_1843, amdemod_d_11__N_1838, 
        amdemod_d_11__N_1833, n16684, n16763, n16762, n16682, n16765, 
        n16766, n16681, n16679, n16678, n16676, n16675, n16673, 
        n16672, n16660, n16661, n16663, n16664, n16756, n16757, 
        n16666, n16667, n16759, n16760, n16732, n16733, n16669, 
        n16670, n16822, n16823, n16837, n16838, n16825, n16826, 
        n16832, n16831, n16829, n16828, n16835, n16834, n16742;
    
    FD1S3AX mult_result_q_res2_e1__i1 (.D(cic_cosine_out[0]), .CK(cic_sine_clk), 
            .Q(n1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_e1__i1.GSR = "ENABLED";
    FD1S3AX amdemod_out_i1 (.D(amdemod_d[0]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2339[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_out_i1.GSR = "ENABLED";
    LUT4 i1464_2_lut (.A(\square_sum[22] ), .B(\square_sum[23] ), .Z(n11179)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1464_2_lut.init = 16'hbbbb;
    PFUMX i5478 (.BLUT(n16687), .ALUT(n16688), .C0(n16925), .Z(amdemod_d_11__N_1874));
    PFUMX i5607 (.BLUT(n16816), .ALUT(n16817), .C0(amdemod_d_11__N_1829), 
          .Z(amdemod_d_11__N_2023));
    PFUMX i5535 (.BLUT(n16744), .ALUT(n16745), .C0(n16927), .Z(amdemod_d_11__N_2146));
    PFUMX i5538 (.BLUT(n16747), .ALUT(n16748), .C0(n16927), .Z(amdemod_d_11__N_2149));
    PFUMX i5610 (.BLUT(n16819), .ALUT(n16820), .C0(amdemod_d_11__N_1829), 
          .Z(amdemod_d_11__N_2020));
    PFUMX i5577 (.BLUT(n16786), .ALUT(n16787), .C0(n16925), .Z(amdemod_d_11__N_2281));
    PFUMX i5595 (.BLUT(n16804), .ALUT(n16805), .C0(n16925), .Z(amdemod_d_11__N_2284));
    PFUMX i5604 (.BLUT(n16813), .ALUT(n16814), .C0(amdemod_d_11__N_1829), 
          .Z(amdemod_d_11__N_2026));
    PFUMX i5541 (.BLUT(n16750), .ALUT(n16751), .C0(n16927), .Z(amdemod_d_11__N_2152));
    LUT4 i676_2_lut_4_lut_4_lut (.A(\square_sum[21] ), .B(\square_sum[23] ), 
         .C(\square_sum[22] ), .D(\square_sum[20] ), .Z(n4)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+(C+!(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(62[20:38])
    defparam i676_2_lut_4_lut_4_lut.init = 16'hab02;
    LUT4 amdemod_d_11__I_19_1_lut (.A(amdemod_d_11__N_1874), .Z(amdemod_d_11__N_1873)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(67[34:48])
    defparam amdemod_d_11__I_19_1_lut.init = 16'h5555;
    LUT4 amdemod_d_11__I_18_rep_235_3_lut (.A(\amdemod_d_11__N_1870[13] ), 
         .B(\amdemod_d_11__N_1871[13] ), .C(n17128), .Z(n16923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_18_rep_235_3_lut.init = 16'hcaca;
    MULT18X18D mult_result_q_res2_mult_2 (.A17(n1[12]), .A16(n1[12]), .A15(n1[12]), 
            .A14(n1[12]), .A13(n1[12]), .A12(n1[12]), .A11(n1[12]), 
            .A10(n1[10]), .A9(n1[9]), .A8(n1[8]), .A7(n1[7]), .A6(n1[6]), 
            .A5(n1[5]), .A4(n1[4]), .A3(n1[3]), .A2(n1[2]), .A1(n1[1]), 
            .A0(n1[0]), .B17(n1[12]), .B16(n1[12]), .B15(n1[12]), .B14(n1[12]), 
            .B13(n1[12]), .B12(n1[12]), .B11(n1[12]), .B10(n1[10]), 
            .B9(n1[9]), .B8(n1[8]), .B7(n1[7]), .B6(n1[6]), .B5(n1[5]), 
            .B4(n1[4]), .B3(n1[3]), .B2(n1[2]), .B1(n1[1]), .B0(n1[0]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .P23(n57), .P22(n58), 
            .P21(n59), .P20(n60), .P19(n61), .P18(n62), .P17(n63), 
            .P16(n64), .P15(n65), .P14(n66), .P13(n67), .P12(n68), 
            .P11(n69), .P10(n70), .P9(n71), .P8(n72), .P7(n73), .P6(n74), 
            .P5(n75), .P4(n76), .P3(n77), .P2(n78), .P1(n79), .P0(n80));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_result_q_res2_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_result_q_res2_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_result_q_res2_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_result_q_res2_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_result_q_res2_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_result_q_res2_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_result_q_res2_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_result_q_res2_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_result_q_res2_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_result_q_res2_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_result_q_res2_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_result_q_res2_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_result_q_res2_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_result_q_res2_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_result_q_res2_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_result_q_res2_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_result_q_res2_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_result_q_res2_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_result_q_res2_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_result_q_res2_mult_2.GSR = "ENABLED";
    defparam mult_result_q_res2_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_result_q_res2_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_result_q_res2_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_result_q_res2_mult_2.RESETMODE = "SYNC";
    LUT4 square_sum_23__bdd_4_lut_5815 (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(\square_sum[20] ), .D(\square_sum[21] ), .Z(n17146)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+!(C+(D)))) */ ;
    defparam square_sum_23__bdd_4_lut_5815.init = 16'h9110;
    LUT4 i1_2_lut_rep_360 (.A(\square_sum[23] ), .B(\square_sum[22] ), .Z(n17157)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_360.init = 16'h6666;
    LUT4 i5560_3_lut (.A(n34), .B(n34_adj_225), .C(n17134), .Z(n16771)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5560_3_lut.init = 16'hcaca;
    LUT4 i5561_3_lut (.A(n32), .B(n32_adj_226), .C(n17134), .Z(n16772)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5561_3_lut.init = 16'hcaca;
    FD1S3AX amdemod_d__0_i1 (.D(amdemod_d_11__N_1879), .CK(cic_sine_clk), 
            .Q(amdemod_d[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_d__0_i1.GSR = "ENABLED";
    LUT4 i5600_3_lut (.A(n71_adj_227), .B(n71_adj_228), .C(n17134), .Z(n16811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5600_3_lut.init = 16'hcaca;
    LUT4 i5599_3_lut (.A(n73_adj_229), .B(n73_adj_230), .C(n17134), .Z(n16810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5599_3_lut.init = 16'hcaca;
    LUT4 i5597_3_lut (.A(n68_adj_231), .B(n68_adj_232), .C(n17134), .Z(n16808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5597_3_lut.init = 16'hcaca;
    LUT4 i5596_3_lut (.A(n70_adj_233), .B(n70_adj_234), .C(n17134), .Z(n16807)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5596_3_lut.init = 16'hcaca;
    LUT4 i5591_3_lut (.A(n65_adj_235), .B(n65_adj_236), .C(n17134), .Z(n16802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5591_3_lut.init = 16'hcaca;
    LUT4 i5590_3_lut (.A(n67_adj_237), .B(n67_adj_238), .C(n17134), .Z(n16801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5590_3_lut.init = 16'hcaca;
    LUT4 i5588_3_lut (.A(n62_adj_239), .B(n62_adj_240), .C(n17134), .Z(n16799)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5588_3_lut.init = 16'hcaca;
    LUT4 i5587_3_lut (.A(n64_adj_241), .B(n64_adj_242), .C(n17134), .Z(n16798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5587_3_lut.init = 16'hcaca;
    LUT4 i5585_3_lut (.A(n59_adj_243), .B(n59_adj_244), .C(n17134), .Z(n16796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5585_3_lut.init = 16'hcaca;
    LUT4 i5584_3_lut (.A(n61_adj_245), .B(n61_adj_246), .C(n17134), .Z(n16795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5584_3_lut.init = 16'hcaca;
    LUT4 i5558_3_lut (.A(n53), .B(n53_adj_247), .C(n17134), .Z(n16769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5558_3_lut.init = 16'hcaca;
    LUT4 i5557_3_lut (.A(n55), .B(n55_adj_248), .C(n17134), .Z(n16768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5557_3_lut.init = 16'hcaca;
    LUT4 i5530_3_lut (.A(n46), .B(n46_adj_249), .C(n17132), .Z(n16741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5530_3_lut.init = 16'hcaca;
    LUT4 i5582_3_lut (.A(n56), .B(n56_adj_250), .C(n17134), .Z(n16793)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5582_3_lut.init = 16'hcaca;
    LUT4 i5581_3_lut (.A(n58_adj_251), .B(n58_adj_252), .C(n17134), .Z(n16792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5581_3_lut.init = 16'hcaca;
    LUT4 i5528_3_lut (.A(n41), .B(n41_adj_253), .C(n17132), .Z(n16739)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5528_3_lut.init = 16'hcaca;
    LUT4 i5579_3_lut (.A(n50), .B(n50_adj_254), .C(n17134), .Z(n16790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5579_3_lut.init = 16'hcaca;
    LUT4 i5578_3_lut (.A(n52), .B(n52_adj_255), .C(n17134), .Z(n16789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5578_3_lut.init = 16'hcaca;
    MULT18X18D mult_result_i_e3 (.A17(mult_i_b[11]), .A16(mult_i_b[11]), 
            .A15(mult_i_b[11]), .A14(mult_i_b[11]), .A13(mult_i_b[11]), 
            .A12(mult_i_b[11]), .A11(mult_i_b[11]), .A10(mult_i_b[10]), 
            .A9(mult_i_b[9]), .A8(mult_i_b[8]), .A7(mult_i_b[7]), .A6(mult_i_b[6]), 
            .A5(mult_i_b[5]), .A4(mult_i_b[4]), .A3(mult_i_b[3]), .A2(mult_i_b[2]), 
            .A1(mult_i_b[1]), .A0(mult_i_b[0]), .B17(mult_i_b[11]), .B16(mult_i_b[11]), 
            .B15(mult_i_b[11]), .B14(mult_i_b[11]), .B13(mult_i_b[11]), 
            .B12(mult_i_b[11]), .B11(mult_i_b[11]), .B10(mult_i_b[10]), 
            .B9(mult_i_b[9]), .B8(mult_i_b[8]), .B7(mult_i_b[7]), .B6(mult_i_b[6]), 
            .B5(mult_i_b[5]), .B4(mult_i_b[4]), .B3(mult_i_b[3]), .B2(mult_i_b[2]), 
            .B1(mult_i_b[1]), .B0(mult_i_b[0]), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(cic_sine_clk), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(VCC_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .P23(mult_result_i[23]), .P22(mult_result_i[22]), .P21(mult_result_i[21]), 
            .P20(mult_result_i[20]), .P19(mult_result_i[19]), .P18(mult_result_i[18]), 
            .P17(mult_result_i[17]), .P16(mult_result_i[16]), .P15(mult_result_i[15]), 
            .P14(mult_result_i[14]), .P13(mult_result_i[13]), .P12(mult_result_i[12]), 
            .P11(mult_result_i[11]), .P10(mult_result_i[10]), .P9(mult_result_i[9]), 
            .P8(mult_result_i[8]), .P7(mult_result_i[7]), .P6(mult_result_i[6]), 
            .P5(mult_result_i[5]), .P4(mult_result_i[4]), .P3(mult_result_i[3]), 
            .P2(mult_result_i[2]), .P1(mult_result_i[1]), .P0(mult_result_i[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(86[22:41])
    defparam mult_result_i_e3.REG_INPUTA_CLK = "CLK3";
    defparam mult_result_i_e3.REG_INPUTA_CE = "CE3";
    defparam mult_result_i_e3.REG_INPUTA_RST = "RST3";
    defparam mult_result_i_e3.REG_INPUTB_CLK = "CLK3";
    defparam mult_result_i_e3.REG_INPUTB_CE = "CE3";
    defparam mult_result_i_e3.REG_INPUTB_RST = "RST3";
    defparam mult_result_i_e3.REG_INPUTC_CLK = "NONE";
    defparam mult_result_i_e3.REG_INPUTC_CE = "CE0";
    defparam mult_result_i_e3.REG_INPUTC_RST = "RST0";
    defparam mult_result_i_e3.REG_PIPELINE_CLK = "NONE";
    defparam mult_result_i_e3.REG_PIPELINE_CE = "CE0";
    defparam mult_result_i_e3.REG_PIPELINE_RST = "RST0";
    defparam mult_result_i_e3.REG_OUTPUT_CLK = "CLK3";
    defparam mult_result_i_e3.REG_OUTPUT_CE = "CE3";
    defparam mult_result_i_e3.REG_OUTPUT_RST = "RST3";
    defparam mult_result_i_e3.CLK0_DIV = "ENABLED";
    defparam mult_result_i_e3.CLK1_DIV = "ENABLED";
    defparam mult_result_i_e3.CLK2_DIV = "ENABLED";
    defparam mult_result_i_e3.CLK3_DIV = "ENABLED";
    defparam mult_result_i_e3.HIGHSPEED_CLK = "NONE";
    defparam mult_result_i_e3.GSR = "ENABLED";
    defparam mult_result_i_e3.CAS_MATCH_REG = "FALSE";
    defparam mult_result_i_e3.SOURCEB_MODE = "B_SHIFT";
    defparam mult_result_i_e3.MULT_BYPASS = "DISABLED";
    defparam mult_result_i_e3.RESETMODE = "ASYNC";
    LUT4 i5527_3_lut (.A(n43), .B(n43_adj_256), .C(n17132), .Z(n16738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5527_3_lut.init = 16'hcaca;
    LUT4 i5573_3_lut (.A(n47), .B(n47_adj_257), .C(n17134), .Z(n16784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5573_3_lut.init = 16'hcaca;
    LUT4 i5572_3_lut (.A(n49), .B(n49_adj_258), .C(n17134), .Z(n16783)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5572_3_lut.init = 16'hcaca;
    LUT4 i5525_3_lut (.A(n38), .B(n38_adj_259), .C(n17132), .Z(n16736)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5525_3_lut.init = 16'hcaca;
    LUT4 i5524_3_lut (.A(n40), .B(n40_adj_260), .C(n17132), .Z(n16735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5524_3_lut.init = 16'hcaca;
    LUT4 i5570_3_lut (.A(n44), .B(n44_adj_261), .C(n17134), .Z(n16781)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5570_3_lut.init = 16'hcaca;
    LUT4 i5569_3_lut (.A(n46_adj_262), .B(n46_adj_263), .C(n17134), .Z(n16780)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5569_3_lut.init = 16'hcaca;
    LUT4 i5513_3_lut (.A(n71_adj_264), .B(n71_adj_265), .C(n17130), .Z(n16724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5513_3_lut.init = 16'hcaca;
    LUT4 i5567_3_lut (.A(n41_adj_266), .B(n41_adj_267), .C(n17134), .Z(n16778)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5567_3_lut.init = 16'hcaca;
    LUT4 i5566_3_lut (.A(n43_adj_268), .B(n43_adj_269), .C(n17134), .Z(n16777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5566_3_lut.init = 16'hcaca;
    LUT4 i5512_3_lut (.A(n73_adj_270), .B(n73_adj_271), .C(n17130), .Z(n16723)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5512_3_lut.init = 16'hcaca;
    LUT4 i5510_3_lut (.A(n68_adj_272), .B(n68_adj_273), .C(n17130), .Z(n16721)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5510_3_lut.init = 16'hcaca;
    LUT4 i5509_3_lut (.A(n70_adj_274), .B(n70_adj_275), .C(n17130), .Z(n16720)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5509_3_lut.init = 16'hcaca;
    LUT4 i5507_3_lut (.A(n65_adj_276), .B(n65_adj_277), .C(n17130), .Z(n16718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5507_3_lut.init = 16'hcaca;
    LUT4 i5506_3_lut (.A(n67_adj_278), .B(n67_adj_279), .C(n17130), .Z(n16717)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5506_3_lut.init = 16'hcaca;
    LUT4 i5504_3_lut (.A(n62_adj_280), .B(n62_adj_281), .C(n17130), .Z(n16715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5504_3_lut.init = 16'hcaca;
    LUT4 amdemod_d_11__I_10_3_lut_rep_334 (.A(\amdemod_d_11__N_1850[13] ), 
         .B(\amdemod_d_11__N_1851[13] ), .C(n17132), .Z(n17131)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_10_3_lut_rep_334.init = 16'hcaca;
    LUT4 i5517_3_lut_rep_331 (.A(n16726), .B(n16727), .C(n17129), .Z(n17128)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5517_3_lut_rep_331.init = 16'hcaca;
    LUT4 i5503_3_lut (.A(n64_adj_282), .B(n64_adj_283), .C(n17130), .Z(n16714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5503_3_lut.init = 16'hcaca;
    LUT4 i5501_3_lut (.A(n59_adj_284), .B(n59_adj_285), .C(n17130), .Z(n16712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5501_3_lut.init = 16'hcaca;
    LUT4 amdemod_d_11__I_15_1_lut_3_lut (.A(n16726), .B(n16727), .C(n17129), 
         .Z(amdemod_d_11__N_1863)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam amdemod_d_11__I_15_1_lut_3_lut.init = 16'h3535;
    LUT4 i5564_3_lut (.A(n38_adj_286), .B(n38_adj_287), .C(n17134), .Z(n16775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5564_3_lut.init = 16'hcaca;
    LUT4 i5500_3_lut (.A(n61_adj_288), .B(n61_adj_289), .C(n17130), .Z(n16711)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5500_3_lut.init = 16'hcaca;
    LUT4 i5563_3_lut (.A(n40_adj_290), .B(n40_adj_291), .C(n17134), .Z(n16774)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5563_3_lut.init = 16'hcaca;
    LUT4 amdemod_d_11__I_22_3_lut (.A(\amdemod_d_11__N_1880[13] ), .B(\amdemod_d_11__N_1881[13] ), 
         .C(amdemod_d_11__N_1874), .Z(amdemod_d_11__N_1879)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_22_3_lut.init = 16'h3535;
    LUT4 i5498_3_lut (.A(n56_adj_292), .B(n56_adj_293), .C(n17130), .Z(n16709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5498_3_lut.init = 16'hcaca;
    LUT4 i5519_3_lut (.A(n71_adj_294), .B(n71_adj_295), .C(n17132), .Z(n16730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5519_3_lut.init = 16'hcaca;
    LUT4 i5518_3_lut (.A(n73_adj_296), .B(n73_adj_297), .C(n17132), .Z(n16729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5518_3_lut.init = 16'hcaca;
    LUT4 i5497_3_lut (.A(n58_adj_298), .B(n58_adj_299), .C(n17130), .Z(n16708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5497_3_lut.init = 16'hcaca;
    LUT4 i5495_3_lut (.A(n53_adj_300), .B(n53_adj_301), .C(n17130), .Z(n16706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5495_3_lut.init = 16'hcaca;
    LUT4 i5494_3_lut (.A(n55_adj_302), .B(n55_adj_303), .C(n17130), .Z(n16705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5494_3_lut.init = 16'hcaca;
    LUT4 i5492_3_lut (.A(n50_adj_304), .B(n50_adj_305), .C(n17130), .Z(n16703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5492_3_lut.init = 16'hcaca;
    FD1S3AX mult_result_q_res2_e1__i2 (.D(cic_cosine_out[1]), .CK(cic_sine_clk), 
            .Q(n1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_e1__i2.GSR = "ENABLED";
    FD1S3AX mult_result_q_res2_e1__i3 (.D(cic_cosine_out[2]), .CK(cic_sine_clk), 
            .Q(n1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_e1__i3.GSR = "ENABLED";
    FD1S3AX mult_result_q_res2_e1__i4 (.D(cic_cosine_out[3]), .CK(cic_sine_clk), 
            .Q(n1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_e1__i4.GSR = "ENABLED";
    FD1S3AX mult_result_q_res2_e1__i5 (.D(cic_cosine_out[4]), .CK(cic_sine_clk), 
            .Q(n1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_e1__i5.GSR = "ENABLED";
    FD1S3AX mult_result_q_res2_e1__i6 (.D(cic_cosine_out[5]), .CK(cic_sine_clk), 
            .Q(n1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_e1__i6.GSR = "ENABLED";
    FD1S3AX mult_result_q_res2_e1__i7 (.D(cic_cosine_out[6]), .CK(cic_sine_clk), 
            .Q(n1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_e1__i7.GSR = "ENABLED";
    FD1S3AX mult_result_q_res2_e1__i8 (.D(cic_cosine_out[7]), .CK(cic_sine_clk), 
            .Q(n1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_e1__i8.GSR = "ENABLED";
    FD1S3AX mult_result_q_res2_e1__i9 (.D(cic_cosine_out[8]), .CK(cic_sine_clk), 
            .Q(n1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_e1__i9.GSR = "ENABLED";
    FD1S3AX mult_result_q_res2_e1__i10 (.D(cic_cosine_out[9]), .CK(cic_sine_clk), 
            .Q(n1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_e1__i10.GSR = "ENABLED";
    FD1S3AX mult_result_q_res2_e1__i11 (.D(cic_cosine_out[10]), .CK(cic_sine_clk), 
            .Q(n1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_e1__i11.GSR = "ENABLED";
    FD1S3AX mult_result_q_res2_e1__i12 (.D(cic_cosine_out[11]), .CK(cic_sine_clk), 
            .Q(n1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(87[22:41])
    defparam mult_result_q_res2_e1__i12.GSR = "ENABLED";
    LUT4 i5476_3_lut (.A(n34_adj_306), .B(n34_adj_307), .C(n17128), .Z(n16687)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5476_3_lut.init = 16'hcaca;
    PFUMX i5544 (.BLUT(n16753), .ALUT(n16754), .C0(n16927), .Z(amdemod_d_11__N_2155));
    FD1S3AX amdemod_out_i2 (.D(amdemod_d[1]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2339[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_out_i2.GSR = "ENABLED";
    LUT4 amdemod_d_11__I_10_rep_238_3_lut (.A(\amdemod_d_11__N_1850[13] ), 
         .B(\amdemod_d_11__N_1851[13] ), .C(n17132), .Z(n16926)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_10_rep_238_3_lut.init = 16'hcaca;
    FD1S3AX amdemod_out_i3 (.D(amdemod_d[2]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2339[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_out_i3.GSR = "ENABLED";
    FD1S3AX amdemod_out_i4 (.D(amdemod_d[3]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2339[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_out_i4.GSR = "ENABLED";
    FD1S3AX amdemod_out_i5 (.D(amdemod_d[4]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2339[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_out_i5.GSR = "ENABLED";
    FD1S3AX amdemod_out_i6 (.D(amdemod_d[5]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2339[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_out_i6.GSR = "ENABLED";
    FD1S3AX amdemod_out_i7 (.D(amdemod_d[6]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2339[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_out_i7.GSR = "ENABLED";
    FD1S3AX amdemod_out_i8 (.D(amdemod_d[7]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2339[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_out_i8.GSR = "ENABLED";
    FD1S3AX amdemod_out_i9 (.D(amdemod_d[8]), .CK(cic_sine_clk), .Q(\data_in_reg_11__N_2339[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_out_i9.GSR = "ENABLED";
    FD1S3AX amdemod_out_i10 (.D(amdemod_d[9]), .CK(cic_sine_clk), .Q(\amdemod_out[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=184, LSE_RLINE=189 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_out_i10.GSR = "ENABLED";
    LUT4 amdemod_d_11__I_18_rep_236_3_lut (.A(\amdemod_d_11__N_1870[13] ), 
         .B(\amdemod_d_11__N_1871[13] ), .C(n17128), .Z(n16924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_18_rep_236_3_lut.init = 16'hcaca;
    LUT4 amdemod_d_11__I_14_rep_240_3_lut (.A(\amdemod_d_11__N_1860[13] ), 
         .B(\amdemod_d_11__N_1861[13] ), .C(n17130), .Z(n16928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_14_rep_240_3_lut.init = 16'hcaca;
    PFUMX i5448 (.BLUT(n16657), .ALUT(n16658), .C0(n17127), .Z(amdemod_d_11__N_2287));
    LUT4 amdemod_d_11__I_14_rep_241_3_lut (.A(\amdemod_d_11__N_1860[13] ), 
         .B(\amdemod_d_11__N_1861[13] ), .C(n17130), .Z(n16929)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_14_rep_241_3_lut.init = 16'hcaca;
    LUT4 amdemod_d_11__I_6_rep_242_3_lut (.A(\amdemod_d_11__N_1840[11] ), 
         .B(\amdemod_d_11__N_1841[11] ), .C(n17134), .Z(n16930)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_6_rep_242_3_lut.init = 16'hcaca;
    LUT4 amdemod_d_11__I_6_rep_243_3_lut (.A(\amdemod_d_11__N_1840[11] ), 
         .B(\amdemod_d_11__N_1841[11] ), .C(n17134), .Z(n16931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_6_rep_243_3_lut.init = 16'hcaca;
    LUT4 i5491_3_lut (.A(n52_adj_308), .B(n52_adj_309), .C(n17130), .Z(n16702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5491_3_lut.init = 16'hcaca;
    LUT4 i11_3_lut_rep_340_4_lut_4_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n17281), .D(n17163), .Z(n17137)) /* synthesis lut_function=(A (B+!(C))+!A !(B (C)+!B !(D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i11_3_lut_rep_340_4_lut_4_lut_4_lut.init = 16'h9f8e;
    LUT4 i5489_3_lut (.A(n47_adj_310), .B(n47_adj_311), .C(n17130), .Z(n16700)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5489_3_lut.init = 16'hcaca;
    LUT4 i5488_3_lut (.A(n49_adj_312), .B(n49_adj_313), .C(n17130), .Z(n16699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5488_3_lut.init = 16'hcaca;
    LUT4 i5486_3_lut (.A(n44_adj_314), .B(n44_adj_315), .C(n17130), .Z(n16697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5486_3_lut.init = 16'hcaca;
    LUT4 amdemod_d_11__I_9_1_lut_3_lut (.A(\amdemod_d_11__N_1850[13] ), .B(\amdemod_d_11__N_1851[13] ), 
         .C(n17132), .Z(amdemod_d_11__N_1848)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_9_1_lut_3_lut.init = 16'h3535;
    LUT4 amdemod_d_11__I_14_rep_332 (.A(\amdemod_d_11__N_1860[13] ), .B(\amdemod_d_11__N_1861[13] ), 
         .C(n17130), .Z(n17129)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_14_rep_332.init = 16'hcaca;
    LUT4 i5485_3_lut (.A(n46_adj_316), .B(n46_adj_317), .C(n17130), .Z(n16696)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5485_3_lut.init = 16'hcaca;
    LUT4 i2582_1_lut_3_lut_4_lut_4_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n17281), .D(n17163), .Z(amdemod_d_11__N_1829)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)+!B !(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i2582_1_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h6071;
    LUT4 i5483_3_lut (.A(n41_adj_318), .B(n41_adj_319), .C(n17130), .Z(n16694)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5483_3_lut.init = 16'hcaca;
    LUT4 i5482_3_lut (.A(n43_adj_320), .B(n43_adj_321), .C(n17130), .Z(n16693)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5482_3_lut.init = 16'hcaca;
    LUT4 amdemod_d_11__I_17_1_lut_3_lut (.A(\amdemod_d_11__N_1870[13] ), .B(\amdemod_d_11__N_1871[13] ), 
         .C(n17128), .Z(amdemod_d_11__N_1868)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_17_1_lut_3_lut.init = 16'h3535;
    LUT4 i5480_3_lut (.A(n38_adj_322), .B(n38_adj_323), .C(n17130), .Z(n16691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5480_3_lut.init = 16'hcaca;
    LUT4 i5479_3_lut (.A(n40_adj_324), .B(n40_adj_325), .C(n17130), .Z(n16690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5479_3_lut.init = 16'hcaca;
    LUT4 i5562_3_lut_rep_335 (.A(n16771), .B(n16772), .C(n17133), .Z(n17132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5562_3_lut_rep_335.init = 16'hcaca;
    LUT4 amdemod_d_11__I_13_1_lut_3_lut (.A(\amdemod_d_11__N_1860[13] ), .B(\amdemod_d_11__N_1861[13] ), 
         .C(n17130), .Z(amdemod_d_11__N_1858)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_13_1_lut_3_lut.init = 16'h3535;
    FD1S3AX amdemod_d__0_i2 (.D(amdemod_d_11__N_1873), .CK(cic_sine_clk), 
            .Q(amdemod_d[1]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_d__0_i2.GSR = "ENABLED";
    LUT4 i5474_3_lut (.A(n71_adj_326), .B(n71_adj_327), .C(n17128), .Z(n16685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5474_3_lut.init = 16'hcaca;
    FD1S3AX amdemod_d__0_i3 (.D(amdemod_d_11__N_1868), .CK(cic_sine_clk), 
            .Q(amdemod_d[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_d__0_i3.GSR = "ENABLED";
    FD1S3AX amdemod_d__0_i4 (.D(amdemod_d_11__N_1863), .CK(cic_sine_clk), 
            .Q(amdemod_d[3]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_d__0_i4.GSR = "ENABLED";
    FD1S3AX amdemod_d__0_i5 (.D(amdemod_d_11__N_1858), .CK(cic_sine_clk), 
            .Q(amdemod_d[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_d__0_i5.GSR = "ENABLED";
    FD1S3AX amdemod_d__0_i6 (.D(amdemod_d_11__N_1853), .CK(cic_sine_clk), 
            .Q(amdemod_d[5]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_d__0_i6.GSR = "ENABLED";
    FD1S3AX amdemod_d__0_i7 (.D(amdemod_d_11__N_1848), .CK(cic_sine_clk), 
            .Q(amdemod_d[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_d__0_i7.GSR = "ENABLED";
    FD1S3AX amdemod_d__0_i8 (.D(amdemod_d_11__N_1843), .CK(cic_sine_clk), 
            .Q(amdemod_d[7]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_d__0_i8.GSR = "ENABLED";
    FD1S3AX amdemod_d__0_i9 (.D(amdemod_d_11__N_1838), .CK(cic_sine_clk), 
            .Q(amdemod_d[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_d__0_i9.GSR = "ENABLED";
    FD1S3AX amdemod_d__0_i10 (.D(amdemod_d_11__N_1833), .CK(cic_sine_clk), 
            .Q(amdemod_d[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(78[10] 97[6])
    defparam amdemod_d__0_i10.GSR = "ENABLED";
    LUT4 i5473_3_lut (.A(n73_adj_328), .B(n73_adj_329), .C(n17128), .Z(n16684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5473_3_lut.init = 16'hcaca;
    LUT4 i5552_3_lut (.A(n65_adj_330), .B(n65_adj_331), .C(n17132), .Z(n16763)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5552_3_lut.init = 16'hcaca;
    LUT4 i5551_3_lut (.A(n67_adj_332), .B(n67_adj_333), .C(n17132), .Z(n16762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5551_3_lut.init = 16'hcaca;
    LUT4 i5471_3_lut (.A(n68_adj_334), .B(n68_adj_335), .C(n17128), .Z(n16682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5471_3_lut.init = 16'hcaca;
    LUT4 amdemod_d_11__I_7_1_lut_3_lut (.A(n16771), .B(n16772), .C(n17133), 
         .Z(amdemod_d_11__N_1843)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam amdemod_d_11__I_7_1_lut_3_lut.init = 16'h3535;
    LUT4 i5556_3_lut_rep_333 (.A(n16765), .B(n16766), .C(n17131), .Z(n17130)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5556_3_lut_rep_333.init = 16'hcaca;
    LUT4 i5470_3_lut (.A(n70_adj_336), .B(n70_adj_337), .C(n17128), .Z(n16681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5470_3_lut.init = 16'hcaca;
    LUT4 i5468_3_lut (.A(n65_adj_338), .B(n65_adj_339), .C(n17128), .Z(n16679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5468_3_lut.init = 16'hcaca;
    LUT4 i5467_3_lut (.A(n67_adj_340), .B(n67_adj_341), .C(n17128), .Z(n16678)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5467_3_lut.init = 16'hcaca;
    LUT4 i5465_3_lut (.A(n62_adj_342), .B(n62_adj_343), .C(n17128), .Z(n16676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5465_3_lut.init = 16'hcaca;
    LUT4 i5464_3_lut (.A(n64_adj_344), .B(n64_adj_345), .C(n17128), .Z(n16675)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5464_3_lut.init = 16'hcaca;
    LUT4 i5462_3_lut (.A(n59_adj_346), .B(n59_adj_347), .C(n17128), .Z(n16673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5462_3_lut.init = 16'hcaca;
    LUT4 i5461_3_lut (.A(n61_adj_348), .B(n61_adj_349), .C(n17128), .Z(n16672)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5461_3_lut.init = 16'hcaca;
    PFUMX i5451 (.BLUT(n16660), .ALUT(n16661), .C0(n16923), .Z(amdemod_d_11__N_2290));
    PFUMX i5454 (.BLUT(n16663), .ALUT(n16664), .C0(n16923), .Z(amdemod_d_11__N_2293));
    PFUMX i5547 (.BLUT(n16756), .ALUT(n16757), .C0(n17131), .Z(amdemod_d_11__N_2158));
    PFUMX i5457 (.BLUT(n16666), .ALUT(n16667), .C0(n16923), .Z(amdemod_d_11__N_2296));
    PFUMX i5550 (.BLUT(n16759), .ALUT(n16760), .C0(n17131), .Z(amdemod_d_11__N_2161));
    LUT4 i5543_3_lut (.A(n56_adj_350), .B(n56_adj_351), .C(n17132), .Z(n16754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5543_3_lut.init = 16'hcaca;
    PFUMX i5523 (.BLUT(n16732), .ALUT(n16733), .C0(n16926), .Z(amdemod_d_11__N_2167));
    PFUMX i5460 (.BLUT(n16669), .ALUT(n16670), .C0(n16923), .Z(amdemod_d_11__N_2299));
    LUT4 i5515_3_lut (.A(n34_adj_352), .B(n34_adj_353), .C(n17130), .Z(n16726)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5515_3_lut.init = 16'hcaca;
    LUT4 i5522_3_lut (.A(n68_adj_354), .B(n68_adj_355), .C(n17132), .Z(n16733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5522_3_lut.init = 16'hcaca;
    LUT4 i719_2_lut_rep_365 (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .Z(n17162)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i719_2_lut_rep_365.init = 16'heeee;
    PFUMX i5463 (.BLUT(n16672), .ALUT(n16673), .C0(n16924), .Z(amdemod_d_11__N_2302));
    PFUMX i5553 (.BLUT(n16762), .ALUT(n16763), .C0(n17131), .Z(amdemod_d_11__N_2164));
    LUT4 i5542_3_lut (.A(n58_adj_356), .B(n58_adj_357), .C(n17132), .Z(n16753)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5542_3_lut.init = 16'hcaca;
    LUT4 i5611_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n39), .D(n39_adj_358), .Z(n16822)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5611_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5612_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n52_adj_441[3]), .D(n52_adj_442[3]), .Z(n16823)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5612_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5447_3_lut (.A(n44_adj_372), .B(n44_adj_373), .C(n17128), .Z(n16658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5447_3_lut.init = 16'hcaca;
    LUT4 i5446_3_lut (.A(n46_adj_374), .B(n46_adj_375), .C(n17128), .Z(n16657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5446_3_lut.init = 16'hcaca;
    LUT4 i5516_3_lut (.A(n32_adj_376), .B(n32_adj_377), .C(n17130), .Z(n16727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5516_3_lut.init = 16'hcaca;
    PFUMX i5466 (.BLUT(n16675), .ALUT(n16676), .C0(n16924), .Z(amdemod_d_11__N_2305));
    LUT4 amdemod_d_11__I_5_1_lut_3_lut (.A(\amdemod_d_11__N_1840[11] ), .B(\amdemod_d_11__N_1841[11] ), 
         .C(n17134), .Z(amdemod_d_11__N_1838)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_5_1_lut_3_lut.init = 16'h3535;
    LUT4 i5628_3_lut_rep_337 (.A(n16837), .B(n16838), .C(n17137), .Z(n17134)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i5628_3_lut_rep_337.init = 16'hacac;
    LUT4 i5521_3_lut (.A(n70_adj_378), .B(n70_adj_379), .C(n17132), .Z(n16732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5521_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), .C(\square_sum[21] ), 
         .D(\square_sum[20] ), .Z(\amdemod_d_11__N_1830[1] )) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i1_3_lut_4_lut.init = 16'he11e;
    LUT4 i5554_3_lut (.A(n34_adj_380), .B(n34_adj_381), .C(n17132), .Z(n16765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5554_3_lut.init = 16'hcaca;
    LUT4 i5555_3_lut (.A(n32_adj_382), .B(n32_adj_383), .C(n17132), .Z(n16766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5555_3_lut.init = 16'hcaca;
    LUT4 amdemod_d_11__I_18_rep_237_3_lut (.A(\amdemod_d_11__N_1870[13] ), 
         .B(\amdemod_d_11__N_1871[13] ), .C(n17128), .Z(n16925)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_18_rep_237_3_lut.init = 16'hcaca;
    LUT4 i5602_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n48), .D(n48_adj_384), .Z(n16813)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5602_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5540_3_lut (.A(n53_adj_385), .B(n53_adj_386), .C(n17132), .Z(n16751)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5540_3_lut.init = 16'hcaca;
    PFUMX i5469 (.BLUT(n16678), .ALUT(n16679), .C0(n16924), .Z(amdemod_d_11__N_2308));
    LUT4 i5603_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n52_adj_441[0]), .D(n52_adj_442[0]), .Z(n16814)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5603_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i5472 (.BLUT(n16681), .ALUT(n16682), .C0(n16924), .Z(amdemod_d_11__N_2311));
    LUT4 i5594_3_lut (.A(n41_adj_387), .B(n41_adj_388), .C(n17128), .Z(n16805)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5594_3_lut.init = 16'hcaca;
    LUT4 i5614_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n36), .D(n36_adj_389), .Z(n16825)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5614_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5608_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n42), .D(n42_adj_390), .Z(n16819)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5608_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i5475 (.BLUT(n16684), .ALUT(n16685), .C0(n16925), .Z(amdemod_d_11__N_2314));
    PFUMX i5481 (.BLUT(n16690), .ALUT(n16691), .C0(n17129), .Z(amdemod_d_11__N_2209));
    LUT4 i5627_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n52_adj_441[8]), .D(n52_adj_442[8]), .Z(n16838)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5627_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5609_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n52_adj_441[2]), .D(n52_adj_442[2]), .Z(n16820)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5609_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i5520 (.BLUT(n16729), .ALUT(n16730), .C0(n17131), .Z(amdemod_d_11__N_2170));
    LUT4 i5606_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n52_adj_441[1]), .D(n52_adj_442[1]), .Z(n16817)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5606_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5615_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n52_adj_441[4]), .D(n52_adj_442[4]), .Z(n16826)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5615_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5626_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n24), .D(n24_adj_391), .Z(n16837)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5626_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i5484 (.BLUT(n16693), .ALUT(n16694), .C0(n16928), .Z(amdemod_d_11__N_2212));
    LUT4 i5621_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n52_adj_441[6]), .D(n52_adj_442[6]), .Z(n16832)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5621_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5605_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n45), .D(n45_adj_392), .Z(n16816)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5605_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5620_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n30), .D(n30_adj_393), .Z(n16831)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5620_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5618_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n52_adj_441[5]), .D(n52_adj_442[5]), .Z(n16829)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5618_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5617_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n33), .D(n33_adj_394), .Z(n16828)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5617_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i5487 (.BLUT(n16696), .ALUT(n16697), .C0(n16928), .Z(amdemod_d_11__N_2215));
    LUT4 i5624_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n52_adj_441[7]), .D(n52_adj_442[7]), .Z(n16835)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5624_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5623_3_lut_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(n27), .D(n27_adj_395), .Z(n16834)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i5623_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i5490 (.BLUT(n16699), .ALUT(n16700), .C0(n16928), .Z(amdemod_d_11__N_2218));
    LUT4 amdemod_d_11__I_10_rep_239_3_lut (.A(\amdemod_d_11__N_1850[13] ), 
         .B(\amdemod_d_11__N_1851[13] ), .C(n17132), .Z(n16927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_10_rep_239_3_lut.init = 16'hcaca;
    PFUMX i5493 (.BLUT(n16702), .ALUT(n16703), .C0(n16928), .Z(amdemod_d_11__N_2221));
    LUT4 amdemod_d_11__I_3_1_lut_3_lut (.A(n16837), .B(n16838), .C(n17137), 
         .Z(amdemod_d_11__N_1833)) /* synthesis lut_function=(!(A (B+(C))+!A !((C)+!B))) */ ;
    defparam amdemod_d_11__I_3_1_lut_3_lut.init = 16'h5353;
    PFUMX i5496 (.BLUT(n16705), .ALUT(n16706), .C0(n16929), .Z(amdemod_d_11__N_2224));
    LUT4 i5459_3_lut (.A(n56_adj_396), .B(n56_adj_397), .C(n17128), .Z(n16670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5459_3_lut.init = 16'hcaca;
    PFUMX i5499 (.BLUT(n16708), .ALUT(n16709), .C0(n16929), .Z(amdemod_d_11__N_2227));
    PFUMX i5502 (.BLUT(n16711), .ALUT(n16712), .C0(n16929), .Z(amdemod_d_11__N_2230));
    LUT4 square_sum_23__bdd_4_lut (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(\square_sum[20] ), .D(\square_sum[21] ), .Z(n6)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B))) */ ;
    defparam square_sum_23__bdd_4_lut.init = 16'h3331;
    PFUMX i5565 (.BLUT(n16774), .ALUT(n16775), .C0(n16930), .Z(amdemod_d_11__N_2065));
    LUT4 amdemod_d_11__I_18_rep_330 (.A(\amdemod_d_11__N_1870[13] ), .B(\amdemod_d_11__N_1871[13] ), 
         .C(n17128), .Z(n17127)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_18_rep_330.init = 16'hcaca;
    PFUMX i5505 (.BLUT(n16714), .ALUT(n16715), .C0(n16929), .Z(amdemod_d_11__N_2233));
    LUT4 i5458_3_lut (.A(n58_adj_398), .B(n58_adj_399), .C(n17128), .Z(n16669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5458_3_lut.init = 16'hcaca;
    PFUMX i5508 (.BLUT(n16717), .ALUT(n16718), .C0(n17129), .Z(amdemod_d_11__N_2236));
    PFUMX i5568 (.BLUT(n16777), .ALUT(n16778), .C0(n16930), .Z(amdemod_d_11__N_2068));
    PFUMX i5511 (.BLUT(n16720), .ALUT(n16721), .C0(n17129), .Z(amdemod_d_11__N_2239));
    LUT4 i1_3_lut_4_lut_4_lut_rep_368_4_lut (.A(\square_sum[22] ), .B(\square_sum[23] ), 
         .C(\square_sum[20] ), .D(\square_sum[21] ), .Z(n17279)) /* synthesis lut_function=(A (B)+!A ((C+(D))+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i1_3_lut_4_lut_4_lut_rep_368_4_lut.init = 16'hddd9;
    LUT4 square_sum_23__bdd_4_lut_5868 (.A(\square_sum[23] ), .B(\square_sum[22] ), 
         .C(\square_sum[20] ), .D(\square_sum[21] ), .Z(n17163)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B (C (D))+!B (C+(D)))) */ ;
    defparam square_sum_23__bdd_4_lut_5868.init = 16'hf332;
    PFUMX i5514 (.BLUT(n16723), .ALUT(n16724), .C0(n17129), .Z(amdemod_d_11__N_2242));
    LUT4 i5456_3_lut (.A(n53_adj_400), .B(n53_adj_401), .C(n17128), .Z(n16667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5456_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_4_lut (.A(\square_sum[21] ), .B(\square_sum[23] ), 
         .C(\square_sum[22] ), .D(\square_sum[20] ), .Z(n4_adj_402)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i1_4_lut_4_lut_4_lut.init = 16'h0e58;
    PFUMX i5571 (.BLUT(n16780), .ALUT(n16781), .C0(n16930), .Z(amdemod_d_11__N_2071));
    PFUMX i5526 (.BLUT(n16735), .ALUT(n16736), .C0(n16926), .Z(amdemod_d_11__N_2137));
    PFUMX i5574 (.BLUT(n16783), .ALUT(n16784), .C0(n16930), .Z(amdemod_d_11__N_2074));
    LUT4 i5549_3_lut (.A(n62_adj_403), .B(n62_adj_404), .C(n17132), .Z(n16760)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5549_3_lut.init = 16'hcaca;
    LUT4 i5548_3_lut (.A(n64_adj_405), .B(n64_adj_406), .C(n17132), .Z(n16759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5548_3_lut.init = 16'hcaca;
    PFUMX i5529 (.BLUT(n16738), .ALUT(n16739), .C0(n16926), .Z(amdemod_d_11__N_2140));
    LUT4 amdemod_d_11__I_6_rep_336 (.A(\amdemod_d_11__N_1840[11] ), .B(\amdemod_d_11__N_1841[11] ), 
         .C(n17134), .Z(n17133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(63[18] 65[12])
    defparam amdemod_d_11__I_6_rep_336.init = 16'hcaca;
    PFUMX i5580 (.BLUT(n16789), .ALUT(n16790), .C0(n16931), .Z(amdemod_d_11__N_2077));
    LUT4 i5593_3_lut (.A(n43_adj_407), .B(n43_adj_408), .C(n17128), .Z(n16804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5593_3_lut.init = 16'hcaca;
    LUT4 i5539_3_lut (.A(n55_adj_409), .B(n55_adj_410), .C(n17132), .Z(n16750)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5539_3_lut.init = 16'hcaca;
    LUT4 i5537_3_lut (.A(n50_adj_411), .B(n50_adj_412), .C(n17132), .Z(n16748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5537_3_lut.init = 16'hcaca;
    PFUMX i5532 (.BLUT(n16741), .ALUT(n16742), .C0(n16926), .Z(amdemod_d_11__N_2143));
    PFUMX i5583 (.BLUT(n16792), .ALUT(n16793), .C0(n16931), .Z(amdemod_d_11__N_2083));
    PFUMX i5559 (.BLUT(n16768), .ALUT(n16769), .C0(n17133), .Z(amdemod_d_11__N_2080));
    LUT4 amdemod_d_11__I_11_1_lut_3_lut (.A(n16765), .B(n16766), .C(n17131), 
         .Z(amdemod_d_11__N_1853)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam amdemod_d_11__I_11_1_lut_3_lut.init = 16'h3535;
    LUT4 i5455_3_lut (.A(n55_adj_413), .B(n55_adj_414), .C(n17128), .Z(n16666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5455_3_lut.init = 16'hcaca;
    LUT4 i1_rep_370 (.A(\square_sum[22] ), .B(\square_sum[23] ), .C(\square_sum[20] ), 
         .D(\square_sum[21] ), .Z(n17281)) /* synthesis lut_function=(A+!((C+(D))+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/AMDemod.v(64[20:38])
    defparam i1_rep_370.init = 16'haaae;
    PFUMX i5586 (.BLUT(n16795), .ALUT(n16796), .C0(n16931), .Z(amdemod_d_11__N_2086));
    LUT4 i5576_3_lut (.A(n38_adj_415), .B(n38_adj_416), .C(n17128), .Z(n16787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5576_3_lut.init = 16'hcaca;
    LUT4 i5546_3_lut (.A(n59_adj_417), .B(n59_adj_418), .C(n17132), .Z(n16757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5546_3_lut.init = 16'hcaca;
    PFUMX i5589 (.BLUT(n16798), .ALUT(n16799), .C0(n16931), .Z(amdemod_d_11__N_2089));
    LUT4 i5575_3_lut (.A(n40_adj_419), .B(n40_adj_420), .C(n17128), .Z(n16786)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5575_3_lut.init = 16'hcaca;
    PFUMX i5592 (.BLUT(n16801), .ALUT(n16802), .C0(n17133), .Z(amdemod_d_11__N_2092));
    LUT4 i5545_3_lut (.A(n61_adj_421), .B(n61_adj_422), .C(n17132), .Z(n16756)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5545_3_lut.init = 16'hcaca;
    PFUMX i5598 (.BLUT(n16807), .ALUT(n16808), .C0(n17133), .Z(amdemod_d_11__N_2095));
    PFUMX i5601 (.BLUT(n16810), .ALUT(n16811), .C0(n17133), .Z(amdemod_d_11__N_2098));
    PFUMX i5625 (.BLUT(n16834), .ALUT(n16835), .C0(amdemod_d_11__N_1829), 
          .Z(amdemod_d_11__N_2005));
    LUT4 i5453_3_lut (.A(n50_adj_423), .B(n50_adj_424), .C(n17128), .Z(n16664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5453_3_lut.init = 16'hcaca;
    LUT4 i5452_3_lut (.A(n52_adj_425), .B(n52_adj_426), .C(n17128), .Z(n16663)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5452_3_lut.init = 16'hcaca;
    LUT4 i5536_3_lut (.A(n52_adj_427), .B(n52_adj_428), .C(n17132), .Z(n16747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5536_3_lut.init = 16'hcaca;
    LUT4 i5477_3_lut (.A(n32_adj_429), .B(n32_adj_430), .C(n17128), .Z(n16688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5477_3_lut.init = 16'hcaca;
    PFUMX i5619 (.BLUT(n16828), .ALUT(n16829), .C0(amdemod_d_11__N_1829), 
          .Z(amdemod_d_11__N_2011));
    LUT4 i5534_3_lut (.A(n47_adj_431), .B(n47_adj_432), .C(n17132), .Z(n16745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5534_3_lut.init = 16'hcaca;
    LUT4 i5450_3_lut (.A(n47_adj_433), .B(n47_adj_434), .C(n17128), .Z(n16661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5450_3_lut.init = 16'hcaca;
    LUT4 i5533_3_lut (.A(n49_adj_435), .B(n49_adj_436), .C(n17132), .Z(n16744)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5533_3_lut.init = 16'hcaca;
    LUT4 i5449_3_lut (.A(n49_adj_437), .B(n49_adj_438), .C(n17128), .Z(n16660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5449_3_lut.init = 16'hcaca;
    LUT4 i5531_3_lut (.A(n44_adj_439), .B(n44_adj_440), .C(n17132), .Z(n16742)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5531_3_lut.init = 16'hcaca;
    PFUMX i5622 (.BLUT(n16831), .ALUT(n16832), .C0(amdemod_d_11__N_1829), 
          .Z(amdemod_d_11__N_2008));
    PFUMX i5613 (.BLUT(n16822), .ALUT(n16823), .C0(amdemod_d_11__N_1829), 
          .Z(amdemod_d_11__N_2017));
    PFUMX i5616 (.BLUT(n16825), .ALUT(n16826), .C0(amdemod_d_11__N_1829), 
          .Z(amdemod_d_11__N_2014));
    
endmodule
//
// Verilog Description of module PLL
//

module PLL (clk_25mhz_c, clk_80mhz, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk_25mhz_c;
    output clk_80mhz;
    input GND_net;
    
    wire clk_25mhz_c /* synthesis is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(39[16:25])
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(64[10:19])
    
    EHXPLLL PLLInst_0 (.CLKI(clk_25mhz_c), .CLKFB(clk_80mhz), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .PHASELOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .CLKOP(clk_80mhz)) /* synthesis FREQUENCY_PIN_CLKOP="83.333333", FREQUENCY_PIN_CLKI="25.000000", ICP_CURRENT="5", LPF_RESISTOR="16", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=102, LSE_RLINE=105 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(102[9] 105[6])
    defparam PLLInst_0.CLKI_DIV = 3;
    defparam PLLInst_0.CLKFB_DIV = 10;
    defparam PLLInst_0.CLKOP_DIV = 7;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 6;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.CLKOP_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.PLL_LOCK_DELAY = 200;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.REFIN_RESET = "DISABLED";
    defparam PLLInst_0.SYNC_ENABLE = "DISABLED";
    defparam PLLInst_0.INT_LOCK_STICKY = "ENABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module Mixer
//

module Mixer (mix_sinewave, clk_80mhz, diff_out_c, mix_cosinewave, rf_in_c, 
            \lo_cosinewave[10] , cosinewave_out_11__N_250, \lo_sinewave[4] , 
            sinewave_out_11__N_236, \lo_cosinewave[11] , \lo_sinewave[5] , 
            \lo_sinewave[6] , \lo_cosinewave[1] , \lo_sinewave[7] , \lo_sinewave[8] , 
            \lo_sinewave[9] , \lo_sinewave[10] , \lo_sinewave[11] , \lo_sinewave[12] , 
            \lo_cosinewave[2] , \lo_cosinewave[3] , \lo_cosinewave[4] , 
            \lo_cosinewave[5] , \lo_cosinewave[6] , \lo_cosinewave[12] , 
            \lo_cosinewave[7] , \lo_cosinewave[8] , \lo_sinewave[2] , 
            \lo_sinewave[1] , \lo_cosinewave[9] , \lo_sinewave[3] ) /* synthesis syn_module_defined=1 */ ;
    output [11:0]mix_sinewave;
    input clk_80mhz;
    output diff_out_c;
    output [11:0]mix_cosinewave;
    input rf_in_c;
    input \lo_cosinewave[10] ;
    input [11:0]cosinewave_out_11__N_250;
    input \lo_sinewave[4] ;
    input [11:0]sinewave_out_11__N_236;
    input \lo_cosinewave[11] ;
    input \lo_sinewave[5] ;
    input \lo_sinewave[6] ;
    input \lo_cosinewave[1] ;
    input \lo_sinewave[7] ;
    input \lo_sinewave[8] ;
    input \lo_sinewave[9] ;
    input \lo_sinewave[10] ;
    input \lo_sinewave[11] ;
    input \lo_sinewave[12] ;
    input \lo_cosinewave[2] ;
    input \lo_cosinewave[3] ;
    input \lo_cosinewave[4] ;
    input \lo_cosinewave[5] ;
    input \lo_cosinewave[6] ;
    input \lo_cosinewave[12] ;
    input \lo_cosinewave[7] ;
    input \lo_cosinewave[8] ;
    input \lo_sinewave[2] ;
    input \lo_sinewave[1] ;
    input \lo_cosinewave[9] ;
    input \lo_sinewave[3] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(64[10:19])
    wire [11:0]sinewave_out_11__N_212;
    
    wire rf_in_delayed_2;
    wire [11:0]cosinewave_out_11__N_224;
    
    FD1S3AX sinewave_out_i0 (.D(sinewave_out_11__N_212[0]), .CK(clk_80mhz), 
            .Q(mix_sinewave[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam sinewave_out_i0.GSR = "ENABLED";
    FD1S3AY rf_in_delayed_2_14 (.D(diff_out_c), .CK(clk_80mhz), .Q(rf_in_delayed_2)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(34[10] 37[6])
    defparam rf_in_delayed_2_14.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i0 (.D(cosinewave_out_11__N_224[0]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam cosinewave_out_i0.GSR = "ENABLED";
    FD1S3AY rf_in_delayed_1_13 (.D(rf_in_c), .CK(clk_80mhz), .Q(diff_out_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(34[10] 37[6])
    defparam rf_in_delayed_1_13.GSR = "ENABLED";
    LUT4 cosinewave_out_11__I_0_i10_3_lut (.A(\lo_cosinewave[10] ), .B(cosinewave_out_11__N_250[9]), 
         .C(rf_in_delayed_2), .Z(cosinewave_out_11__N_224[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam cosinewave_out_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 sinewave_out_11__I_0_i4_3_lut (.A(\lo_sinewave[4] ), .B(sinewave_out_11__N_236[3]), 
         .C(rf_in_delayed_2), .Z(sinewave_out_11__N_212[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam sinewave_out_11__I_0_i4_3_lut.init = 16'hcaca;
    FD1S3AX sinewave_out_i1 (.D(sinewave_out_11__N_212[1]), .CK(clk_80mhz), 
            .Q(mix_sinewave[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam sinewave_out_i1.GSR = "ENABLED";
    FD1S3AX sinewave_out_i2 (.D(sinewave_out_11__N_212[2]), .CK(clk_80mhz), 
            .Q(mix_sinewave[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam sinewave_out_i2.GSR = "ENABLED";
    FD1S3AX sinewave_out_i3 (.D(sinewave_out_11__N_212[3]), .CK(clk_80mhz), 
            .Q(mix_sinewave[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam sinewave_out_i3.GSR = "ENABLED";
    FD1S3AX sinewave_out_i4 (.D(sinewave_out_11__N_212[4]), .CK(clk_80mhz), 
            .Q(mix_sinewave[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam sinewave_out_i4.GSR = "ENABLED";
    FD1S3AX sinewave_out_i5 (.D(sinewave_out_11__N_212[5]), .CK(clk_80mhz), 
            .Q(mix_sinewave[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam sinewave_out_i5.GSR = "ENABLED";
    FD1S3AX sinewave_out_i6 (.D(sinewave_out_11__N_212[6]), .CK(clk_80mhz), 
            .Q(mix_sinewave[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam sinewave_out_i6.GSR = "ENABLED";
    FD1S3AX sinewave_out_i7 (.D(sinewave_out_11__N_212[7]), .CK(clk_80mhz), 
            .Q(mix_sinewave[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam sinewave_out_i7.GSR = "ENABLED";
    FD1S3AX sinewave_out_i8 (.D(sinewave_out_11__N_212[8]), .CK(clk_80mhz), 
            .Q(mix_sinewave[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam sinewave_out_i8.GSR = "ENABLED";
    FD1S3AX sinewave_out_i9 (.D(sinewave_out_11__N_212[9]), .CK(clk_80mhz), 
            .Q(mix_sinewave[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam sinewave_out_i9.GSR = "ENABLED";
    FD1S3AX sinewave_out_i10 (.D(sinewave_out_11__N_212[10]), .CK(clk_80mhz), 
            .Q(mix_sinewave[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam sinewave_out_i10.GSR = "ENABLED";
    FD1S3AX sinewave_out_i11 (.D(sinewave_out_11__N_212[11]), .CK(clk_80mhz), 
            .Q(mix_sinewave[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam sinewave_out_i11.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i1 (.D(cosinewave_out_11__N_224[1]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam cosinewave_out_i1.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i2 (.D(cosinewave_out_11__N_224[2]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam cosinewave_out_i2.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i3 (.D(cosinewave_out_11__N_224[3]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam cosinewave_out_i3.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i4 (.D(cosinewave_out_11__N_224[4]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam cosinewave_out_i4.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i5 (.D(cosinewave_out_11__N_224[5]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam cosinewave_out_i5.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i6 (.D(cosinewave_out_11__N_224[6]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam cosinewave_out_i6.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i7 (.D(cosinewave_out_11__N_224[7]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam cosinewave_out_i7.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i8 (.D(cosinewave_out_11__N_224[8]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam cosinewave_out_i8.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i9 (.D(cosinewave_out_11__N_224[9]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam cosinewave_out_i9.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i10 (.D(cosinewave_out_11__N_224[10]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam cosinewave_out_i10.GSR = "ENABLED";
    FD1S3AX cosinewave_out_i11 (.D(cosinewave_out_11__N_224[11]), .CK(clk_80mhz), 
            .Q(mix_cosinewave[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=137, LSE_RLINE=145 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(43[10] 51[6])
    defparam cosinewave_out_i11.GSR = "ENABLED";
    LUT4 cosinewave_out_11__I_0_i11_3_lut (.A(\lo_cosinewave[11] ), .B(cosinewave_out_11__N_250[10]), 
         .C(rf_in_delayed_2), .Z(cosinewave_out_11__N_224[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam cosinewave_out_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 sinewave_out_11__I_0_i5_3_lut (.A(\lo_sinewave[5] ), .B(sinewave_out_11__N_236[4]), 
         .C(rf_in_delayed_2), .Z(sinewave_out_11__N_212[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam sinewave_out_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 sinewave_out_11__I_0_i6_3_lut (.A(\lo_sinewave[6] ), .B(sinewave_out_11__N_236[5]), 
         .C(rf_in_delayed_2), .Z(sinewave_out_11__N_212[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam sinewave_out_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 cosinewave_out_11__I_0_i1_3_lut (.A(\lo_cosinewave[1] ), .B(cosinewave_out_11__N_250[0]), 
         .C(rf_in_delayed_2), .Z(cosinewave_out_11__N_224[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam cosinewave_out_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 sinewave_out_11__I_0_i7_3_lut (.A(\lo_sinewave[7] ), .B(sinewave_out_11__N_236[6]), 
         .C(rf_in_delayed_2), .Z(sinewave_out_11__N_212[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam sinewave_out_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 sinewave_out_11__I_0_i8_3_lut (.A(\lo_sinewave[8] ), .B(sinewave_out_11__N_236[7]), 
         .C(rf_in_delayed_2), .Z(sinewave_out_11__N_212[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam sinewave_out_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 sinewave_out_11__I_0_i9_3_lut (.A(\lo_sinewave[9] ), .B(sinewave_out_11__N_236[8]), 
         .C(rf_in_delayed_2), .Z(sinewave_out_11__N_212[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam sinewave_out_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 sinewave_out_11__I_0_i10_3_lut (.A(\lo_sinewave[10] ), .B(sinewave_out_11__N_236[9]), 
         .C(rf_in_delayed_2), .Z(sinewave_out_11__N_212[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam sinewave_out_11__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 sinewave_out_11__I_0_i11_3_lut (.A(\lo_sinewave[11] ), .B(sinewave_out_11__N_236[10]), 
         .C(rf_in_delayed_2), .Z(sinewave_out_11__N_212[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam sinewave_out_11__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 sinewave_out_11__I_0_i12_3_lut (.A(\lo_sinewave[12] ), .B(sinewave_out_11__N_236[11]), 
         .C(rf_in_delayed_2), .Z(sinewave_out_11__N_212[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam sinewave_out_11__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 cosinewave_out_11__I_0_i2_3_lut (.A(\lo_cosinewave[2] ), .B(cosinewave_out_11__N_250[1]), 
         .C(rf_in_delayed_2), .Z(cosinewave_out_11__N_224[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam cosinewave_out_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 cosinewave_out_11__I_0_i3_3_lut (.A(\lo_cosinewave[3] ), .B(cosinewave_out_11__N_250[2]), 
         .C(rf_in_delayed_2), .Z(cosinewave_out_11__N_224[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam cosinewave_out_11__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 cosinewave_out_11__I_0_i4_3_lut (.A(\lo_cosinewave[4] ), .B(cosinewave_out_11__N_250[3]), 
         .C(rf_in_delayed_2), .Z(cosinewave_out_11__N_224[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam cosinewave_out_11__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 cosinewave_out_11__I_0_i5_3_lut (.A(\lo_cosinewave[5] ), .B(cosinewave_out_11__N_250[4]), 
         .C(rf_in_delayed_2), .Z(cosinewave_out_11__N_224[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam cosinewave_out_11__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 cosinewave_out_11__I_0_i6_3_lut (.A(\lo_cosinewave[6] ), .B(cosinewave_out_11__N_250[5]), 
         .C(rf_in_delayed_2), .Z(cosinewave_out_11__N_224[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam cosinewave_out_11__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 cosinewave_out_11__I_0_i12_3_lut (.A(\lo_cosinewave[12] ), .B(cosinewave_out_11__N_250[11]), 
         .C(rf_in_delayed_2), .Z(cosinewave_out_11__N_224[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam cosinewave_out_11__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 cosinewave_out_11__I_0_i7_3_lut (.A(\lo_cosinewave[7] ), .B(cosinewave_out_11__N_250[6]), 
         .C(rf_in_delayed_2), .Z(cosinewave_out_11__N_224[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam cosinewave_out_11__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 cosinewave_out_11__I_0_i8_3_lut (.A(\lo_cosinewave[8] ), .B(cosinewave_out_11__N_250[7]), 
         .C(rf_in_delayed_2), .Z(cosinewave_out_11__N_224[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam cosinewave_out_11__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 sinewave_out_11__I_0_i2_3_lut (.A(\lo_sinewave[2] ), .B(sinewave_out_11__N_236[1]), 
         .C(rf_in_delayed_2), .Z(sinewave_out_11__N_212[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam sinewave_out_11__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 sinewave_out_11__I_0_i1_3_lut (.A(\lo_sinewave[1] ), .B(sinewave_out_11__N_236[0]), 
         .C(rf_in_delayed_2), .Z(sinewave_out_11__N_212[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam sinewave_out_11__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 cosinewave_out_11__I_0_i9_3_lut (.A(\lo_cosinewave[9] ), .B(cosinewave_out_11__N_250[8]), 
         .C(rf_in_delayed_2), .Z(cosinewave_out_11__N_224[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam cosinewave_out_11__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 sinewave_out_11__I_0_i3_3_lut (.A(\lo_sinewave[3] ), .B(sinewave_out_11__N_236[2]), 
         .C(rf_in_delayed_2), .Z(sinewave_out_11__N_212[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/Mixer.v(47[14] 50[8])
    defparam sinewave_out_11__I_0_i3_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module \CIC(REGISTER_WIDTH=72,DECIMATION_RATIO=4096) 
//

module \CIC(REGISTER_WIDTH=72,DECIMATION_RATIO=4096)  (integrator_d_tmp, clk_80mhz, 
            integrator_tmp, n30, integrator5, integrator2, integrator2_71__N_490, 
            n33, integrator3, integrator3_71__N_562, integrator4, integrator4_71__N_634, 
            integrator5_71__N_706, comb6, comb6_71__N_1451, cic_sine_clk, 
            comb_d6, comb7, comb7_71__N_1523, comb_d7, comb8, comb8_71__N_1595, 
            comb_d8, comb9, comb9_71__N_1667, comb_d9, mult_i_b, integrator1, 
            integrator1_71__N_418, count, n32, n35, n34, n37, n36, 
            n67, \cic_gain[0] , \comb10[66] , \comb10[67] , \comb10[69] , 
            \comb10[68] , \comb10[65] , \cic_gain[1] , \comb10[70] , 
            \comb10[71] , n63, \data_out_11__N_1811[2] , n64, \data_out_11__N_1811[3] , 
            n65, \data_out_11__N_1811[4] , n66, \data_out_11__N_1811[5] , 
            \data_out_11__N_1811[6] , \data_out_11__N_1811[7] , n118, 
            n120, cout, n115, n117, n112, n114, n109, n111, 
            n106, n108, n103, n105, n100, n102, \comb10[64] , 
            \comb10[62] , \comb10[63] , n97, n99, \comb10[61] , n94, 
            n96, n91, n93, n16607, \comb10[59] , n62, \comb10[60] , 
            n88, n90, n85, n87, n82, n84, n79, n81, n76, n78, 
            n3, n2, n5, n4, n7, n6, n9, n8, n11, n10, n13, 
            n12, n15, n14, n17, n16, n19, n18, n21, n20, n23, 
            n22, n25, n24, n27, n26, n29, n28_adj_115, n31_adj_116, 
            n30_adj_117, n33_adj_118, n32_adj_119, n35_adj_120, n34_adj_121, 
            n37_adj_122, n36_adj_123, n3_adj_124, n2_adj_125, n5_adj_126, 
            n4_adj_127, n3_adj_128, n2_adj_129, n5_adj_130, n4_adj_131, 
            n7_adj_132, n6_adj_133, n9_adj_134, n8_adj_135, n11_adj_136, 
            n10_adj_137, n13_adj_138, n12_adj_139, n15_adj_140, n14_adj_141, 
            n17_adj_142, n16_adj_143, n19_adj_144, n18_adj_145, n21_adj_146, 
            n20_adj_147, n7_adj_148, n6_adj_149, n9_adj_150, n8_adj_151, 
            n11_adj_152, n10_adj_153, n13_adj_154, n12_adj_155, n15_adj_156, 
            n14_adj_157, n17_adj_158, n16_adj_159, n19_adj_160, \data_out_11__N_1811[10] , 
            n18_adj_161, n21_adj_162, n20_adj_163, n23_adj_164, n22_adj_165, 
            n23_adj_166, n22_adj_167, n25_adj_168, n24_adj_169, n27_adj_170, 
            \data_out_11__N_1811[11] , n26_adj_171, n29_adj_172, n28_adj_173, 
            n31_adj_174, n30_adj_175, n25_adj_176, n24_adj_177, n33_adj_178, 
            n32_adj_179, n35_adj_180, n34_adj_181, n37_adj_182, n36_adj_183, 
            n27_adj_184, n26_adj_185, n29_adj_186, n28_adj_187, n31_adj_188, 
            n30_adj_189, n33_adj_190, n32_adj_191, n35_adj_192, n34_adj_193, 
            n37_adj_194, n36_adj_195, \data_out_11__N_1811[8] , n3_adj_196, 
            n2_adj_197, n5_adj_198, n4_adj_199, n7_adj_200, \data_out_11__N_1811[9] , 
            n6_adj_201, n9_adj_202, n8_adj_203, n11_adj_204, n10_adj_205, 
            n13_adj_206, n12_adj_207, n15_adj_208, n14_adj_209, n17_adj_210, 
            n16_adj_211, n19_adj_212, n18_adj_213, n21_adj_214, n20_adj_215, 
            n23_adj_216, n22_adj_217, n25_adj_218, n24_adj_219, n27_adj_220, 
            n26_adj_221, n29_adj_222, n28_adj_223, n31_adj_224) /* synthesis syn_module_defined=1 */ ;
    output [71:0]integrator_d_tmp;
    input clk_80mhz;
    output [71:0]integrator_tmp;
    output n30;
    output [71:0]integrator5;
    output [71:0]integrator2;
    input [71:0]integrator2_71__N_490;
    output n33;
    output [71:0]integrator3;
    input [71:0]integrator3_71__N_562;
    output [71:0]integrator4;
    input [71:0]integrator4_71__N_634;
    input [71:0]integrator5_71__N_706;
    output [71:0]comb6;
    input [71:0]comb6_71__N_1451;
    output cic_sine_clk;
    output [71:0]comb_d6;
    output [71:0]comb7;
    input [71:0]comb7_71__N_1523;
    output [71:0]comb_d7;
    output [71:0]comb8;
    input [71:0]comb8_71__N_1595;
    output [71:0]comb_d8;
    output [71:0]comb9;
    input [71:0]comb9_71__N_1667;
    output [71:0]comb_d9;
    output [11:0]mult_i_b;
    output [71:0]integrator1;
    input [71:0]integrator1_71__N_418;
    output [11:0]count;
    output n32;
    output n35;
    output n34;
    output n37;
    output n36;
    input [11:0]n67;
    input \cic_gain[0] ;
    input \comb10[66] ;
    input \comb10[67] ;
    input \comb10[69] ;
    input \comb10[68] ;
    input \comb10[65] ;
    input \cic_gain[1] ;
    input \comb10[70] ;
    input \comb10[71] ;
    input n63;
    output \data_out_11__N_1811[2] ;
    input n64;
    output \data_out_11__N_1811[3] ;
    input n65;
    output \data_out_11__N_1811[4] ;
    input n66;
    output \data_out_11__N_1811[5] ;
    output \data_out_11__N_1811[6] ;
    output \data_out_11__N_1811[7] ;
    input n118;
    input n120;
    input cout;
    input n115;
    input n117;
    input n112;
    input n114;
    input n109;
    input n111;
    input n106;
    input n108;
    input n103;
    input n105;
    input n100;
    input n102;
    input \comb10[64] ;
    input \comb10[62] ;
    input \comb10[63] ;
    input n97;
    input n99;
    input \comb10[61] ;
    input n94;
    input n96;
    input n91;
    input n93;
    input n16607;
    input \comb10[59] ;
    input n62;
    input \comb10[60] ;
    input n88;
    input n90;
    input n85;
    input n87;
    input n82;
    input n84;
    input n79;
    input n81;
    input n76;
    input n78;
    output n3;
    output n2;
    output n5;
    output n4;
    output n7;
    output n6;
    output n9;
    output n8;
    output n11;
    output n10;
    output n13;
    output n12;
    output n15;
    output n14;
    output n17;
    output n16;
    output n19;
    output n18;
    output n21;
    output n20;
    output n23;
    output n22;
    output n25;
    output n24;
    output n27;
    output n26;
    output n29;
    output n28_adj_115;
    output n31_adj_116;
    output n30_adj_117;
    output n33_adj_118;
    output n32_adj_119;
    output n35_adj_120;
    output n34_adj_121;
    output n37_adj_122;
    output n36_adj_123;
    output n3_adj_124;
    output n2_adj_125;
    output n5_adj_126;
    output n4_adj_127;
    output n3_adj_128;
    output n2_adj_129;
    output n5_adj_130;
    output n4_adj_131;
    output n7_adj_132;
    output n6_adj_133;
    output n9_adj_134;
    output n8_adj_135;
    output n11_adj_136;
    output n10_adj_137;
    output n13_adj_138;
    output n12_adj_139;
    output n15_adj_140;
    output n14_adj_141;
    output n17_adj_142;
    output n16_adj_143;
    output n19_adj_144;
    output n18_adj_145;
    output n21_adj_146;
    output n20_adj_147;
    output n7_adj_148;
    output n6_adj_149;
    output n9_adj_150;
    output n8_adj_151;
    output n11_adj_152;
    output n10_adj_153;
    output n13_adj_154;
    output n12_adj_155;
    output n15_adj_156;
    output n14_adj_157;
    output n17_adj_158;
    output n16_adj_159;
    output n19_adj_160;
    output \data_out_11__N_1811[10] ;
    output n18_adj_161;
    output n21_adj_162;
    output n20_adj_163;
    output n23_adj_164;
    output n22_adj_165;
    output n23_adj_166;
    output n22_adj_167;
    output n25_adj_168;
    output n24_adj_169;
    output n27_adj_170;
    output \data_out_11__N_1811[11] ;
    output n26_adj_171;
    output n29_adj_172;
    output n28_adj_173;
    output n31_adj_174;
    output n30_adj_175;
    output n25_adj_176;
    output n24_adj_177;
    output n33_adj_178;
    output n32_adj_179;
    output n35_adj_180;
    output n34_adj_181;
    output n37_adj_182;
    output n36_adj_183;
    output n27_adj_184;
    output n26_adj_185;
    output n29_adj_186;
    output n28_adj_187;
    output n31_adj_188;
    output n30_adj_189;
    output n33_adj_190;
    output n32_adj_191;
    output n35_adj_192;
    output n34_adj_193;
    output n37_adj_194;
    output n36_adj_195;
    output \data_out_11__N_1811[8] ;
    output n3_adj_196;
    output n2_adj_197;
    output n5_adj_198;
    output n4_adj_199;
    output n7_adj_200;
    output \data_out_11__N_1811[9] ;
    output n6_adj_201;
    output n9_adj_202;
    output n8_adj_203;
    output n11_adj_204;
    output n10_adj_205;
    output n13_adj_206;
    output n12_adj_207;
    output n15_adj_208;
    output n14_adj_209;
    output n17_adj_210;
    output n16_adj_211;
    output n19_adj_212;
    output n18_adj_213;
    output n21_adj_214;
    output n20_adj_215;
    output n23_adj_216;
    output n22_adj_217;
    output n25_adj_218;
    output n24_adj_219;
    output n27_adj_220;
    output n26_adj_221;
    output n29_adj_222;
    output n28_adj_223;
    output n31_adj_224;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(64[10:19])
    wire cic_sine_clk /* synthesis SET_AS_NETWORK=cic_sine_clk, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(86[10:22])
    
    wire clk_80mhz_enable_1508, clk_80mhz_enable_99, decimation_clk, n11887, 
        valid_comb, clk_80mhz_enable_38;
    wire [71:0]data_out_11__N_1811;
    wire [11:0]count_11__N_1438;
    
    wire clk_80mhz_enable_186, clk_80mhz_enable_149, n11935, n17180, 
        n17179, n17183, n17182;
    wire [71:0]comb10;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[105:111])
    
    wire n17186, n17185, n17189, n17188, n17192, n17191, n16626, 
        n17195, n17194, n17198, n17197, n17201, n17200, n17204, 
        n16640, n17203, n17207, n16650, n17206, n63_c, n131, n64_c, 
        n132, n65_c, n133, n66_c, n134, n135, n136, n131_adj_2589, 
        n132_adj_2592, n133_adj_2595, n134_adj_2598, n135_adj_2600, 
        n136_adj_2602;
    wire [71:0]comb10_71__N_1739;
    
    wire clk_80mhz_enable_744, clk_80mhz_enable_236, clk_80mhz_enable_286, 
        clk_80mhz_enable_336, clk_80mhz_enable_386, clk_80mhz_enable_436, 
        clk_80mhz_enable_486, clk_80mhz_enable_536, clk_80mhz_enable_586, 
        clk_80mhz_enable_636, clk_80mhz_enable_686, clk_80mhz_enable_736, 
        clk_80mhz_enable_737, clk_80mhz_enable_738, clk_80mhz_enable_739, 
        clk_80mhz_enable_740, clk_80mhz_enable_741, clk_80mhz_enable_742, 
        clk_80mhz_enable_743, clk_80mhz_enable_745, clk_80mhz_enable_746, 
        clk_80mhz_enable_747, decimation_clk_N_1823, n73, n16525, n16509, 
        n16517, n16521, n16569, n16553, n17316, n16565, n16551;
    
    FD1P3AX integrator_d_tmp_i0_i55 (.D(integrator_tmp[55]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i54 (.D(integrator_tmp[54]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i53 (.D(integrator_tmp[53]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i52 (.D(integrator_tmp[52]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i51 (.D(integrator_tmp[51]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i50 (.D(integrator_tmp[50]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i49 (.D(integrator_tmp[49]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i48 (.D(integrator_tmp[48]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i47 (.D(integrator_tmp[47]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i46 (.D(integrator_tmp[46]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i46.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i44_1_lut (.A(integrator_d_tmp[43]), .Z(n30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i44_1_lut.init = 16'h5555;
    FD1P3AX integrator_d_tmp_i0_i45 (.D(integrator_tmp[45]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i0 (.D(integrator5[0]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i0 (.D(integrator_tmp[0]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i44 (.D(integrator_tmp[44]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i43 (.D(integrator_tmp[43]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i42 (.D(integrator_tmp[42]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i41 (.D(integrator_tmp[41]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i40 (.D(integrator_tmp[40]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i39 (.D(integrator_tmp[39]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i38 (.D(integrator_tmp[38]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i37 (.D(integrator_tmp[37]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i36 (.D(integrator_tmp[36]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i36.GSR = "ENABLED";
    FD1S3AX integrator2_i0 (.D(integrator2_71__N_490[0]), .CK(clk_80mhz), 
            .Q(integrator2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i0.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i41_1_lut (.A(integrator_d_tmp[40]), .Z(n33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i41_1_lut.init = 16'h5555;
    FD1P3AX integrator_d_tmp_i0_i35 (.D(integrator_tmp[35]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i34 (.D(integrator_tmp[34]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i34.GSR = "ENABLED";
    FD1S3AX integrator3_i0 (.D(integrator3_71__N_562[0]), .CK(clk_80mhz), 
            .Q(integrator3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i0.GSR = "ENABLED";
    FD1S3AX integrator4_i0 (.D(integrator4_71__N_634[0]), .CK(clk_80mhz), 
            .Q(integrator4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i0.GSR = "ENABLED";
    FD1S3AX integrator5_i0 (.D(integrator5_71__N_706[0]), .CK(clk_80mhz), 
            .Q(integrator5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i0.GSR = "ENABLED";
    FD1P3AX comb6_i0_i0 (.D(comb6_71__N_1451[0]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(comb6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i0.GSR = "ENABLED";
    FD1S3JX decimation_clk_65 (.D(n11887), .CK(clk_80mhz), .PD(clk_80mhz_enable_99), 
            .Q(decimation_clk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam decimation_clk_65.GSR = "ENABLED";
    FD1S3AX valid_comb_66 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), .Q(valid_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66.GSR = "ENABLED";
    FD1S3AX data_clk_67 (.D(decimation_clk), .CK(clk_80mhz), .Q(cic_sine_clk)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_clk_67.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i33 (.D(integrator_tmp[33]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i32 (.D(integrator_tmp[32]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i31 (.D(integrator_tmp[31]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i30 (.D(integrator_tmp[30]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i0 (.D(comb6[0]), .SP(clk_80mhz_enable_1508), .CK(clk_80mhz), 
            .Q(comb_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i0.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i29 (.D(integrator_tmp[29]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX comb7_i0_i0 (.D(comb7_71__N_1523[0]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(comb7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i0 (.D(comb7[0]), .SP(clk_80mhz_enable_1508), .CK(clk_80mhz), 
            .Q(comb_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX comb8_i0_i0 (.D(comb8_71__N_1595[0]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(comb8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i0 (.D(comb8[0]), .SP(clk_80mhz_enable_1508), .CK(clk_80mhz), 
            .Q(comb_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX comb9_i0_i0 (.D(comb9_71__N_1667[0]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(comb9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i0 (.D(comb9[0]), .SP(clk_80mhz_enable_1508), .CK(clk_80mhz), 
            .Q(comb_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i0.GSR = "ENABLED";
    FD1P3AX data_out_i0_i0 (.D(data_out_11__N_1811[0]), .SP(clk_80mhz_enable_38), 
            .CK(clk_80mhz), .Q(mult_i_b[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i0.GSR = "ENABLED";
    FD1S3AX integrator1_i0 (.D(integrator1_71__N_418[0]), .CK(clk_80mhz), 
            .Q(integrator1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i0.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i28 (.D(integrator_tmp[28]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i27 (.D(integrator_tmp[27]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i26 (.D(integrator_tmp[26]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i25 (.D(integrator_tmp[25]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i25.GSR = "ENABLED";
    FD1S3IX count__i0 (.D(count_11__N_1438[0]), .CK(clk_80mhz), .CD(clk_80mhz_enable_99), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i0.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i24 (.D(integrator_tmp[24]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i23 (.D(integrator_tmp[23]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i22 (.D(integrator_tmp[22]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i21 (.D(integrator_tmp[21]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i20 (.D(integrator_tmp[20]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i19 (.D(integrator_tmp[19]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i18 (.D(integrator_tmp[18]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i17 (.D(integrator_tmp[17]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i16 (.D(integrator_tmp[16]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i15 (.D(integrator_tmp[15]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i14 (.D(integrator_tmp[14]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i13 (.D(integrator_tmp[13]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i12 (.D(integrator_tmp[12]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i11 (.D(integrator_tmp[11]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i10 (.D(integrator_tmp[10]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i9 (.D(integrator_tmp[9]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i8 (.D(integrator_tmp[8]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i7 (.D(integrator_tmp[7]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i6 (.D(integrator_tmp[6]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i5 (.D(integrator_tmp[5]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i4 (.D(integrator_tmp[4]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i4.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i42_1_lut (.A(integrator_d_tmp[41]), .Z(n32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i42_1_lut.init = 16'h5555;
    FD1P3AX integrator_d_tmp_i0_i3 (.D(integrator_tmp[3]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i3.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i39_1_lut (.A(integrator_d_tmp[38]), .Z(n35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i39_1_lut.init = 16'h5555;
    FD1P3AX integrator_d_tmp_i0_i2 (.D(integrator_tmp[2]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i2.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i40_1_lut (.A(integrator_d_tmp[39]), .Z(n34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i40_1_lut.init = 16'h5555;
    FD1P3AX integrator_d_tmp_i0_i1 (.D(integrator_tmp[1]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i71 (.D(integrator5[71]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i70 (.D(integrator5[70]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i69 (.D(integrator5[69]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i68 (.D(integrator5[68]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i67 (.D(integrator5[67]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i66 (.D(integrator5[66]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i65 (.D(integrator5[65]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i64 (.D(integrator5[64]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i63 (.D(integrator5[63]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i62 (.D(integrator5[62]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i61 (.D(integrator5[61]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i60 (.D(integrator5[60]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i60.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i37_1_lut (.A(integrator_d_tmp[36]), .Z(n37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i38_1_lut (.A(integrator_d_tmp[37]), .Z(n36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i38_1_lut.init = 16'h5555;
    FD1P3AX integrator_tmp_i0_i59 (.D(integrator5[59]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i58 (.D(integrator5[58]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i57 (.D(integrator5[57]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i56 (.D(integrator5[56]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i55 (.D(integrator5[55]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i54 (.D(integrator5[54]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i53 (.D(integrator5[53]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i52 (.D(integrator5[52]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i51 (.D(integrator5[51]), .SP(clk_80mhz_enable_99), 
            .CK(clk_80mhz), .Q(integrator_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i50 (.D(integrator5[50]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i49 (.D(integrator5[49]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i48 (.D(integrator5[48]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i47 (.D(integrator5[47]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i46 (.D(integrator5[46]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i45 (.D(integrator5[45]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i44 (.D(integrator5[44]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i43 (.D(integrator5[43]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i42 (.D(integrator5[42]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i41 (.D(integrator5[41]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i40 (.D(integrator5[40]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i39 (.D(integrator5[39]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i38 (.D(integrator5[38]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i37 (.D(integrator5[37]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i36 (.D(integrator5[36]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i35 (.D(integrator5[35]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i34 (.D(integrator5[34]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i33 (.D(integrator5[33]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i32 (.D(integrator5[32]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i31 (.D(integrator5[31]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i30 (.D(integrator5[30]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i29 (.D(integrator5[29]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i28 (.D(integrator5[28]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i27 (.D(integrator5[27]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i26 (.D(integrator5[26]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i25 (.D(integrator5[25]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i24 (.D(integrator5[24]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i23 (.D(integrator5[23]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i22 (.D(integrator5[22]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i21 (.D(integrator5[21]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i20 (.D(integrator5[20]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i19 (.D(integrator5[19]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i18 (.D(integrator5[18]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i17 (.D(integrator5[17]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i16 (.D(integrator5[16]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i15 (.D(integrator5[15]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i14 (.D(integrator5[14]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i13 (.D(integrator5[13]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i12 (.D(integrator5[12]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i11 (.D(integrator5[11]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i10 (.D(integrator5[10]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i9 (.D(integrator5[9]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i8 (.D(integrator5[8]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i7 (.D(integrator5[7]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i6 (.D(integrator5[6]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i5 (.D(integrator5[5]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i4 (.D(integrator5[4]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i3 (.D(integrator5[3]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i2 (.D(integrator5[2]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i1 (.D(integrator5[1]), .SP(clk_80mhz_enable_149), 
            .CK(clk_80mhz), .Q(integrator_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i1.GSR = "ENABLED";
    FD1S3IX count__i1 (.D(n67[1]), .CK(clk_80mhz), .CD(n11935), .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i1.GSR = "ENABLED";
    LUT4 shift_right_31_i210_3_lut_4_lut_then_3_lut (.A(\cic_gain[0] ), .B(\comb10[66] ), 
         .C(\comb10[67] ), .Z(n17180)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 shift_right_31_i210_3_lut_4_lut_else_3_lut (.A(\cic_gain[0] ), .B(\comb10[69] ), 
         .C(\comb10[68] ), .Z(n17179)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam shift_right_31_i210_3_lut_4_lut_else_3_lut.init = 16'he4e4;
    LUT4 shift_right_31_i209_3_lut_4_lut_then_3_lut (.A(\cic_gain[0] ), .B(\comb10[65] ), 
         .C(\comb10[66] ), .Z(n17183)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam shift_right_31_i209_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 shift_right_31_i209_3_lut_4_lut_else_3_lut (.A(\cic_gain[0] ), .B(\comb10[68] ), 
         .C(\comb10[67] ), .Z(n17182)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam shift_right_31_i209_3_lut_4_lut_else_3_lut.init = 16'he4e4;
    LUT4 shift_right_31_i209_3_lut_4_lut_then_3_lut_adj_161 (.A(\cic_gain[0] ), 
         .B(comb10[65]), .C(comb10[66]), .Z(n17186)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam shift_right_31_i209_3_lut_4_lut_then_3_lut_adj_161.init = 16'hd8d8;
    LUT4 shift_right_31_i209_3_lut_4_lut_else_3_lut_adj_162 (.A(\cic_gain[0] ), 
         .B(comb10[68]), .C(comb10[67]), .Z(n17185)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam shift_right_31_i209_3_lut_4_lut_else_3_lut_adj_162.init = 16'he4e4;
    LUT4 shift_right_31_i212_3_lut_4_lut_then_3_lut (.A(\cic_gain[1] ), .B(\comb10[68] ), 
         .C(\comb10[70] ), .Z(n17189)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i212_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 shift_right_31_i212_3_lut_4_lut_else_3_lut (.A(\comb10[71] ), .B(\cic_gain[1] ), 
         .C(\comb10[69] ), .Z(n17188)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i212_3_lut_4_lut_else_3_lut.init = 16'he2e2;
    LUT4 i11_3_lut_4_lut_then_3_lut (.A(\cic_gain[1] ), .B(\comb10[67] ), 
         .C(\comb10[69] ), .Z(n17192)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam i11_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 i11_3_lut_4_lut_else_3_lut (.A(\comb10[70] ), .B(\cic_gain[1] ), 
         .C(\comb10[68] ), .Z(n17191)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam i11_3_lut_4_lut_else_3_lut.init = 16'he2e2;
    LUT4 shift_right_31_i212_3_lut_4_lut_then_4_lut (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(comb10[68]), .D(n16626), .Z(n17195)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((D)+!B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i212_3_lut_4_lut_then_4_lut.init = 16'hf791;
    LUT4 shift_right_31_i212_3_lut_4_lut_else_4_lut (.A(\cic_gain[0] ), .B(\cic_gain[1] ), 
         .C(comb10[68]), .D(n16626), .Z(n17194)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (D))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i212_3_lut_4_lut_else_4_lut.init = 16'he680;
    LUT4 i11_3_lut_4_lut_then_3_lut_adj_163 (.A(\cic_gain[1] ), .B(comb10[67]), 
         .C(comb10[69]), .Z(n17198)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam i11_3_lut_4_lut_then_3_lut_adj_163.init = 16'hd8d8;
    LUT4 i11_3_lut_4_lut_else_3_lut_adj_164 (.A(comb10[70]), .B(\cic_gain[1] ), 
         .C(comb10[68]), .Z(n17197)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam i11_3_lut_4_lut_else_3_lut_adj_164.init = 16'he2e2;
    LUT4 i5806_then_3_lut (.A(\cic_gain[1] ), .B(comb10[68]), .C(comb10[66]), 
         .Z(n17201)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5806_then_3_lut.init = 16'he4e4;
    LUT4 i5806_else_3_lut (.A(n16626), .B(\cic_gain[1] ), .C(comb10[67]), 
         .Z(n17200)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5806_else_3_lut.init = 16'he2e2;
    LUT4 i5809_then_3_lut (.A(\cic_gain[1] ), .B(comb10[60]), .C(comb10[58]), 
         .Z(n17204)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5809_then_3_lut.init = 16'he4e4;
    LUT4 i5809_else_3_lut (.A(n16640), .B(\cic_gain[1] ), .C(comb10[59]), 
         .Z(n17203)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5809_else_3_lut.init = 16'he2e2;
    LUT4 i5799_then_3_lut (.A(\cic_gain[1] ), .B(comb10[59]), .C(comb10[57]), 
         .Z(n17207)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5799_then_3_lut.init = 16'he4e4;
    LUT4 i5799_else_3_lut (.A(n16650), .B(\cic_gain[1] ), .C(comb10[58]), 
         .Z(n17206)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5799_else_3_lut.init = 16'he2e2;
    LUT4 shift_right_31_i203_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n63_c), .D(n131), .Z(data_out_11__N_1811[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i204_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n64_c), .D(n132), .Z(data_out_11__N_1811[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i205_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n65_c), .D(n133), .Z(data_out_11__N_1811[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i206_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n66_c), .D(n134), .Z(data_out_11__N_1811[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i207_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(comb10[66]), .D(n135), .Z(data_out_11__N_1811[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i208_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(comb10[67]), .D(n136), .Z(data_out_11__N_1811[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut.init = 16'hfe10;
    LUT4 shift_right_31_i203_3_lut_4_lut_adj_165 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n63), .D(n131_adj_2589), .Z(\data_out_11__N_1811[2] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i203_3_lut_4_lut_adj_165.init = 16'hfe10;
    LUT4 shift_right_31_i204_3_lut_4_lut_adj_166 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n64), .D(n132_adj_2592), .Z(\data_out_11__N_1811[3] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i204_3_lut_4_lut_adj_166.init = 16'hfe10;
    LUT4 shift_right_31_i205_3_lut_4_lut_adj_167 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n65), .D(n133_adj_2595), .Z(\data_out_11__N_1811[4] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i205_3_lut_4_lut_adj_167.init = 16'hfe10;
    LUT4 shift_right_31_i206_3_lut_4_lut_adj_168 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n66), .D(n134_adj_2598), .Z(\data_out_11__N_1811[5] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i206_3_lut_4_lut_adj_168.init = 16'hfe10;
    LUT4 shift_right_31_i207_3_lut_4_lut_adj_169 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(\comb10[66] ), .D(n135_adj_2600), .Z(\data_out_11__N_1811[6] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i207_3_lut_4_lut_adj_169.init = 16'hfe10;
    LUT4 shift_right_31_i208_3_lut_4_lut_adj_170 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(\comb10[67] ), .D(n136_adj_2602), .Z(\data_out_11__N_1811[7] )) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam shift_right_31_i208_3_lut_4_lut_adj_170.init = 16'hfe10;
    LUT4 mux_873_i2_3_lut (.A(n118), .B(n120), .C(cout), .Z(comb10_71__N_1739[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i2_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i135_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n65_c), .D(comb10[63]), .Z(n135)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i134_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n64_c), .D(comb10[62]), .Z(n134)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut.init = 16'hf960;
    LUT4 mux_873_i3_3_lut (.A(n115), .B(n117), .C(cout), .Z(comb10_71__N_1739[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i3_3_lut.init = 16'hcaca;
    LUT4 mux_873_i4_3_lut (.A(n112), .B(n114), .C(cout), .Z(comb10_71__N_1739[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i4_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i133_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n63_c), .D(comb10[61]), .Z(n133)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i132_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n16640), .D(comb10[60]), .Z(n132)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut.init = 16'hf960;
    LUT4 mux_873_i5_3_lut (.A(n109), .B(n111), .C(cout), .Z(comb10_71__N_1739[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i5_3_lut.init = 16'hcaca;
    LUT4 mux_873_i6_3_lut (.A(n106), .B(n108), .C(cout), .Z(comb10_71__N_1739[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i6_3_lut.init = 16'hcaca;
    FD1S3AX valid_comb_66_rep_381 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_744)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_381.GSR = "ENABLED";
    LUT4 mux_873_i7_3_lut (.A(n103), .B(n105), .C(cout), .Z(comb10_71__N_1739[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i7_3_lut.init = 16'hcaca;
    LUT4 mux_873_i8_3_lut (.A(n100), .B(n102), .C(cout), .Z(comb10_71__N_1739[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i8_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i136_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n66), .D(\comb10[64] ), .Z(n136_adj_2602)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i134_3_lut_4_lut_adj_171 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n64), .D(\comb10[62] ), .Z(n134_adj_2598)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i134_3_lut_4_lut_adj_171.init = 16'hf960;
    LUT4 shift_right_31_i135_3_lut_4_lut_adj_172 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n65), .D(\comb10[63] ), .Z(n135_adj_2600)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i135_3_lut_4_lut_adj_172.init = 16'hf960;
    LUT4 mux_873_i9_3_lut (.A(n97), .B(n99), .C(cout), .Z(comb10_71__N_1739[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i9_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i133_3_lut_4_lut_adj_173 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n63), .D(\comb10[61] ), .Z(n133_adj_2595)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i133_3_lut_4_lut_adj_173.init = 16'hf960;
    LUT4 mux_873_i10_3_lut (.A(n94), .B(n96), .C(cout), .Z(comb10_71__N_1739[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i10_3_lut.init = 16'hcaca;
    LUT4 mux_873_i11_3_lut (.A(n91), .B(n93), .C(cout), .Z(comb10_71__N_1739[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i11_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i131_3_lut_4_lut (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n16607), .D(\comb10[59] ), .Z(n131_adj_2589)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut.init = 16'hf960;
    LUT4 shift_right_31_i132_3_lut_4_lut_adj_174 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n62), .D(\comb10[60] ), .Z(n132_adj_2592)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i132_3_lut_4_lut_adj_174.init = 16'hf960;
    LUT4 mux_873_i12_3_lut (.A(n88), .B(n90), .C(cout), .Z(comb10_71__N_1739[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i12_3_lut.init = 16'hcaca;
    LUT4 mux_873_i13_3_lut (.A(n85), .B(n87), .C(cout), .Z(comb10_71__N_1739[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i13_3_lut.init = 16'hcaca;
    LUT4 mux_873_i14_3_lut (.A(n82), .B(n84), .C(cout), .Z(comb10_71__N_1739[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i14_3_lut.init = 16'hcaca;
    LUT4 mux_873_i15_3_lut (.A(n79), .B(n81), .C(cout), .Z(comb10_71__N_1739[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i15_3_lut.init = 16'hcaca;
    LUT4 mux_873_i16_3_lut (.A(n76), .B(n78), .C(cout), .Z(comb10_71__N_1739[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_873_i16_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i62_rep_218_3_lut (.A(comb10[61]), .B(comb10[62]), 
         .C(\cic_gain[0] ), .Z(n16640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i62_rep_218_3_lut.init = 16'hcaca;
    FD1P3AX integrator_d_tmp_i0_i57 (.D(integrator_tmp[57]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i57.GSR = "ENABLED";
    LUT4 shift_right_31_i63_3_lut (.A(comb10[62]), .B(comb10[63]), .C(\cic_gain[0] ), 
         .Z(n63_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    FD1P3AX integrator_d_tmp_i0_i58 (.D(integrator_tmp[58]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i59 (.D(integrator_tmp[59]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i60 (.D(integrator_tmp[60]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i61 (.D(integrator_tmp[61]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i62 (.D(integrator_tmp[62]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i63 (.D(integrator_tmp[63]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i64 (.D(integrator_tmp[64]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i65 (.D(integrator_tmp[65]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i66 (.D(integrator_tmp[66]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i67 (.D(integrator_tmp[67]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i68 (.D(integrator_tmp[68]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i69 (.D(integrator_tmp[69]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i70 (.D(integrator_tmp[70]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i71 (.D(integrator_tmp[71]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i71.GSR = "ENABLED";
    LUT4 shift_right_31_i64_3_lut (.A(comb10[63]), .B(comb10[64]), .C(\cic_gain[0] ), 
         .Z(n64_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i65_3_lut (.A(comb10[64]), .B(comb10[65]), .C(\cic_gain[0] ), 
         .Z(n65_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i131_3_lut_4_lut_adj_175 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n16650), .D(comb10[59]), .Z(n131)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i131_3_lut_4_lut_adj_175.init = 16'hf960;
    LUT4 shift_right_31_i66_3_lut (.A(comb10[65]), .B(comb10[66]), .C(\cic_gain[0] ), 
         .Z(n66_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i136_3_lut_4_lut_adj_176 (.A(\cic_gain[1] ), .B(\cic_gain[0] ), 
         .C(n66_c), .D(comb10[64]), .Z(n136)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam shift_right_31_i136_3_lut_4_lut_adj_176.init = 16'hf960;
    FD1S3AX integrator2_i1 (.D(integrator2_71__N_490[1]), .CK(clk_80mhz), 
            .Q(integrator2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i1.GSR = "ENABLED";
    FD1S3AX integrator2_i2 (.D(integrator2_71__N_490[2]), .CK(clk_80mhz), 
            .Q(integrator2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i2.GSR = "ENABLED";
    FD1S3AX integrator2_i3 (.D(integrator2_71__N_490[3]), .CK(clk_80mhz), 
            .Q(integrator2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i3.GSR = "ENABLED";
    FD1S3AX integrator2_i4 (.D(integrator2_71__N_490[4]), .CK(clk_80mhz), 
            .Q(integrator2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i4.GSR = "ENABLED";
    FD1S3AX integrator2_i5 (.D(integrator2_71__N_490[5]), .CK(clk_80mhz), 
            .Q(integrator2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i5.GSR = "ENABLED";
    FD1S3AX integrator2_i6 (.D(integrator2_71__N_490[6]), .CK(clk_80mhz), 
            .Q(integrator2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i6.GSR = "ENABLED";
    FD1S3AX integrator2_i7 (.D(integrator2_71__N_490[7]), .CK(clk_80mhz), 
            .Q(integrator2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i7.GSR = "ENABLED";
    FD1S3AX integrator2_i8 (.D(integrator2_71__N_490[8]), .CK(clk_80mhz), 
            .Q(integrator2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i8.GSR = "ENABLED";
    FD1S3AX integrator2_i9 (.D(integrator2_71__N_490[9]), .CK(clk_80mhz), 
            .Q(integrator2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i9.GSR = "ENABLED";
    FD1S3AX integrator2_i10 (.D(integrator2_71__N_490[10]), .CK(clk_80mhz), 
            .Q(integrator2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i10.GSR = "ENABLED";
    FD1S3AX integrator2_i11 (.D(integrator2_71__N_490[11]), .CK(clk_80mhz), 
            .Q(integrator2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i11.GSR = "ENABLED";
    FD1S3AX integrator2_i12 (.D(integrator2_71__N_490[12]), .CK(clk_80mhz), 
            .Q(integrator2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i12.GSR = "ENABLED";
    FD1S3AX integrator2_i13 (.D(integrator2_71__N_490[13]), .CK(clk_80mhz), 
            .Q(integrator2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i13.GSR = "ENABLED";
    FD1S3AX integrator2_i14 (.D(integrator2_71__N_490[14]), .CK(clk_80mhz), 
            .Q(integrator2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i14.GSR = "ENABLED";
    FD1S3AX integrator2_i15 (.D(integrator2_71__N_490[15]), .CK(clk_80mhz), 
            .Q(integrator2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i15.GSR = "ENABLED";
    FD1S3AX integrator2_i16 (.D(integrator2_71__N_490[16]), .CK(clk_80mhz), 
            .Q(integrator2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i16.GSR = "ENABLED";
    FD1S3AX integrator2_i17 (.D(integrator2_71__N_490[17]), .CK(clk_80mhz), 
            .Q(integrator2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i17.GSR = "ENABLED";
    FD1S3AX integrator2_i18 (.D(integrator2_71__N_490[18]), .CK(clk_80mhz), 
            .Q(integrator2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i18.GSR = "ENABLED";
    FD1S3AX integrator2_i19 (.D(integrator2_71__N_490[19]), .CK(clk_80mhz), 
            .Q(integrator2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i19.GSR = "ENABLED";
    FD1S3AX integrator2_i20 (.D(integrator2_71__N_490[20]), .CK(clk_80mhz), 
            .Q(integrator2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i20.GSR = "ENABLED";
    FD1S3AX integrator2_i21 (.D(integrator2_71__N_490[21]), .CK(clk_80mhz), 
            .Q(integrator2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i21.GSR = "ENABLED";
    FD1S3AX integrator2_i22 (.D(integrator2_71__N_490[22]), .CK(clk_80mhz), 
            .Q(integrator2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i22.GSR = "ENABLED";
    FD1S3AX integrator2_i23 (.D(integrator2_71__N_490[23]), .CK(clk_80mhz), 
            .Q(integrator2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i23.GSR = "ENABLED";
    FD1S3AX integrator2_i24 (.D(integrator2_71__N_490[24]), .CK(clk_80mhz), 
            .Q(integrator2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i24.GSR = "ENABLED";
    FD1S3AX integrator2_i25 (.D(integrator2_71__N_490[25]), .CK(clk_80mhz), 
            .Q(integrator2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i25.GSR = "ENABLED";
    FD1S3AX integrator2_i26 (.D(integrator2_71__N_490[26]), .CK(clk_80mhz), 
            .Q(integrator2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i26.GSR = "ENABLED";
    FD1S3AX integrator2_i27 (.D(integrator2_71__N_490[27]), .CK(clk_80mhz), 
            .Q(integrator2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i27.GSR = "ENABLED";
    FD1S3AX integrator2_i28 (.D(integrator2_71__N_490[28]), .CK(clk_80mhz), 
            .Q(integrator2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i28.GSR = "ENABLED";
    FD1S3AX integrator2_i29 (.D(integrator2_71__N_490[29]), .CK(clk_80mhz), 
            .Q(integrator2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i29.GSR = "ENABLED";
    FD1S3AX integrator2_i30 (.D(integrator2_71__N_490[30]), .CK(clk_80mhz), 
            .Q(integrator2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i30.GSR = "ENABLED";
    FD1S3AX integrator2_i31 (.D(integrator2_71__N_490[31]), .CK(clk_80mhz), 
            .Q(integrator2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i31.GSR = "ENABLED";
    FD1S3AX integrator2_i32 (.D(integrator2_71__N_490[32]), .CK(clk_80mhz), 
            .Q(integrator2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i32.GSR = "ENABLED";
    FD1S3AX integrator2_i33 (.D(integrator2_71__N_490[33]), .CK(clk_80mhz), 
            .Q(integrator2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i33.GSR = "ENABLED";
    FD1S3AX integrator2_i34 (.D(integrator2_71__N_490[34]), .CK(clk_80mhz), 
            .Q(integrator2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i34.GSR = "ENABLED";
    FD1S3AX integrator2_i35 (.D(integrator2_71__N_490[35]), .CK(clk_80mhz), 
            .Q(integrator2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i35.GSR = "ENABLED";
    FD1S3AX integrator2_i36 (.D(integrator2_71__N_490[36]), .CK(clk_80mhz), 
            .Q(integrator2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i36.GSR = "ENABLED";
    FD1S3AX integrator2_i37 (.D(integrator2_71__N_490[37]), .CK(clk_80mhz), 
            .Q(integrator2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i37.GSR = "ENABLED";
    FD1S3AX integrator2_i38 (.D(integrator2_71__N_490[38]), .CK(clk_80mhz), 
            .Q(integrator2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i38.GSR = "ENABLED";
    FD1S3AX integrator2_i39 (.D(integrator2_71__N_490[39]), .CK(clk_80mhz), 
            .Q(integrator2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i39.GSR = "ENABLED";
    FD1S3AX integrator2_i40 (.D(integrator2_71__N_490[40]), .CK(clk_80mhz), 
            .Q(integrator2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i40.GSR = "ENABLED";
    FD1S3AX integrator2_i41 (.D(integrator2_71__N_490[41]), .CK(clk_80mhz), 
            .Q(integrator2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i41.GSR = "ENABLED";
    FD1S3AX integrator2_i42 (.D(integrator2_71__N_490[42]), .CK(clk_80mhz), 
            .Q(integrator2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i42.GSR = "ENABLED";
    FD1S3AX integrator2_i43 (.D(integrator2_71__N_490[43]), .CK(clk_80mhz), 
            .Q(integrator2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i43.GSR = "ENABLED";
    FD1S3AX integrator2_i44 (.D(integrator2_71__N_490[44]), .CK(clk_80mhz), 
            .Q(integrator2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i44.GSR = "ENABLED";
    FD1S3AX integrator2_i45 (.D(integrator2_71__N_490[45]), .CK(clk_80mhz), 
            .Q(integrator2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i45.GSR = "ENABLED";
    FD1S3AX integrator2_i46 (.D(integrator2_71__N_490[46]), .CK(clk_80mhz), 
            .Q(integrator2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i46.GSR = "ENABLED";
    FD1S3AX integrator2_i47 (.D(integrator2_71__N_490[47]), .CK(clk_80mhz), 
            .Q(integrator2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i47.GSR = "ENABLED";
    FD1S3AX integrator2_i48 (.D(integrator2_71__N_490[48]), .CK(clk_80mhz), 
            .Q(integrator2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i48.GSR = "ENABLED";
    FD1S3AX integrator2_i49 (.D(integrator2_71__N_490[49]), .CK(clk_80mhz), 
            .Q(integrator2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i49.GSR = "ENABLED";
    FD1S3AX integrator2_i50 (.D(integrator2_71__N_490[50]), .CK(clk_80mhz), 
            .Q(integrator2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i50.GSR = "ENABLED";
    FD1S3AX integrator2_i51 (.D(integrator2_71__N_490[51]), .CK(clk_80mhz), 
            .Q(integrator2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i51.GSR = "ENABLED";
    FD1S3AX integrator2_i52 (.D(integrator2_71__N_490[52]), .CK(clk_80mhz), 
            .Q(integrator2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i52.GSR = "ENABLED";
    FD1S3AX integrator2_i53 (.D(integrator2_71__N_490[53]), .CK(clk_80mhz), 
            .Q(integrator2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i53.GSR = "ENABLED";
    FD1S3AX integrator2_i54 (.D(integrator2_71__N_490[54]), .CK(clk_80mhz), 
            .Q(integrator2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i54.GSR = "ENABLED";
    FD1S3AX integrator2_i55 (.D(integrator2_71__N_490[55]), .CK(clk_80mhz), 
            .Q(integrator2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i55.GSR = "ENABLED";
    FD1S3AX integrator2_i56 (.D(integrator2_71__N_490[56]), .CK(clk_80mhz), 
            .Q(integrator2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i56.GSR = "ENABLED";
    FD1S3AX integrator2_i57 (.D(integrator2_71__N_490[57]), .CK(clk_80mhz), 
            .Q(integrator2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i57.GSR = "ENABLED";
    FD1S3AX integrator2_i58 (.D(integrator2_71__N_490[58]), .CK(clk_80mhz), 
            .Q(integrator2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i58.GSR = "ENABLED";
    FD1S3AX integrator2_i59 (.D(integrator2_71__N_490[59]), .CK(clk_80mhz), 
            .Q(integrator2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i59.GSR = "ENABLED";
    FD1S3AX integrator2_i60 (.D(integrator2_71__N_490[60]), .CK(clk_80mhz), 
            .Q(integrator2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i60.GSR = "ENABLED";
    FD1S3AX integrator2_i61 (.D(integrator2_71__N_490[61]), .CK(clk_80mhz), 
            .Q(integrator2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i61.GSR = "ENABLED";
    FD1S3AX integrator2_i62 (.D(integrator2_71__N_490[62]), .CK(clk_80mhz), 
            .Q(integrator2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i62.GSR = "ENABLED";
    FD1S3AX integrator2_i63 (.D(integrator2_71__N_490[63]), .CK(clk_80mhz), 
            .Q(integrator2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i63.GSR = "ENABLED";
    FD1S3AX integrator2_i64 (.D(integrator2_71__N_490[64]), .CK(clk_80mhz), 
            .Q(integrator2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i64.GSR = "ENABLED";
    FD1S3AX integrator2_i65 (.D(integrator2_71__N_490[65]), .CK(clk_80mhz), 
            .Q(integrator2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i65.GSR = "ENABLED";
    FD1S3AX integrator2_i66 (.D(integrator2_71__N_490[66]), .CK(clk_80mhz), 
            .Q(integrator2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i66.GSR = "ENABLED";
    FD1S3AX integrator2_i67 (.D(integrator2_71__N_490[67]), .CK(clk_80mhz), 
            .Q(integrator2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i67.GSR = "ENABLED";
    FD1S3AX integrator2_i68 (.D(integrator2_71__N_490[68]), .CK(clk_80mhz), 
            .Q(integrator2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i68.GSR = "ENABLED";
    FD1S3AX integrator2_i69 (.D(integrator2_71__N_490[69]), .CK(clk_80mhz), 
            .Q(integrator2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i69.GSR = "ENABLED";
    FD1S3AX integrator2_i70 (.D(integrator2_71__N_490[70]), .CK(clk_80mhz), 
            .Q(integrator2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i70.GSR = "ENABLED";
    FD1S3AX integrator2_i71 (.D(integrator2_71__N_490[71]), .CK(clk_80mhz), 
            .Q(integrator2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i71.GSR = "ENABLED";
    FD1S3AX integrator3_i1 (.D(integrator3_71__N_562[1]), .CK(clk_80mhz), 
            .Q(integrator3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i1.GSR = "ENABLED";
    FD1S3AX integrator3_i2 (.D(integrator3_71__N_562[2]), .CK(clk_80mhz), 
            .Q(integrator3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i2.GSR = "ENABLED";
    FD1S3AX integrator3_i3 (.D(integrator3_71__N_562[3]), .CK(clk_80mhz), 
            .Q(integrator3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i3.GSR = "ENABLED";
    FD1S3AX integrator3_i4 (.D(integrator3_71__N_562[4]), .CK(clk_80mhz), 
            .Q(integrator3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i4.GSR = "ENABLED";
    FD1S3AX integrator3_i5 (.D(integrator3_71__N_562[5]), .CK(clk_80mhz), 
            .Q(integrator3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i5.GSR = "ENABLED";
    FD1S3AX integrator3_i6 (.D(integrator3_71__N_562[6]), .CK(clk_80mhz), 
            .Q(integrator3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i6.GSR = "ENABLED";
    FD1S3AX integrator3_i7 (.D(integrator3_71__N_562[7]), .CK(clk_80mhz), 
            .Q(integrator3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i7.GSR = "ENABLED";
    FD1S3AX integrator3_i8 (.D(integrator3_71__N_562[8]), .CK(clk_80mhz), 
            .Q(integrator3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i8.GSR = "ENABLED";
    FD1S3AX integrator3_i9 (.D(integrator3_71__N_562[9]), .CK(clk_80mhz), 
            .Q(integrator3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i9.GSR = "ENABLED";
    FD1S3AX integrator3_i10 (.D(integrator3_71__N_562[10]), .CK(clk_80mhz), 
            .Q(integrator3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i10.GSR = "ENABLED";
    FD1S3AX integrator3_i11 (.D(integrator3_71__N_562[11]), .CK(clk_80mhz), 
            .Q(integrator3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i11.GSR = "ENABLED";
    FD1S3AX integrator3_i12 (.D(integrator3_71__N_562[12]), .CK(clk_80mhz), 
            .Q(integrator3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i12.GSR = "ENABLED";
    FD1S3AX integrator3_i13 (.D(integrator3_71__N_562[13]), .CK(clk_80mhz), 
            .Q(integrator3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i13.GSR = "ENABLED";
    FD1S3AX integrator3_i14 (.D(integrator3_71__N_562[14]), .CK(clk_80mhz), 
            .Q(integrator3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i14.GSR = "ENABLED";
    FD1S3AX integrator3_i15 (.D(integrator3_71__N_562[15]), .CK(clk_80mhz), 
            .Q(integrator3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i15.GSR = "ENABLED";
    FD1S3AX integrator3_i16 (.D(integrator3_71__N_562[16]), .CK(clk_80mhz), 
            .Q(integrator3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i16.GSR = "ENABLED";
    FD1S3AX integrator3_i17 (.D(integrator3_71__N_562[17]), .CK(clk_80mhz), 
            .Q(integrator3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i17.GSR = "ENABLED";
    FD1S3AX integrator3_i18 (.D(integrator3_71__N_562[18]), .CK(clk_80mhz), 
            .Q(integrator3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i18.GSR = "ENABLED";
    FD1S3AX integrator3_i19 (.D(integrator3_71__N_562[19]), .CK(clk_80mhz), 
            .Q(integrator3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i19.GSR = "ENABLED";
    FD1S3AX integrator3_i20 (.D(integrator3_71__N_562[20]), .CK(clk_80mhz), 
            .Q(integrator3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i20.GSR = "ENABLED";
    FD1S3AX integrator3_i21 (.D(integrator3_71__N_562[21]), .CK(clk_80mhz), 
            .Q(integrator3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i21.GSR = "ENABLED";
    FD1S3AX integrator3_i22 (.D(integrator3_71__N_562[22]), .CK(clk_80mhz), 
            .Q(integrator3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i22.GSR = "ENABLED";
    FD1S3AX integrator3_i23 (.D(integrator3_71__N_562[23]), .CK(clk_80mhz), 
            .Q(integrator3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i23.GSR = "ENABLED";
    FD1S3AX integrator3_i24 (.D(integrator3_71__N_562[24]), .CK(clk_80mhz), 
            .Q(integrator3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i24.GSR = "ENABLED";
    FD1S3AX integrator3_i25 (.D(integrator3_71__N_562[25]), .CK(clk_80mhz), 
            .Q(integrator3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i25.GSR = "ENABLED";
    FD1S3AX integrator3_i26 (.D(integrator3_71__N_562[26]), .CK(clk_80mhz), 
            .Q(integrator3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i26.GSR = "ENABLED";
    FD1S3AX integrator3_i27 (.D(integrator3_71__N_562[27]), .CK(clk_80mhz), 
            .Q(integrator3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i27.GSR = "ENABLED";
    FD1S3AX integrator3_i28 (.D(integrator3_71__N_562[28]), .CK(clk_80mhz), 
            .Q(integrator3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i28.GSR = "ENABLED";
    FD1S3AX integrator3_i29 (.D(integrator3_71__N_562[29]), .CK(clk_80mhz), 
            .Q(integrator3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i29.GSR = "ENABLED";
    FD1S3AX integrator3_i30 (.D(integrator3_71__N_562[30]), .CK(clk_80mhz), 
            .Q(integrator3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i30.GSR = "ENABLED";
    FD1S3AX integrator3_i31 (.D(integrator3_71__N_562[31]), .CK(clk_80mhz), 
            .Q(integrator3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i31.GSR = "ENABLED";
    FD1S3AX integrator3_i32 (.D(integrator3_71__N_562[32]), .CK(clk_80mhz), 
            .Q(integrator3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i32.GSR = "ENABLED";
    FD1S3AX integrator3_i33 (.D(integrator3_71__N_562[33]), .CK(clk_80mhz), 
            .Q(integrator3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i33.GSR = "ENABLED";
    FD1S3AX integrator3_i34 (.D(integrator3_71__N_562[34]), .CK(clk_80mhz), 
            .Q(integrator3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i34.GSR = "ENABLED";
    FD1S3AX integrator3_i35 (.D(integrator3_71__N_562[35]), .CK(clk_80mhz), 
            .Q(integrator3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i35.GSR = "ENABLED";
    FD1S3AX integrator3_i36 (.D(integrator3_71__N_562[36]), .CK(clk_80mhz), 
            .Q(integrator3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i36.GSR = "ENABLED";
    FD1S3AX integrator3_i37 (.D(integrator3_71__N_562[37]), .CK(clk_80mhz), 
            .Q(integrator3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i37.GSR = "ENABLED";
    FD1S3AX integrator3_i38 (.D(integrator3_71__N_562[38]), .CK(clk_80mhz), 
            .Q(integrator3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i38.GSR = "ENABLED";
    FD1S3AX integrator3_i39 (.D(integrator3_71__N_562[39]), .CK(clk_80mhz), 
            .Q(integrator3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i39.GSR = "ENABLED";
    FD1S3AX integrator3_i40 (.D(integrator3_71__N_562[40]), .CK(clk_80mhz), 
            .Q(integrator3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i40.GSR = "ENABLED";
    FD1S3AX integrator3_i41 (.D(integrator3_71__N_562[41]), .CK(clk_80mhz), 
            .Q(integrator3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i41.GSR = "ENABLED";
    FD1S3AX integrator3_i42 (.D(integrator3_71__N_562[42]), .CK(clk_80mhz), 
            .Q(integrator3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i42.GSR = "ENABLED";
    FD1S3AX integrator3_i43 (.D(integrator3_71__N_562[43]), .CK(clk_80mhz), 
            .Q(integrator3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i43.GSR = "ENABLED";
    FD1S3AX integrator3_i44 (.D(integrator3_71__N_562[44]), .CK(clk_80mhz), 
            .Q(integrator3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i44.GSR = "ENABLED";
    FD1S3AX integrator3_i45 (.D(integrator3_71__N_562[45]), .CK(clk_80mhz), 
            .Q(integrator3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i45.GSR = "ENABLED";
    FD1S3AX integrator3_i46 (.D(integrator3_71__N_562[46]), .CK(clk_80mhz), 
            .Q(integrator3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i46.GSR = "ENABLED";
    FD1S3AX integrator3_i47 (.D(integrator3_71__N_562[47]), .CK(clk_80mhz), 
            .Q(integrator3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i47.GSR = "ENABLED";
    FD1S3AX integrator3_i48 (.D(integrator3_71__N_562[48]), .CK(clk_80mhz), 
            .Q(integrator3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i48.GSR = "ENABLED";
    FD1S3AX integrator3_i49 (.D(integrator3_71__N_562[49]), .CK(clk_80mhz), 
            .Q(integrator3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i49.GSR = "ENABLED";
    FD1S3AX integrator3_i50 (.D(integrator3_71__N_562[50]), .CK(clk_80mhz), 
            .Q(integrator3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i50.GSR = "ENABLED";
    FD1S3AX integrator3_i51 (.D(integrator3_71__N_562[51]), .CK(clk_80mhz), 
            .Q(integrator3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i51.GSR = "ENABLED";
    FD1S3AX integrator3_i52 (.D(integrator3_71__N_562[52]), .CK(clk_80mhz), 
            .Q(integrator3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i52.GSR = "ENABLED";
    FD1S3AX integrator3_i53 (.D(integrator3_71__N_562[53]), .CK(clk_80mhz), 
            .Q(integrator3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i53.GSR = "ENABLED";
    FD1S3AX integrator3_i54 (.D(integrator3_71__N_562[54]), .CK(clk_80mhz), 
            .Q(integrator3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i54.GSR = "ENABLED";
    FD1S3AX integrator3_i55 (.D(integrator3_71__N_562[55]), .CK(clk_80mhz), 
            .Q(integrator3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i55.GSR = "ENABLED";
    FD1S3AX integrator3_i56 (.D(integrator3_71__N_562[56]), .CK(clk_80mhz), 
            .Q(integrator3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i56.GSR = "ENABLED";
    FD1S3AX integrator3_i57 (.D(integrator3_71__N_562[57]), .CK(clk_80mhz), 
            .Q(integrator3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i57.GSR = "ENABLED";
    FD1S3AX integrator3_i58 (.D(integrator3_71__N_562[58]), .CK(clk_80mhz), 
            .Q(integrator3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i58.GSR = "ENABLED";
    FD1S3AX integrator3_i59 (.D(integrator3_71__N_562[59]), .CK(clk_80mhz), 
            .Q(integrator3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i59.GSR = "ENABLED";
    FD1S3AX integrator3_i60 (.D(integrator3_71__N_562[60]), .CK(clk_80mhz), 
            .Q(integrator3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i60.GSR = "ENABLED";
    FD1S3AX integrator3_i61 (.D(integrator3_71__N_562[61]), .CK(clk_80mhz), 
            .Q(integrator3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i61.GSR = "ENABLED";
    FD1S3AX integrator3_i62 (.D(integrator3_71__N_562[62]), .CK(clk_80mhz), 
            .Q(integrator3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i62.GSR = "ENABLED";
    FD1S3AX integrator3_i63 (.D(integrator3_71__N_562[63]), .CK(clk_80mhz), 
            .Q(integrator3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i63.GSR = "ENABLED";
    FD1S3AX integrator3_i64 (.D(integrator3_71__N_562[64]), .CK(clk_80mhz), 
            .Q(integrator3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i64.GSR = "ENABLED";
    FD1S3AX integrator3_i65 (.D(integrator3_71__N_562[65]), .CK(clk_80mhz), 
            .Q(integrator3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i65.GSR = "ENABLED";
    FD1S3AX integrator3_i66 (.D(integrator3_71__N_562[66]), .CK(clk_80mhz), 
            .Q(integrator3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i66.GSR = "ENABLED";
    FD1S3AX integrator3_i67 (.D(integrator3_71__N_562[67]), .CK(clk_80mhz), 
            .Q(integrator3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i67.GSR = "ENABLED";
    FD1S3AX integrator3_i68 (.D(integrator3_71__N_562[68]), .CK(clk_80mhz), 
            .Q(integrator3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i68.GSR = "ENABLED";
    FD1S3AX integrator3_i69 (.D(integrator3_71__N_562[69]), .CK(clk_80mhz), 
            .Q(integrator3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i69.GSR = "ENABLED";
    FD1S3AX integrator3_i70 (.D(integrator3_71__N_562[70]), .CK(clk_80mhz), 
            .Q(integrator3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i70.GSR = "ENABLED";
    FD1S3AX integrator3_i71 (.D(integrator3_71__N_562[71]), .CK(clk_80mhz), 
            .Q(integrator3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i71.GSR = "ENABLED";
    FD1S3AX integrator4_i1 (.D(integrator4_71__N_634[1]), .CK(clk_80mhz), 
            .Q(integrator4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i1.GSR = "ENABLED";
    FD1S3AX integrator4_i2 (.D(integrator4_71__N_634[2]), .CK(clk_80mhz), 
            .Q(integrator4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i2.GSR = "ENABLED";
    FD1S3AX integrator4_i3 (.D(integrator4_71__N_634[3]), .CK(clk_80mhz), 
            .Q(integrator4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i3.GSR = "ENABLED";
    FD1S3AX integrator4_i4 (.D(integrator4_71__N_634[4]), .CK(clk_80mhz), 
            .Q(integrator4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i4.GSR = "ENABLED";
    FD1S3AX integrator4_i5 (.D(integrator4_71__N_634[5]), .CK(clk_80mhz), 
            .Q(integrator4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i5.GSR = "ENABLED";
    FD1S3AX integrator4_i6 (.D(integrator4_71__N_634[6]), .CK(clk_80mhz), 
            .Q(integrator4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i6.GSR = "ENABLED";
    FD1S3AX integrator4_i7 (.D(integrator4_71__N_634[7]), .CK(clk_80mhz), 
            .Q(integrator4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i7.GSR = "ENABLED";
    FD1S3AX integrator4_i8 (.D(integrator4_71__N_634[8]), .CK(clk_80mhz), 
            .Q(integrator4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i8.GSR = "ENABLED";
    FD1S3AX integrator4_i9 (.D(integrator4_71__N_634[9]), .CK(clk_80mhz), 
            .Q(integrator4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i9.GSR = "ENABLED";
    FD1S3AX integrator4_i10 (.D(integrator4_71__N_634[10]), .CK(clk_80mhz), 
            .Q(integrator4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i10.GSR = "ENABLED";
    FD1S3AX integrator4_i11 (.D(integrator4_71__N_634[11]), .CK(clk_80mhz), 
            .Q(integrator4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i11.GSR = "ENABLED";
    FD1S3AX integrator4_i12 (.D(integrator4_71__N_634[12]), .CK(clk_80mhz), 
            .Q(integrator4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i12.GSR = "ENABLED";
    FD1S3AX integrator4_i13 (.D(integrator4_71__N_634[13]), .CK(clk_80mhz), 
            .Q(integrator4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i13.GSR = "ENABLED";
    FD1S3AX integrator4_i14 (.D(integrator4_71__N_634[14]), .CK(clk_80mhz), 
            .Q(integrator4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i14.GSR = "ENABLED";
    FD1S3AX integrator4_i15 (.D(integrator4_71__N_634[15]), .CK(clk_80mhz), 
            .Q(integrator4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i15.GSR = "ENABLED";
    FD1S3AX integrator4_i16 (.D(integrator4_71__N_634[16]), .CK(clk_80mhz), 
            .Q(integrator4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i16.GSR = "ENABLED";
    FD1S3AX integrator4_i17 (.D(integrator4_71__N_634[17]), .CK(clk_80mhz), 
            .Q(integrator4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i17.GSR = "ENABLED";
    FD1S3AX integrator4_i18 (.D(integrator4_71__N_634[18]), .CK(clk_80mhz), 
            .Q(integrator4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i18.GSR = "ENABLED";
    FD1S3AX integrator4_i19 (.D(integrator4_71__N_634[19]), .CK(clk_80mhz), 
            .Q(integrator4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i19.GSR = "ENABLED";
    FD1S3AX integrator4_i20 (.D(integrator4_71__N_634[20]), .CK(clk_80mhz), 
            .Q(integrator4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i20.GSR = "ENABLED";
    FD1S3AX integrator4_i21 (.D(integrator4_71__N_634[21]), .CK(clk_80mhz), 
            .Q(integrator4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i21.GSR = "ENABLED";
    FD1S3AX integrator4_i22 (.D(integrator4_71__N_634[22]), .CK(clk_80mhz), 
            .Q(integrator4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i22.GSR = "ENABLED";
    FD1S3AX integrator4_i23 (.D(integrator4_71__N_634[23]), .CK(clk_80mhz), 
            .Q(integrator4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i23.GSR = "ENABLED";
    FD1S3AX integrator4_i24 (.D(integrator4_71__N_634[24]), .CK(clk_80mhz), 
            .Q(integrator4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i24.GSR = "ENABLED";
    FD1S3AX integrator4_i25 (.D(integrator4_71__N_634[25]), .CK(clk_80mhz), 
            .Q(integrator4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i25.GSR = "ENABLED";
    FD1S3AX integrator4_i26 (.D(integrator4_71__N_634[26]), .CK(clk_80mhz), 
            .Q(integrator4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i26.GSR = "ENABLED";
    FD1S3AX integrator4_i27 (.D(integrator4_71__N_634[27]), .CK(clk_80mhz), 
            .Q(integrator4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i27.GSR = "ENABLED";
    FD1S3AX integrator4_i28 (.D(integrator4_71__N_634[28]), .CK(clk_80mhz), 
            .Q(integrator4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i28.GSR = "ENABLED";
    FD1S3AX integrator4_i29 (.D(integrator4_71__N_634[29]), .CK(clk_80mhz), 
            .Q(integrator4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i29.GSR = "ENABLED";
    FD1S3AX integrator4_i30 (.D(integrator4_71__N_634[30]), .CK(clk_80mhz), 
            .Q(integrator4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i30.GSR = "ENABLED";
    FD1S3AX integrator4_i31 (.D(integrator4_71__N_634[31]), .CK(clk_80mhz), 
            .Q(integrator4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i31.GSR = "ENABLED";
    FD1S3AX integrator4_i32 (.D(integrator4_71__N_634[32]), .CK(clk_80mhz), 
            .Q(integrator4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i32.GSR = "ENABLED";
    FD1S3AX integrator4_i33 (.D(integrator4_71__N_634[33]), .CK(clk_80mhz), 
            .Q(integrator4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i33.GSR = "ENABLED";
    FD1S3AX integrator4_i34 (.D(integrator4_71__N_634[34]), .CK(clk_80mhz), 
            .Q(integrator4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i34.GSR = "ENABLED";
    FD1S3AX integrator4_i35 (.D(integrator4_71__N_634[35]), .CK(clk_80mhz), 
            .Q(integrator4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i35.GSR = "ENABLED";
    FD1S3AX integrator4_i36 (.D(integrator4_71__N_634[36]), .CK(clk_80mhz), 
            .Q(integrator4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i36.GSR = "ENABLED";
    FD1S3AX integrator4_i37 (.D(integrator4_71__N_634[37]), .CK(clk_80mhz), 
            .Q(integrator4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i37.GSR = "ENABLED";
    FD1S3AX integrator4_i38 (.D(integrator4_71__N_634[38]), .CK(clk_80mhz), 
            .Q(integrator4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i38.GSR = "ENABLED";
    FD1S3AX integrator4_i39 (.D(integrator4_71__N_634[39]), .CK(clk_80mhz), 
            .Q(integrator4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i39.GSR = "ENABLED";
    FD1S3AX integrator4_i40 (.D(integrator4_71__N_634[40]), .CK(clk_80mhz), 
            .Q(integrator4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i40.GSR = "ENABLED";
    FD1S3AX integrator4_i41 (.D(integrator4_71__N_634[41]), .CK(clk_80mhz), 
            .Q(integrator4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i41.GSR = "ENABLED";
    FD1S3AX integrator4_i42 (.D(integrator4_71__N_634[42]), .CK(clk_80mhz), 
            .Q(integrator4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i42.GSR = "ENABLED";
    FD1S3AX integrator4_i43 (.D(integrator4_71__N_634[43]), .CK(clk_80mhz), 
            .Q(integrator4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i43.GSR = "ENABLED";
    FD1S3AX integrator4_i44 (.D(integrator4_71__N_634[44]), .CK(clk_80mhz), 
            .Q(integrator4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i44.GSR = "ENABLED";
    FD1S3AX integrator4_i45 (.D(integrator4_71__N_634[45]), .CK(clk_80mhz), 
            .Q(integrator4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i45.GSR = "ENABLED";
    FD1S3AX integrator4_i46 (.D(integrator4_71__N_634[46]), .CK(clk_80mhz), 
            .Q(integrator4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i46.GSR = "ENABLED";
    FD1S3AX integrator4_i47 (.D(integrator4_71__N_634[47]), .CK(clk_80mhz), 
            .Q(integrator4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i47.GSR = "ENABLED";
    FD1S3AX integrator4_i48 (.D(integrator4_71__N_634[48]), .CK(clk_80mhz), 
            .Q(integrator4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i48.GSR = "ENABLED";
    FD1S3AX integrator4_i49 (.D(integrator4_71__N_634[49]), .CK(clk_80mhz), 
            .Q(integrator4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i49.GSR = "ENABLED";
    FD1S3AX integrator4_i50 (.D(integrator4_71__N_634[50]), .CK(clk_80mhz), 
            .Q(integrator4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i50.GSR = "ENABLED";
    FD1S3AX integrator4_i51 (.D(integrator4_71__N_634[51]), .CK(clk_80mhz), 
            .Q(integrator4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i51.GSR = "ENABLED";
    FD1S3AX integrator4_i52 (.D(integrator4_71__N_634[52]), .CK(clk_80mhz), 
            .Q(integrator4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i52.GSR = "ENABLED";
    FD1S3AX integrator4_i53 (.D(integrator4_71__N_634[53]), .CK(clk_80mhz), 
            .Q(integrator4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i53.GSR = "ENABLED";
    FD1S3AX integrator4_i54 (.D(integrator4_71__N_634[54]), .CK(clk_80mhz), 
            .Q(integrator4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i54.GSR = "ENABLED";
    FD1S3AX integrator4_i55 (.D(integrator4_71__N_634[55]), .CK(clk_80mhz), 
            .Q(integrator4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i55.GSR = "ENABLED";
    FD1S3AX integrator4_i56 (.D(integrator4_71__N_634[56]), .CK(clk_80mhz), 
            .Q(integrator4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i56.GSR = "ENABLED";
    FD1S3AX integrator4_i57 (.D(integrator4_71__N_634[57]), .CK(clk_80mhz), 
            .Q(integrator4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i57.GSR = "ENABLED";
    FD1S3AX integrator4_i58 (.D(integrator4_71__N_634[58]), .CK(clk_80mhz), 
            .Q(integrator4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i58.GSR = "ENABLED";
    FD1S3AX integrator4_i59 (.D(integrator4_71__N_634[59]), .CK(clk_80mhz), 
            .Q(integrator4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i59.GSR = "ENABLED";
    FD1S3AX integrator4_i60 (.D(integrator4_71__N_634[60]), .CK(clk_80mhz), 
            .Q(integrator4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i60.GSR = "ENABLED";
    FD1S3AX integrator4_i61 (.D(integrator4_71__N_634[61]), .CK(clk_80mhz), 
            .Q(integrator4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i61.GSR = "ENABLED";
    FD1S3AX integrator4_i62 (.D(integrator4_71__N_634[62]), .CK(clk_80mhz), 
            .Q(integrator4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i62.GSR = "ENABLED";
    FD1S3AX integrator4_i63 (.D(integrator4_71__N_634[63]), .CK(clk_80mhz), 
            .Q(integrator4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i63.GSR = "ENABLED";
    FD1S3AX integrator4_i64 (.D(integrator4_71__N_634[64]), .CK(clk_80mhz), 
            .Q(integrator4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i64.GSR = "ENABLED";
    FD1S3AX integrator4_i65 (.D(integrator4_71__N_634[65]), .CK(clk_80mhz), 
            .Q(integrator4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i65.GSR = "ENABLED";
    FD1S3AX integrator4_i66 (.D(integrator4_71__N_634[66]), .CK(clk_80mhz), 
            .Q(integrator4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i66.GSR = "ENABLED";
    FD1S3AX integrator4_i67 (.D(integrator4_71__N_634[67]), .CK(clk_80mhz), 
            .Q(integrator4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i67.GSR = "ENABLED";
    FD1S3AX integrator4_i68 (.D(integrator4_71__N_634[68]), .CK(clk_80mhz), 
            .Q(integrator4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i68.GSR = "ENABLED";
    FD1S3AX integrator4_i69 (.D(integrator4_71__N_634[69]), .CK(clk_80mhz), 
            .Q(integrator4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i69.GSR = "ENABLED";
    FD1S3AX integrator4_i70 (.D(integrator4_71__N_634[70]), .CK(clk_80mhz), 
            .Q(integrator4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i70.GSR = "ENABLED";
    FD1S3AX integrator4_i71 (.D(integrator4_71__N_634[71]), .CK(clk_80mhz), 
            .Q(integrator4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i71.GSR = "ENABLED";
    FD1S3AX integrator5_i1 (.D(integrator5_71__N_706[1]), .CK(clk_80mhz), 
            .Q(integrator5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i1.GSR = "ENABLED";
    FD1S3AX integrator5_i2 (.D(integrator5_71__N_706[2]), .CK(clk_80mhz), 
            .Q(integrator5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i2.GSR = "ENABLED";
    FD1S3AX integrator5_i3 (.D(integrator5_71__N_706[3]), .CK(clk_80mhz), 
            .Q(integrator5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i3.GSR = "ENABLED";
    FD1S3AX integrator5_i4 (.D(integrator5_71__N_706[4]), .CK(clk_80mhz), 
            .Q(integrator5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i4.GSR = "ENABLED";
    FD1S3AX integrator5_i5 (.D(integrator5_71__N_706[5]), .CK(clk_80mhz), 
            .Q(integrator5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i5.GSR = "ENABLED";
    FD1S3AX integrator5_i6 (.D(integrator5_71__N_706[6]), .CK(clk_80mhz), 
            .Q(integrator5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i6.GSR = "ENABLED";
    FD1S3AX integrator5_i7 (.D(integrator5_71__N_706[7]), .CK(clk_80mhz), 
            .Q(integrator5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i7.GSR = "ENABLED";
    FD1S3AX integrator5_i8 (.D(integrator5_71__N_706[8]), .CK(clk_80mhz), 
            .Q(integrator5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i8.GSR = "ENABLED";
    FD1S3AX integrator5_i9 (.D(integrator5_71__N_706[9]), .CK(clk_80mhz), 
            .Q(integrator5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i9.GSR = "ENABLED";
    FD1S3AX integrator5_i10 (.D(integrator5_71__N_706[10]), .CK(clk_80mhz), 
            .Q(integrator5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i10.GSR = "ENABLED";
    FD1S3AX integrator5_i11 (.D(integrator5_71__N_706[11]), .CK(clk_80mhz), 
            .Q(integrator5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i11.GSR = "ENABLED";
    FD1S3AX integrator5_i12 (.D(integrator5_71__N_706[12]), .CK(clk_80mhz), 
            .Q(integrator5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i12.GSR = "ENABLED";
    FD1S3AX integrator5_i13 (.D(integrator5_71__N_706[13]), .CK(clk_80mhz), 
            .Q(integrator5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i13.GSR = "ENABLED";
    FD1S3AX integrator5_i14 (.D(integrator5_71__N_706[14]), .CK(clk_80mhz), 
            .Q(integrator5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i14.GSR = "ENABLED";
    FD1S3AX integrator5_i15 (.D(integrator5_71__N_706[15]), .CK(clk_80mhz), 
            .Q(integrator5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i15.GSR = "ENABLED";
    FD1S3AX integrator5_i16 (.D(integrator5_71__N_706[16]), .CK(clk_80mhz), 
            .Q(integrator5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i16.GSR = "ENABLED";
    FD1S3AX integrator5_i17 (.D(integrator5_71__N_706[17]), .CK(clk_80mhz), 
            .Q(integrator5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i17.GSR = "ENABLED";
    FD1S3AX integrator5_i18 (.D(integrator5_71__N_706[18]), .CK(clk_80mhz), 
            .Q(integrator5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i18.GSR = "ENABLED";
    FD1S3AX integrator5_i19 (.D(integrator5_71__N_706[19]), .CK(clk_80mhz), 
            .Q(integrator5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i19.GSR = "ENABLED";
    FD1S3AX integrator5_i20 (.D(integrator5_71__N_706[20]), .CK(clk_80mhz), 
            .Q(integrator5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i20.GSR = "ENABLED";
    FD1S3AX integrator5_i21 (.D(integrator5_71__N_706[21]), .CK(clk_80mhz), 
            .Q(integrator5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i21.GSR = "ENABLED";
    FD1S3AX integrator5_i22 (.D(integrator5_71__N_706[22]), .CK(clk_80mhz), 
            .Q(integrator5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i22.GSR = "ENABLED";
    FD1S3AX integrator5_i23 (.D(integrator5_71__N_706[23]), .CK(clk_80mhz), 
            .Q(integrator5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i23.GSR = "ENABLED";
    FD1S3AX integrator5_i24 (.D(integrator5_71__N_706[24]), .CK(clk_80mhz), 
            .Q(integrator5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i24.GSR = "ENABLED";
    FD1S3AX integrator5_i25 (.D(integrator5_71__N_706[25]), .CK(clk_80mhz), 
            .Q(integrator5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i25.GSR = "ENABLED";
    FD1S3AX integrator5_i26 (.D(integrator5_71__N_706[26]), .CK(clk_80mhz), 
            .Q(integrator5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i26.GSR = "ENABLED";
    FD1S3AX integrator5_i27 (.D(integrator5_71__N_706[27]), .CK(clk_80mhz), 
            .Q(integrator5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i27.GSR = "ENABLED";
    FD1S3AX integrator5_i28 (.D(integrator5_71__N_706[28]), .CK(clk_80mhz), 
            .Q(integrator5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i28.GSR = "ENABLED";
    FD1S3AX integrator5_i29 (.D(integrator5_71__N_706[29]), .CK(clk_80mhz), 
            .Q(integrator5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i29.GSR = "ENABLED";
    FD1S3AX integrator5_i30 (.D(integrator5_71__N_706[30]), .CK(clk_80mhz), 
            .Q(integrator5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i30.GSR = "ENABLED";
    FD1S3AX integrator5_i31 (.D(integrator5_71__N_706[31]), .CK(clk_80mhz), 
            .Q(integrator5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i31.GSR = "ENABLED";
    FD1S3AX integrator5_i32 (.D(integrator5_71__N_706[32]), .CK(clk_80mhz), 
            .Q(integrator5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i32.GSR = "ENABLED";
    FD1S3AX integrator5_i33 (.D(integrator5_71__N_706[33]), .CK(clk_80mhz), 
            .Q(integrator5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i33.GSR = "ENABLED";
    FD1S3AX integrator5_i34 (.D(integrator5_71__N_706[34]), .CK(clk_80mhz), 
            .Q(integrator5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i34.GSR = "ENABLED";
    FD1S3AX integrator5_i35 (.D(integrator5_71__N_706[35]), .CK(clk_80mhz), 
            .Q(integrator5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i35.GSR = "ENABLED";
    FD1S3AX integrator5_i36 (.D(integrator5_71__N_706[36]), .CK(clk_80mhz), 
            .Q(integrator5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i36.GSR = "ENABLED";
    FD1S3AX integrator5_i37 (.D(integrator5_71__N_706[37]), .CK(clk_80mhz), 
            .Q(integrator5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i37.GSR = "ENABLED";
    FD1S3AX integrator5_i38 (.D(integrator5_71__N_706[38]), .CK(clk_80mhz), 
            .Q(integrator5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i38.GSR = "ENABLED";
    FD1S3AX integrator5_i39 (.D(integrator5_71__N_706[39]), .CK(clk_80mhz), 
            .Q(integrator5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i39.GSR = "ENABLED";
    FD1S3AX integrator5_i40 (.D(integrator5_71__N_706[40]), .CK(clk_80mhz), 
            .Q(integrator5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i40.GSR = "ENABLED";
    FD1S3AX integrator5_i41 (.D(integrator5_71__N_706[41]), .CK(clk_80mhz), 
            .Q(integrator5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i41.GSR = "ENABLED";
    FD1S3AX integrator5_i42 (.D(integrator5_71__N_706[42]), .CK(clk_80mhz), 
            .Q(integrator5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i42.GSR = "ENABLED";
    FD1S3AX integrator5_i43 (.D(integrator5_71__N_706[43]), .CK(clk_80mhz), 
            .Q(integrator5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i43.GSR = "ENABLED";
    FD1S3AX integrator5_i44 (.D(integrator5_71__N_706[44]), .CK(clk_80mhz), 
            .Q(integrator5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i44.GSR = "ENABLED";
    FD1S3AX integrator5_i45 (.D(integrator5_71__N_706[45]), .CK(clk_80mhz), 
            .Q(integrator5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i45.GSR = "ENABLED";
    FD1S3AX integrator5_i46 (.D(integrator5_71__N_706[46]), .CK(clk_80mhz), 
            .Q(integrator5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i46.GSR = "ENABLED";
    FD1S3AX integrator5_i47 (.D(integrator5_71__N_706[47]), .CK(clk_80mhz), 
            .Q(integrator5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i47.GSR = "ENABLED";
    FD1S3AX integrator5_i48 (.D(integrator5_71__N_706[48]), .CK(clk_80mhz), 
            .Q(integrator5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i48.GSR = "ENABLED";
    FD1S3AX integrator5_i49 (.D(integrator5_71__N_706[49]), .CK(clk_80mhz), 
            .Q(integrator5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i49.GSR = "ENABLED";
    FD1S3AX integrator5_i50 (.D(integrator5_71__N_706[50]), .CK(clk_80mhz), 
            .Q(integrator5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i50.GSR = "ENABLED";
    FD1S3AX integrator5_i51 (.D(integrator5_71__N_706[51]), .CK(clk_80mhz), 
            .Q(integrator5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i51.GSR = "ENABLED";
    FD1S3AX integrator5_i52 (.D(integrator5_71__N_706[52]), .CK(clk_80mhz), 
            .Q(integrator5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i52.GSR = "ENABLED";
    FD1S3AX integrator5_i53 (.D(integrator5_71__N_706[53]), .CK(clk_80mhz), 
            .Q(integrator5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i53.GSR = "ENABLED";
    FD1S3AX integrator5_i54 (.D(integrator5_71__N_706[54]), .CK(clk_80mhz), 
            .Q(integrator5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i54.GSR = "ENABLED";
    FD1S3AX integrator5_i55 (.D(integrator5_71__N_706[55]), .CK(clk_80mhz), 
            .Q(integrator5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i55.GSR = "ENABLED";
    FD1S3AX integrator5_i56 (.D(integrator5_71__N_706[56]), .CK(clk_80mhz), 
            .Q(integrator5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i56.GSR = "ENABLED";
    FD1S3AX integrator5_i57 (.D(integrator5_71__N_706[57]), .CK(clk_80mhz), 
            .Q(integrator5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i57.GSR = "ENABLED";
    FD1S3AX integrator5_i58 (.D(integrator5_71__N_706[58]), .CK(clk_80mhz), 
            .Q(integrator5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i58.GSR = "ENABLED";
    FD1S3AX integrator5_i59 (.D(integrator5_71__N_706[59]), .CK(clk_80mhz), 
            .Q(integrator5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i59.GSR = "ENABLED";
    FD1S3AX integrator5_i60 (.D(integrator5_71__N_706[60]), .CK(clk_80mhz), 
            .Q(integrator5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i60.GSR = "ENABLED";
    FD1S3AX integrator5_i61 (.D(integrator5_71__N_706[61]), .CK(clk_80mhz), 
            .Q(integrator5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i61.GSR = "ENABLED";
    FD1S3AX integrator5_i62 (.D(integrator5_71__N_706[62]), .CK(clk_80mhz), 
            .Q(integrator5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i62.GSR = "ENABLED";
    FD1S3AX integrator5_i63 (.D(integrator5_71__N_706[63]), .CK(clk_80mhz), 
            .Q(integrator5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i63.GSR = "ENABLED";
    FD1S3AX integrator5_i64 (.D(integrator5_71__N_706[64]), .CK(clk_80mhz), 
            .Q(integrator5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i64.GSR = "ENABLED";
    FD1S3AX integrator5_i65 (.D(integrator5_71__N_706[65]), .CK(clk_80mhz), 
            .Q(integrator5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i65.GSR = "ENABLED";
    FD1S3AX integrator5_i66 (.D(integrator5_71__N_706[66]), .CK(clk_80mhz), 
            .Q(integrator5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i66.GSR = "ENABLED";
    FD1S3AX integrator5_i67 (.D(integrator5_71__N_706[67]), .CK(clk_80mhz), 
            .Q(integrator5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i67.GSR = "ENABLED";
    FD1S3AX integrator5_i68 (.D(integrator5_71__N_706[68]), .CK(clk_80mhz), 
            .Q(integrator5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i68.GSR = "ENABLED";
    FD1S3AX integrator5_i69 (.D(integrator5_71__N_706[69]), .CK(clk_80mhz), 
            .Q(integrator5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i69.GSR = "ENABLED";
    FD1S3AX integrator5_i70 (.D(integrator5_71__N_706[70]), .CK(clk_80mhz), 
            .Q(integrator5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i70.GSR = "ENABLED";
    FD1S3AX integrator5_i71 (.D(integrator5_71__N_706[71]), .CK(clk_80mhz), 
            .Q(integrator5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i71.GSR = "ENABLED";
    FD1P3AX comb6_i0_i1 (.D(comb6_71__N_1451[1]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i1.GSR = "ENABLED";
    FD1P3AX comb6_i0_i2 (.D(comb6_71__N_1451[2]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i2.GSR = "ENABLED";
    FD1P3AX comb6_i0_i3 (.D(comb6_71__N_1451[3]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i3.GSR = "ENABLED";
    FD1P3AX comb6_i0_i4 (.D(comb6_71__N_1451[4]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i4.GSR = "ENABLED";
    FD1P3AX comb6_i0_i5 (.D(comb6_71__N_1451[5]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i5.GSR = "ENABLED";
    FD1P3AX comb6_i0_i6 (.D(comb6_71__N_1451[6]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i6.GSR = "ENABLED";
    FD1P3AX comb6_i0_i7 (.D(comb6_71__N_1451[7]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i7.GSR = "ENABLED";
    FD1P3AX comb6_i0_i8 (.D(comb6_71__N_1451[8]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i8.GSR = "ENABLED";
    FD1P3AX comb6_i0_i9 (.D(comb6_71__N_1451[9]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i9.GSR = "ENABLED";
    FD1P3AX comb6_i0_i10 (.D(comb6_71__N_1451[10]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i10.GSR = "ENABLED";
    FD1P3AX comb6_i0_i11 (.D(comb6_71__N_1451[11]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i11.GSR = "ENABLED";
    FD1P3AX comb6_i0_i12 (.D(comb6_71__N_1451[12]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i12.GSR = "ENABLED";
    FD1P3AX comb6_i0_i13 (.D(comb6_71__N_1451[13]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i13.GSR = "ENABLED";
    FD1P3AX comb6_i0_i14 (.D(comb6_71__N_1451[14]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i14.GSR = "ENABLED";
    FD1P3AX comb6_i0_i15 (.D(comb6_71__N_1451[15]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i15.GSR = "ENABLED";
    FD1P3AX comb6_i0_i16 (.D(comb6_71__N_1451[16]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i16.GSR = "ENABLED";
    FD1P3AX comb6_i0_i17 (.D(comb6_71__N_1451[17]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i17.GSR = "ENABLED";
    FD1P3AX comb6_i0_i18 (.D(comb6_71__N_1451[18]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i18.GSR = "ENABLED";
    FD1P3AX comb6_i0_i19 (.D(comb6_71__N_1451[19]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i19.GSR = "ENABLED";
    FD1P3AX comb6_i0_i20 (.D(comb6_71__N_1451[20]), .SP(clk_80mhz_enable_186), 
            .CK(clk_80mhz), .Q(comb6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i20.GSR = "ENABLED";
    FD1P3AX comb6_i0_i21 (.D(comb6_71__N_1451[21]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i21.GSR = "ENABLED";
    FD1P3AX comb6_i0_i22 (.D(comb6_71__N_1451[22]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i22.GSR = "ENABLED";
    FD1P3AX comb6_i0_i23 (.D(comb6_71__N_1451[23]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i23.GSR = "ENABLED";
    FD1P3AX comb6_i0_i24 (.D(comb6_71__N_1451[24]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i24.GSR = "ENABLED";
    FD1P3AX comb6_i0_i25 (.D(comb6_71__N_1451[25]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i25.GSR = "ENABLED";
    FD1P3AX comb6_i0_i26 (.D(comb6_71__N_1451[26]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i26.GSR = "ENABLED";
    FD1P3AX comb6_i0_i27 (.D(comb6_71__N_1451[27]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i27.GSR = "ENABLED";
    FD1P3AX comb6_i0_i28 (.D(comb6_71__N_1451[28]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i28.GSR = "ENABLED";
    FD1P3AX comb6_i0_i29 (.D(comb6_71__N_1451[29]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i29.GSR = "ENABLED";
    FD1P3AX comb6_i0_i30 (.D(comb6_71__N_1451[30]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i30.GSR = "ENABLED";
    FD1P3AX comb6_i0_i31 (.D(comb6_71__N_1451[31]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i31.GSR = "ENABLED";
    FD1P3AX comb6_i0_i32 (.D(comb6_71__N_1451[32]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i32.GSR = "ENABLED";
    FD1P3AX comb6_i0_i33 (.D(comb6_71__N_1451[33]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i33.GSR = "ENABLED";
    FD1P3AX comb6_i0_i34 (.D(comb6_71__N_1451[34]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i34.GSR = "ENABLED";
    FD1P3AX comb6_i0_i35 (.D(comb6_71__N_1451[35]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i35.GSR = "ENABLED";
    FD1P3AX comb6_i0_i36 (.D(comb6_71__N_1451[36]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i36.GSR = "ENABLED";
    FD1P3AX comb6_i0_i37 (.D(comb6_71__N_1451[37]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i37.GSR = "ENABLED";
    FD1P3AX comb6_i0_i38 (.D(comb6_71__N_1451[38]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i38.GSR = "ENABLED";
    FD1P3AX comb6_i0_i39 (.D(comb6_71__N_1451[39]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i39.GSR = "ENABLED";
    FD1P3AX comb6_i0_i40 (.D(comb6_71__N_1451[40]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i40.GSR = "ENABLED";
    FD1P3AX comb6_i0_i41 (.D(comb6_71__N_1451[41]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i41.GSR = "ENABLED";
    FD1P3AX comb6_i0_i42 (.D(comb6_71__N_1451[42]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i42.GSR = "ENABLED";
    FD1P3AX comb6_i0_i43 (.D(comb6_71__N_1451[43]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i43.GSR = "ENABLED";
    FD1P3AX comb6_i0_i44 (.D(comb6_71__N_1451[44]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i44.GSR = "ENABLED";
    FD1P3AX comb6_i0_i45 (.D(comb6_71__N_1451[45]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i45.GSR = "ENABLED";
    FD1P3AX comb6_i0_i46 (.D(comb6_71__N_1451[46]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i46.GSR = "ENABLED";
    FD1P3AX comb6_i0_i47 (.D(comb6_71__N_1451[47]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i47.GSR = "ENABLED";
    FD1P3AX comb6_i0_i48 (.D(comb6_71__N_1451[48]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i48.GSR = "ENABLED";
    FD1P3AX comb6_i0_i49 (.D(comb6_71__N_1451[49]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i49.GSR = "ENABLED";
    FD1P3AX comb6_i0_i50 (.D(comb6_71__N_1451[50]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i50.GSR = "ENABLED";
    FD1P3AX comb6_i0_i51 (.D(comb6_71__N_1451[51]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i51.GSR = "ENABLED";
    FD1P3AX comb6_i0_i52 (.D(comb6_71__N_1451[52]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i52.GSR = "ENABLED";
    FD1P3AX comb6_i0_i53 (.D(comb6_71__N_1451[53]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i53.GSR = "ENABLED";
    FD1P3AX comb6_i0_i54 (.D(comb6_71__N_1451[54]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i54.GSR = "ENABLED";
    FD1P3AX comb6_i0_i55 (.D(comb6_71__N_1451[55]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i55.GSR = "ENABLED";
    FD1P3AX comb6_i0_i56 (.D(comb6_71__N_1451[56]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i56.GSR = "ENABLED";
    FD1P3AX comb6_i0_i57 (.D(comb6_71__N_1451[57]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i57.GSR = "ENABLED";
    FD1P3AX comb6_i0_i58 (.D(comb6_71__N_1451[58]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i58.GSR = "ENABLED";
    FD1P3AX comb6_i0_i59 (.D(comb6_71__N_1451[59]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i59.GSR = "ENABLED";
    FD1P3AX comb6_i0_i60 (.D(comb6_71__N_1451[60]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i60.GSR = "ENABLED";
    FD1P3AX comb6_i0_i61 (.D(comb6_71__N_1451[61]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i61.GSR = "ENABLED";
    FD1P3AX comb6_i0_i62 (.D(comb6_71__N_1451[62]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i62.GSR = "ENABLED";
    FD1P3AX comb6_i0_i63 (.D(comb6_71__N_1451[63]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i63.GSR = "ENABLED";
    FD1P3AX comb6_i0_i64 (.D(comb6_71__N_1451[64]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i64.GSR = "ENABLED";
    FD1P3AX comb6_i0_i65 (.D(comb6_71__N_1451[65]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i65.GSR = "ENABLED";
    FD1P3AX comb6_i0_i66 (.D(comb6_71__N_1451[66]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i66.GSR = "ENABLED";
    FD1P3AX comb6_i0_i67 (.D(comb6_71__N_1451[67]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i67.GSR = "ENABLED";
    FD1P3AX comb6_i0_i68 (.D(comb6_71__N_1451[68]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i68.GSR = "ENABLED";
    FD1P3AX comb6_i0_i69 (.D(comb6_71__N_1451[69]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i69.GSR = "ENABLED";
    FD1P3AX comb6_i0_i70 (.D(comb6_71__N_1451[70]), .SP(clk_80mhz_enable_236), 
            .CK(clk_80mhz), .Q(comb6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i70.GSR = "ENABLED";
    FD1P3AX comb6_i0_i71 (.D(comb6_71__N_1451[71]), .SP(clk_80mhz_enable_286), 
            .CK(clk_80mhz), .Q(comb6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i1 (.D(comb6[1]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i2 (.D(comb6[2]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i3 (.D(comb6[3]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i4 (.D(comb6[4]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i5 (.D(comb6[5]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i6 (.D(comb6[6]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i7 (.D(comb6[7]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i8 (.D(comb6[8]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i9 (.D(comb6[9]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i10 (.D(comb6[10]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i11 (.D(comb6[11]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i12 (.D(comb6[12]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i13 (.D(comb6[13]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i14 (.D(comb6[14]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i15 (.D(comb6[15]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i16 (.D(comb6[16]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i17 (.D(comb6[17]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i18 (.D(comb6[18]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i19 (.D(comb6[19]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i20 (.D(comb6[20]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i21 (.D(comb6[21]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i22 (.D(comb6[22]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i23 (.D(comb6[23]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i24 (.D(comb6[24]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i25 (.D(comb6[25]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i26 (.D(comb6[26]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i27 (.D(comb6[27]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i28 (.D(comb6[28]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i29 (.D(comb6[29]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i30 (.D(comb6[30]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i31 (.D(comb6[31]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i32 (.D(comb6[32]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i33 (.D(comb6[33]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i34 (.D(comb6[34]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i35 (.D(comb6[35]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i36 (.D(comb6[36]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i37 (.D(comb6[37]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i38 (.D(comb6[38]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i39 (.D(comb6[39]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i40 (.D(comb6[40]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i41 (.D(comb6[41]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i42 (.D(comb6[42]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i43 (.D(comb6[43]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i44 (.D(comb6[44]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i45 (.D(comb6[45]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i46 (.D(comb6[46]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i47 (.D(comb6[47]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i48 (.D(comb6[48]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i49 (.D(comb6[49]), .SP(clk_80mhz_enable_286), .CK(clk_80mhz), 
            .Q(comb_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i50 (.D(comb6[50]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i51 (.D(comb6[51]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i52 (.D(comb6[52]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i53 (.D(comb6[53]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i54 (.D(comb6[54]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i55 (.D(comb6[55]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i56 (.D(comb6[56]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i57 (.D(comb6[57]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i58 (.D(comb6[58]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i59 (.D(comb6[59]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i60 (.D(comb6[60]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i61 (.D(comb6[61]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i62 (.D(comb6[62]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i63 (.D(comb6[63]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i64 (.D(comb6[64]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i65 (.D(comb6[65]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i66 (.D(comb6[66]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i67 (.D(comb6[67]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i68 (.D(comb6[68]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i69 (.D(comb6[69]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i70 (.D(comb6[70]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i71 (.D(comb6[71]), .SP(clk_80mhz_enable_336), .CK(clk_80mhz), 
            .Q(comb_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX comb7_i0_i1 (.D(comb7_71__N_1523[1]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i1.GSR = "ENABLED";
    FD1P3AX comb7_i0_i2 (.D(comb7_71__N_1523[2]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i2.GSR = "ENABLED";
    FD1P3AX comb7_i0_i3 (.D(comb7_71__N_1523[3]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i3.GSR = "ENABLED";
    FD1P3AX comb7_i0_i4 (.D(comb7_71__N_1523[4]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i4.GSR = "ENABLED";
    FD1P3AX comb7_i0_i5 (.D(comb7_71__N_1523[5]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i5.GSR = "ENABLED";
    FD1P3AX comb7_i0_i6 (.D(comb7_71__N_1523[6]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i6.GSR = "ENABLED";
    FD1P3AX comb7_i0_i7 (.D(comb7_71__N_1523[7]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i7.GSR = "ENABLED";
    FD1P3AX comb7_i0_i8 (.D(comb7_71__N_1523[8]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i8.GSR = "ENABLED";
    FD1P3AX comb7_i0_i9 (.D(comb7_71__N_1523[9]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i9.GSR = "ENABLED";
    FD1P3AX comb7_i0_i10 (.D(comb7_71__N_1523[10]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i10.GSR = "ENABLED";
    FD1P3AX comb7_i0_i11 (.D(comb7_71__N_1523[11]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i11.GSR = "ENABLED";
    FD1P3AX comb7_i0_i12 (.D(comb7_71__N_1523[12]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i12.GSR = "ENABLED";
    FD1P3AX comb7_i0_i13 (.D(comb7_71__N_1523[13]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i13.GSR = "ENABLED";
    FD1P3AX comb7_i0_i14 (.D(comb7_71__N_1523[14]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i14.GSR = "ENABLED";
    FD1P3AX comb7_i0_i15 (.D(comb7_71__N_1523[15]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i15.GSR = "ENABLED";
    FD1P3AX comb7_i0_i16 (.D(comb7_71__N_1523[16]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i16.GSR = "ENABLED";
    FD1P3AX comb7_i0_i17 (.D(comb7_71__N_1523[17]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i17.GSR = "ENABLED";
    FD1P3AX comb7_i0_i18 (.D(comb7_71__N_1523[18]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i18.GSR = "ENABLED";
    FD1P3AX comb7_i0_i19 (.D(comb7_71__N_1523[19]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i19.GSR = "ENABLED";
    FD1P3AX comb7_i0_i20 (.D(comb7_71__N_1523[20]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i20.GSR = "ENABLED";
    FD1P3AX comb7_i0_i21 (.D(comb7_71__N_1523[21]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i21.GSR = "ENABLED";
    FD1P3AX comb7_i0_i22 (.D(comb7_71__N_1523[22]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i22.GSR = "ENABLED";
    FD1P3AX comb7_i0_i23 (.D(comb7_71__N_1523[23]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i23.GSR = "ENABLED";
    FD1P3AX comb7_i0_i24 (.D(comb7_71__N_1523[24]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i24.GSR = "ENABLED";
    FD1P3AX comb7_i0_i25 (.D(comb7_71__N_1523[25]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i25.GSR = "ENABLED";
    FD1P3AX comb7_i0_i26 (.D(comb7_71__N_1523[26]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i26.GSR = "ENABLED";
    FD1P3AX comb7_i0_i27 (.D(comb7_71__N_1523[27]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i27.GSR = "ENABLED";
    FD1P3AX comb7_i0_i28 (.D(comb7_71__N_1523[28]), .SP(clk_80mhz_enable_336), 
            .CK(clk_80mhz), .Q(comb7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i28.GSR = "ENABLED";
    FD1P3AX comb7_i0_i29 (.D(comb7_71__N_1523[29]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i29.GSR = "ENABLED";
    FD1P3AX comb7_i0_i30 (.D(comb7_71__N_1523[30]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i30.GSR = "ENABLED";
    FD1P3AX comb7_i0_i31 (.D(comb7_71__N_1523[31]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i31.GSR = "ENABLED";
    FD1P3AX comb7_i0_i32 (.D(comb7_71__N_1523[32]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i32.GSR = "ENABLED";
    FD1P3AX comb7_i0_i33 (.D(comb7_71__N_1523[33]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i33.GSR = "ENABLED";
    FD1P3AX comb7_i0_i34 (.D(comb7_71__N_1523[34]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i34.GSR = "ENABLED";
    FD1P3AX comb7_i0_i35 (.D(comb7_71__N_1523[35]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i35.GSR = "ENABLED";
    FD1P3AX comb7_i0_i36 (.D(comb7_71__N_1523[36]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i36.GSR = "ENABLED";
    FD1P3AX comb7_i0_i37 (.D(comb7_71__N_1523[37]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i37.GSR = "ENABLED";
    FD1P3AX comb7_i0_i38 (.D(comb7_71__N_1523[38]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i38.GSR = "ENABLED";
    FD1P3AX comb7_i0_i39 (.D(comb7_71__N_1523[39]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i39.GSR = "ENABLED";
    FD1P3AX comb7_i0_i40 (.D(comb7_71__N_1523[40]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i40.GSR = "ENABLED";
    FD1P3AX comb7_i0_i41 (.D(comb7_71__N_1523[41]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i41.GSR = "ENABLED";
    FD1P3AX comb7_i0_i42 (.D(comb7_71__N_1523[42]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i42.GSR = "ENABLED";
    FD1P3AX comb7_i0_i43 (.D(comb7_71__N_1523[43]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i43.GSR = "ENABLED";
    FD1P3AX comb7_i0_i44 (.D(comb7_71__N_1523[44]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i44.GSR = "ENABLED";
    FD1P3AX comb7_i0_i45 (.D(comb7_71__N_1523[45]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i45.GSR = "ENABLED";
    FD1P3AX comb7_i0_i46 (.D(comb7_71__N_1523[46]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i46.GSR = "ENABLED";
    FD1P3AX comb7_i0_i47 (.D(comb7_71__N_1523[47]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i47.GSR = "ENABLED";
    FD1P3AX comb7_i0_i48 (.D(comb7_71__N_1523[48]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i48.GSR = "ENABLED";
    FD1P3AX comb7_i0_i49 (.D(comb7_71__N_1523[49]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i49.GSR = "ENABLED";
    FD1P3AX comb7_i0_i50 (.D(comb7_71__N_1523[50]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i50.GSR = "ENABLED";
    FD1P3AX comb7_i0_i51 (.D(comb7_71__N_1523[51]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i51.GSR = "ENABLED";
    FD1P3AX comb7_i0_i52 (.D(comb7_71__N_1523[52]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i52.GSR = "ENABLED";
    FD1P3AX comb7_i0_i53 (.D(comb7_71__N_1523[53]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i53.GSR = "ENABLED";
    FD1P3AX comb7_i0_i54 (.D(comb7_71__N_1523[54]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i54.GSR = "ENABLED";
    FD1P3AX comb7_i0_i55 (.D(comb7_71__N_1523[55]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i55.GSR = "ENABLED";
    FD1P3AX comb7_i0_i56 (.D(comb7_71__N_1523[56]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i56.GSR = "ENABLED";
    FD1P3AX comb7_i0_i57 (.D(comb7_71__N_1523[57]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i57.GSR = "ENABLED";
    FD1P3AX comb7_i0_i58 (.D(comb7_71__N_1523[58]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i58.GSR = "ENABLED";
    FD1P3AX comb7_i0_i59 (.D(comb7_71__N_1523[59]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i59.GSR = "ENABLED";
    FD1P3AX comb7_i0_i60 (.D(comb7_71__N_1523[60]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i60.GSR = "ENABLED";
    FD1P3AX comb7_i0_i61 (.D(comb7_71__N_1523[61]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i61.GSR = "ENABLED";
    FD1P3AX comb7_i0_i62 (.D(comb7_71__N_1523[62]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i62.GSR = "ENABLED";
    FD1P3AX comb7_i0_i63 (.D(comb7_71__N_1523[63]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i63.GSR = "ENABLED";
    FD1P3AX comb7_i0_i64 (.D(comb7_71__N_1523[64]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i64.GSR = "ENABLED";
    FD1P3AX comb7_i0_i65 (.D(comb7_71__N_1523[65]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i65.GSR = "ENABLED";
    FD1P3AX comb7_i0_i66 (.D(comb7_71__N_1523[66]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i66.GSR = "ENABLED";
    FD1P3AX comb7_i0_i67 (.D(comb7_71__N_1523[67]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i67.GSR = "ENABLED";
    FD1P3AX comb7_i0_i68 (.D(comb7_71__N_1523[68]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i68.GSR = "ENABLED";
    FD1P3AX comb7_i0_i69 (.D(comb7_71__N_1523[69]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i69.GSR = "ENABLED";
    FD1P3AX comb7_i0_i70 (.D(comb7_71__N_1523[70]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i70.GSR = "ENABLED";
    FD1P3AX comb7_i0_i71 (.D(comb7_71__N_1523[71]), .SP(clk_80mhz_enable_386), 
            .CK(clk_80mhz), .Q(comb7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i1 (.D(comb7[1]), .SP(clk_80mhz_enable_386), .CK(clk_80mhz), 
            .Q(comb_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i2 (.D(comb7[2]), .SP(clk_80mhz_enable_386), .CK(clk_80mhz), 
            .Q(comb_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i3 (.D(comb7[3]), .SP(clk_80mhz_enable_386), .CK(clk_80mhz), 
            .Q(comb_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i4 (.D(comb7[4]), .SP(clk_80mhz_enable_386), .CK(clk_80mhz), 
            .Q(comb_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i5 (.D(comb7[5]), .SP(clk_80mhz_enable_386), .CK(clk_80mhz), 
            .Q(comb_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i6 (.D(comb7[6]), .SP(clk_80mhz_enable_386), .CK(clk_80mhz), 
            .Q(comb_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i7 (.D(comb7[7]), .SP(clk_80mhz_enable_386), .CK(clk_80mhz), 
            .Q(comb_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i8 (.D(comb7[8]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i9 (.D(comb7[9]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i10 (.D(comb7[10]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i11 (.D(comb7[11]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i12 (.D(comb7[12]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i13 (.D(comb7[13]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i14 (.D(comb7[14]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i15 (.D(comb7[15]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i16 (.D(comb7[16]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i17 (.D(comb7[17]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i18 (.D(comb7[18]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i19 (.D(comb7[19]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i20 (.D(comb7[20]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i21 (.D(comb7[21]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i22 (.D(comb7[22]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i23 (.D(comb7[23]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i24 (.D(comb7[24]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i25 (.D(comb7[25]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i26 (.D(comb7[26]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i27 (.D(comb7[27]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i28 (.D(comb7[28]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i29 (.D(comb7[29]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i30 (.D(comb7[30]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i31 (.D(comb7[31]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i32 (.D(comb7[32]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i33 (.D(comb7[33]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i34 (.D(comb7[34]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i35 (.D(comb7[35]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i36 (.D(comb7[36]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i37 (.D(comb7[37]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i38 (.D(comb7[38]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i39 (.D(comb7[39]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i40 (.D(comb7[40]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i41 (.D(comb7[41]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i42 (.D(comb7[42]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i43 (.D(comb7[43]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i44 (.D(comb7[44]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i45 (.D(comb7[45]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i46 (.D(comb7[46]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i47 (.D(comb7[47]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i48 (.D(comb7[48]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i49 (.D(comb7[49]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i50 (.D(comb7[50]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i51 (.D(comb7[51]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i52 (.D(comb7[52]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i53 (.D(comb7[53]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i54 (.D(comb7[54]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i55 (.D(comb7[55]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i56 (.D(comb7[56]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i57 (.D(comb7[57]), .SP(clk_80mhz_enable_436), .CK(clk_80mhz), 
            .Q(comb_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i58 (.D(comb7[58]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i59 (.D(comb7[59]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i60 (.D(comb7[60]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i61 (.D(comb7[61]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i62 (.D(comb7[62]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i63 (.D(comb7[63]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i64 (.D(comb7[64]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i65 (.D(comb7[65]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i66 (.D(comb7[66]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i67 (.D(comb7[67]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i68 (.D(comb7[68]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i69 (.D(comb7[69]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i70 (.D(comb7[70]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i71 (.D(comb7[71]), .SP(clk_80mhz_enable_486), .CK(clk_80mhz), 
            .Q(comb_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX comb8_i0_i1 (.D(comb8_71__N_1595[1]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i1.GSR = "ENABLED";
    FD1P3AX comb8_i0_i2 (.D(comb8_71__N_1595[2]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i2.GSR = "ENABLED";
    FD1P3AX comb8_i0_i3 (.D(comb8_71__N_1595[3]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i3.GSR = "ENABLED";
    FD1P3AX comb8_i0_i4 (.D(comb8_71__N_1595[4]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i4.GSR = "ENABLED";
    FD1P3AX comb8_i0_i5 (.D(comb8_71__N_1595[5]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i5.GSR = "ENABLED";
    FD1P3AX comb8_i0_i6 (.D(comb8_71__N_1595[6]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i6.GSR = "ENABLED";
    FD1P3AX comb8_i0_i7 (.D(comb8_71__N_1595[7]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i7.GSR = "ENABLED";
    FD1P3AX comb8_i0_i8 (.D(comb8_71__N_1595[8]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i8.GSR = "ENABLED";
    FD1P3AX comb8_i0_i9 (.D(comb8_71__N_1595[9]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i9.GSR = "ENABLED";
    FD1P3AX comb8_i0_i10 (.D(comb8_71__N_1595[10]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i10.GSR = "ENABLED";
    FD1P3AX comb8_i0_i11 (.D(comb8_71__N_1595[11]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i11.GSR = "ENABLED";
    FD1P3AX comb8_i0_i12 (.D(comb8_71__N_1595[12]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i12.GSR = "ENABLED";
    FD1P3AX comb8_i0_i13 (.D(comb8_71__N_1595[13]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i13.GSR = "ENABLED";
    FD1P3AX comb8_i0_i14 (.D(comb8_71__N_1595[14]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i14.GSR = "ENABLED";
    FD1P3AX comb8_i0_i15 (.D(comb8_71__N_1595[15]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i15.GSR = "ENABLED";
    FD1P3AX comb8_i0_i16 (.D(comb8_71__N_1595[16]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i16.GSR = "ENABLED";
    FD1P3AX comb8_i0_i17 (.D(comb8_71__N_1595[17]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i17.GSR = "ENABLED";
    FD1P3AX comb8_i0_i18 (.D(comb8_71__N_1595[18]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i18.GSR = "ENABLED";
    FD1P3AX comb8_i0_i19 (.D(comb8_71__N_1595[19]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i19.GSR = "ENABLED";
    FD1P3AX comb8_i0_i20 (.D(comb8_71__N_1595[20]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i20.GSR = "ENABLED";
    FD1P3AX comb8_i0_i21 (.D(comb8_71__N_1595[21]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i21.GSR = "ENABLED";
    FD1P3AX comb8_i0_i22 (.D(comb8_71__N_1595[22]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i22.GSR = "ENABLED";
    FD1P3AX comb8_i0_i23 (.D(comb8_71__N_1595[23]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i23.GSR = "ENABLED";
    FD1P3AX comb8_i0_i24 (.D(comb8_71__N_1595[24]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i24.GSR = "ENABLED";
    FD1P3AX comb8_i0_i25 (.D(comb8_71__N_1595[25]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i25.GSR = "ENABLED";
    FD1P3AX comb8_i0_i26 (.D(comb8_71__N_1595[26]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i26.GSR = "ENABLED";
    FD1P3AX comb8_i0_i27 (.D(comb8_71__N_1595[27]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i27.GSR = "ENABLED";
    FD1P3AX comb8_i0_i28 (.D(comb8_71__N_1595[28]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i28.GSR = "ENABLED";
    FD1P3AX comb8_i0_i29 (.D(comb8_71__N_1595[29]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i29.GSR = "ENABLED";
    FD1P3AX comb8_i0_i30 (.D(comb8_71__N_1595[30]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i30.GSR = "ENABLED";
    FD1P3AX comb8_i0_i31 (.D(comb8_71__N_1595[31]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i31.GSR = "ENABLED";
    FD1P3AX comb8_i0_i32 (.D(comb8_71__N_1595[32]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i32.GSR = "ENABLED";
    FD1P3AX comb8_i0_i33 (.D(comb8_71__N_1595[33]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i33.GSR = "ENABLED";
    FD1P3AX comb8_i0_i34 (.D(comb8_71__N_1595[34]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i34.GSR = "ENABLED";
    FD1P3AX comb8_i0_i35 (.D(comb8_71__N_1595[35]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i35.GSR = "ENABLED";
    FD1P3AX comb8_i0_i36 (.D(comb8_71__N_1595[36]), .SP(clk_80mhz_enable_486), 
            .CK(clk_80mhz), .Q(comb8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i36.GSR = "ENABLED";
    FD1P3AX comb8_i0_i37 (.D(comb8_71__N_1595[37]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i37.GSR = "ENABLED";
    FD1P3AX comb8_i0_i38 (.D(comb8_71__N_1595[38]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i38.GSR = "ENABLED";
    FD1P3AX comb8_i0_i39 (.D(comb8_71__N_1595[39]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i39.GSR = "ENABLED";
    FD1P3AX comb8_i0_i40 (.D(comb8_71__N_1595[40]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i40.GSR = "ENABLED";
    FD1P3AX comb8_i0_i41 (.D(comb8_71__N_1595[41]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i41.GSR = "ENABLED";
    FD1P3AX comb8_i0_i42 (.D(comb8_71__N_1595[42]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i42.GSR = "ENABLED";
    FD1P3AX comb8_i0_i43 (.D(comb8_71__N_1595[43]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i43.GSR = "ENABLED";
    FD1P3AX comb8_i0_i44 (.D(comb8_71__N_1595[44]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i44.GSR = "ENABLED";
    FD1P3AX comb8_i0_i45 (.D(comb8_71__N_1595[45]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i45.GSR = "ENABLED";
    FD1P3AX comb8_i0_i46 (.D(comb8_71__N_1595[46]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i46.GSR = "ENABLED";
    FD1P3AX comb8_i0_i47 (.D(comb8_71__N_1595[47]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i47.GSR = "ENABLED";
    FD1P3AX comb8_i0_i48 (.D(comb8_71__N_1595[48]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i48.GSR = "ENABLED";
    FD1P3AX comb8_i0_i49 (.D(comb8_71__N_1595[49]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i49.GSR = "ENABLED";
    FD1P3AX comb8_i0_i50 (.D(comb8_71__N_1595[50]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i50.GSR = "ENABLED";
    FD1P3AX comb8_i0_i51 (.D(comb8_71__N_1595[51]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i51.GSR = "ENABLED";
    FD1P3AX comb8_i0_i52 (.D(comb8_71__N_1595[52]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i52.GSR = "ENABLED";
    FD1P3AX comb8_i0_i53 (.D(comb8_71__N_1595[53]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i53.GSR = "ENABLED";
    FD1P3AX comb8_i0_i54 (.D(comb8_71__N_1595[54]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i54.GSR = "ENABLED";
    FD1P3AX comb8_i0_i55 (.D(comb8_71__N_1595[55]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i55.GSR = "ENABLED";
    FD1P3AX comb8_i0_i56 (.D(comb8_71__N_1595[56]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i56.GSR = "ENABLED";
    FD1P3AX comb8_i0_i57 (.D(comb8_71__N_1595[57]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i57.GSR = "ENABLED";
    FD1P3AX comb8_i0_i58 (.D(comb8_71__N_1595[58]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i58.GSR = "ENABLED";
    FD1P3AX comb8_i0_i59 (.D(comb8_71__N_1595[59]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i59.GSR = "ENABLED";
    FD1P3AX comb8_i0_i60 (.D(comb8_71__N_1595[60]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i60.GSR = "ENABLED";
    FD1P3AX comb8_i0_i61 (.D(comb8_71__N_1595[61]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i61.GSR = "ENABLED";
    FD1P3AX comb8_i0_i62 (.D(comb8_71__N_1595[62]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i62.GSR = "ENABLED";
    FD1P3AX comb8_i0_i63 (.D(comb8_71__N_1595[63]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i63.GSR = "ENABLED";
    FD1P3AX comb8_i0_i64 (.D(comb8_71__N_1595[64]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i64.GSR = "ENABLED";
    FD1P3AX comb8_i0_i65 (.D(comb8_71__N_1595[65]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i65.GSR = "ENABLED";
    FD1P3AX comb8_i0_i66 (.D(comb8_71__N_1595[66]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i66.GSR = "ENABLED";
    FD1P3AX comb8_i0_i67 (.D(comb8_71__N_1595[67]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i67.GSR = "ENABLED";
    FD1P3AX comb8_i0_i68 (.D(comb8_71__N_1595[68]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i68.GSR = "ENABLED";
    FD1P3AX comb8_i0_i69 (.D(comb8_71__N_1595[69]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i69.GSR = "ENABLED";
    FD1P3AX comb8_i0_i70 (.D(comb8_71__N_1595[70]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i70.GSR = "ENABLED";
    FD1P3AX comb8_i0_i71 (.D(comb8_71__N_1595[71]), .SP(clk_80mhz_enable_536), 
            .CK(clk_80mhz), .Q(comb8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i1 (.D(comb8[1]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i2 (.D(comb8[2]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i3 (.D(comb8[3]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i4 (.D(comb8[4]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i5 (.D(comb8[5]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i6 (.D(comb8[6]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i7 (.D(comb8[7]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i8 (.D(comb8[8]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i9 (.D(comb8[9]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i10 (.D(comb8[10]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i11 (.D(comb8[11]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i12 (.D(comb8[12]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i13 (.D(comb8[13]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i14 (.D(comb8[14]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i15 (.D(comb8[15]), .SP(clk_80mhz_enable_536), .CK(clk_80mhz), 
            .Q(comb_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i16 (.D(comb8[16]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i17 (.D(comb8[17]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i18 (.D(comb8[18]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i19 (.D(comb8[19]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i20 (.D(comb8[20]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i21 (.D(comb8[21]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i22 (.D(comb8[22]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i23 (.D(comb8[23]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i24 (.D(comb8[24]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i25 (.D(comb8[25]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i26 (.D(comb8[26]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i27 (.D(comb8[27]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i28 (.D(comb8[28]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i29 (.D(comb8[29]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i30 (.D(comb8[30]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i31 (.D(comb8[31]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i32 (.D(comb8[32]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i33 (.D(comb8[33]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i34 (.D(comb8[34]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i35 (.D(comb8[35]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i36 (.D(comb8[36]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i37 (.D(comb8[37]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i38 (.D(comb8[38]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i39 (.D(comb8[39]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i40 (.D(comb8[40]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i41 (.D(comb8[41]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i42 (.D(comb8[42]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i43 (.D(comb8[43]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i44 (.D(comb8[44]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i45 (.D(comb8[45]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i46 (.D(comb8[46]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i47 (.D(comb8[47]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i48 (.D(comb8[48]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i49 (.D(comb8[49]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i50 (.D(comb8[50]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i51 (.D(comb8[51]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i52 (.D(comb8[52]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i53 (.D(comb8[53]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i54 (.D(comb8[54]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i55 (.D(comb8[55]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i56 (.D(comb8[56]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i57 (.D(comb8[57]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i58 (.D(comb8[58]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i59 (.D(comb8[59]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i60 (.D(comb8[60]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i61 (.D(comb8[61]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i62 (.D(comb8[62]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i63 (.D(comb8[63]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i64 (.D(comb8[64]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i65 (.D(comb8[65]), .SP(clk_80mhz_enable_586), .CK(clk_80mhz), 
            .Q(comb_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i66 (.D(comb8[66]), .SP(clk_80mhz_enable_636), .CK(clk_80mhz), 
            .Q(comb_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i67 (.D(comb8[67]), .SP(clk_80mhz_enable_636), .CK(clk_80mhz), 
            .Q(comb_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i68 (.D(comb8[68]), .SP(clk_80mhz_enable_636), .CK(clk_80mhz), 
            .Q(comb_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i69 (.D(comb8[69]), .SP(clk_80mhz_enable_636), .CK(clk_80mhz), 
            .Q(comb_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i70 (.D(comb8[70]), .SP(clk_80mhz_enable_636), .CK(clk_80mhz), 
            .Q(comb_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i71 (.D(comb8[71]), .SP(clk_80mhz_enable_636), .CK(clk_80mhz), 
            .Q(comb_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX comb9_i0_i1 (.D(comb9_71__N_1667[1]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i1.GSR = "ENABLED";
    FD1P3AX comb9_i0_i2 (.D(comb9_71__N_1667[2]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i2.GSR = "ENABLED";
    FD1P3AX comb9_i0_i3 (.D(comb9_71__N_1667[3]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i3.GSR = "ENABLED";
    FD1P3AX comb9_i0_i4 (.D(comb9_71__N_1667[4]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i4.GSR = "ENABLED";
    FD1P3AX comb9_i0_i5 (.D(comb9_71__N_1667[5]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i5.GSR = "ENABLED";
    FD1P3AX comb9_i0_i6 (.D(comb9_71__N_1667[6]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i6.GSR = "ENABLED";
    FD1P3AX comb9_i0_i7 (.D(comb9_71__N_1667[7]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i7.GSR = "ENABLED";
    FD1P3AX comb9_i0_i8 (.D(comb9_71__N_1667[8]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i8.GSR = "ENABLED";
    FD1P3AX comb9_i0_i9 (.D(comb9_71__N_1667[9]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i9.GSR = "ENABLED";
    FD1P3AX comb9_i0_i10 (.D(comb9_71__N_1667[10]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i10.GSR = "ENABLED";
    FD1P3AX comb9_i0_i11 (.D(comb9_71__N_1667[11]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i11.GSR = "ENABLED";
    FD1P3AX comb9_i0_i12 (.D(comb9_71__N_1667[12]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i12.GSR = "ENABLED";
    FD1P3AX comb9_i0_i13 (.D(comb9_71__N_1667[13]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i13.GSR = "ENABLED";
    FD1P3AX comb9_i0_i14 (.D(comb9_71__N_1667[14]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i14.GSR = "ENABLED";
    FD1P3AX comb9_i0_i15 (.D(comb9_71__N_1667[15]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i15.GSR = "ENABLED";
    FD1P3AX comb9_i0_i16 (.D(comb9_71__N_1667[16]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i16.GSR = "ENABLED";
    FD1P3AX comb9_i0_i17 (.D(comb9_71__N_1667[17]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i17.GSR = "ENABLED";
    FD1P3AX comb9_i0_i18 (.D(comb9_71__N_1667[18]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i18.GSR = "ENABLED";
    FD1P3AX comb9_i0_i19 (.D(comb9_71__N_1667[19]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i19.GSR = "ENABLED";
    FD1P3AX comb9_i0_i20 (.D(comb9_71__N_1667[20]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i20.GSR = "ENABLED";
    FD1P3AX comb9_i0_i21 (.D(comb9_71__N_1667[21]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i21.GSR = "ENABLED";
    FD1P3AX comb9_i0_i22 (.D(comb9_71__N_1667[22]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i22.GSR = "ENABLED";
    FD1P3AX comb9_i0_i23 (.D(comb9_71__N_1667[23]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i23.GSR = "ENABLED";
    FD1P3AX comb9_i0_i24 (.D(comb9_71__N_1667[24]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i24.GSR = "ENABLED";
    FD1P3AX comb9_i0_i25 (.D(comb9_71__N_1667[25]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i25.GSR = "ENABLED";
    FD1P3AX comb9_i0_i26 (.D(comb9_71__N_1667[26]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i26.GSR = "ENABLED";
    FD1P3AX comb9_i0_i27 (.D(comb9_71__N_1667[27]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i27.GSR = "ENABLED";
    FD1P3AX comb9_i0_i28 (.D(comb9_71__N_1667[28]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i28.GSR = "ENABLED";
    FD1P3AX comb9_i0_i29 (.D(comb9_71__N_1667[29]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i29.GSR = "ENABLED";
    FD1P3AX comb9_i0_i30 (.D(comb9_71__N_1667[30]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i30.GSR = "ENABLED";
    FD1P3AX comb9_i0_i31 (.D(comb9_71__N_1667[31]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i31.GSR = "ENABLED";
    FD1P3AX comb9_i0_i32 (.D(comb9_71__N_1667[32]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i32.GSR = "ENABLED";
    FD1P3AX comb9_i0_i33 (.D(comb9_71__N_1667[33]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i33.GSR = "ENABLED";
    FD1P3AX comb9_i0_i34 (.D(comb9_71__N_1667[34]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i34.GSR = "ENABLED";
    FD1P3AX comb9_i0_i35 (.D(comb9_71__N_1667[35]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i35.GSR = "ENABLED";
    FD1P3AX comb9_i0_i36 (.D(comb9_71__N_1667[36]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i36.GSR = "ENABLED";
    FD1P3AX comb9_i0_i37 (.D(comb9_71__N_1667[37]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i37.GSR = "ENABLED";
    FD1P3AX comb9_i0_i38 (.D(comb9_71__N_1667[38]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i38.GSR = "ENABLED";
    FD1P3AX comb9_i0_i39 (.D(comb9_71__N_1667[39]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i39.GSR = "ENABLED";
    FD1P3AX comb9_i0_i40 (.D(comb9_71__N_1667[40]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i40.GSR = "ENABLED";
    FD1P3AX comb9_i0_i41 (.D(comb9_71__N_1667[41]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i41.GSR = "ENABLED";
    FD1P3AX comb9_i0_i42 (.D(comb9_71__N_1667[42]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i42.GSR = "ENABLED";
    FD1P3AX comb9_i0_i43 (.D(comb9_71__N_1667[43]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i43.GSR = "ENABLED";
    FD1P3AX comb9_i0_i44 (.D(comb9_71__N_1667[44]), .SP(clk_80mhz_enable_636), 
            .CK(clk_80mhz), .Q(comb9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i44.GSR = "ENABLED";
    FD1P3AX comb9_i0_i45 (.D(comb9_71__N_1667[45]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i45.GSR = "ENABLED";
    FD1P3AX comb9_i0_i46 (.D(comb9_71__N_1667[46]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i46.GSR = "ENABLED";
    FD1P3AX comb9_i0_i47 (.D(comb9_71__N_1667[47]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i47.GSR = "ENABLED";
    FD1P3AX comb9_i0_i48 (.D(comb9_71__N_1667[48]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i48.GSR = "ENABLED";
    FD1P3AX comb9_i0_i49 (.D(comb9_71__N_1667[49]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i49.GSR = "ENABLED";
    FD1P3AX comb9_i0_i50 (.D(comb9_71__N_1667[50]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i50.GSR = "ENABLED";
    FD1P3AX comb9_i0_i51 (.D(comb9_71__N_1667[51]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i51.GSR = "ENABLED";
    FD1P3AX comb9_i0_i52 (.D(comb9_71__N_1667[52]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i52.GSR = "ENABLED";
    FD1P3AX comb9_i0_i53 (.D(comb9_71__N_1667[53]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i53.GSR = "ENABLED";
    FD1P3AX comb9_i0_i54 (.D(comb9_71__N_1667[54]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i54.GSR = "ENABLED";
    FD1P3AX comb9_i0_i55 (.D(comb9_71__N_1667[55]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i55.GSR = "ENABLED";
    FD1P3AX comb9_i0_i56 (.D(comb9_71__N_1667[56]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i56.GSR = "ENABLED";
    FD1P3AX comb9_i0_i57 (.D(comb9_71__N_1667[57]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i57.GSR = "ENABLED";
    FD1P3AX comb9_i0_i58 (.D(comb9_71__N_1667[58]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i58.GSR = "ENABLED";
    FD1P3AX comb9_i0_i59 (.D(comb9_71__N_1667[59]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i59.GSR = "ENABLED";
    FD1P3AX comb9_i0_i60 (.D(comb9_71__N_1667[60]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i60.GSR = "ENABLED";
    FD1P3AX comb9_i0_i61 (.D(comb9_71__N_1667[61]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i61.GSR = "ENABLED";
    FD1P3AX comb9_i0_i62 (.D(comb9_71__N_1667[62]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i62.GSR = "ENABLED";
    FD1P3AX comb9_i0_i63 (.D(comb9_71__N_1667[63]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i63.GSR = "ENABLED";
    FD1P3AX comb9_i0_i64 (.D(comb9_71__N_1667[64]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i64.GSR = "ENABLED";
    FD1P3AX comb9_i0_i65 (.D(comb9_71__N_1667[65]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i65.GSR = "ENABLED";
    FD1P3AX comb9_i0_i66 (.D(comb9_71__N_1667[66]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i66.GSR = "ENABLED";
    FD1P3AX comb9_i0_i67 (.D(comb9_71__N_1667[67]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i67.GSR = "ENABLED";
    FD1P3AX comb9_i0_i68 (.D(comb9_71__N_1667[68]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i68.GSR = "ENABLED";
    FD1P3AX comb9_i0_i69 (.D(comb9_71__N_1667[69]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i69.GSR = "ENABLED";
    FD1P3AX comb9_i0_i70 (.D(comb9_71__N_1667[70]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i70.GSR = "ENABLED";
    FD1P3AX comb9_i0_i71 (.D(comb9_71__N_1667[71]), .SP(clk_80mhz_enable_686), 
            .CK(clk_80mhz), .Q(comb9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i1 (.D(comb9[1]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i2 (.D(comb9[2]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i3 (.D(comb9[3]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i4 (.D(comb9[4]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i5 (.D(comb9[5]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i6 (.D(comb9[6]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i7 (.D(comb9[7]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i8 (.D(comb9[8]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i9 (.D(comb9[9]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i10 (.D(comb9[10]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i11 (.D(comb9[11]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i12 (.D(comb9[12]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i13 (.D(comb9[13]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i14 (.D(comb9[14]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i15 (.D(comb9[15]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i16 (.D(comb9[16]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i17 (.D(comb9[17]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i18 (.D(comb9[18]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i19 (.D(comb9[19]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i20 (.D(comb9[20]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i21 (.D(comb9[21]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i22 (.D(comb9[22]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i23 (.D(comb9[23]), .SP(clk_80mhz_enable_686), .CK(clk_80mhz), 
            .Q(comb_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i24 (.D(comb9[24]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i25 (.D(comb9[25]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i26 (.D(comb9[26]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i27 (.D(comb9[27]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i28 (.D(comb9[28]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i29 (.D(comb9[29]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i30 (.D(comb9[30]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i31 (.D(comb9[31]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i32 (.D(comb9[32]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i33 (.D(comb9[33]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i34 (.D(comb9[34]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i35 (.D(comb9[35]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i36 (.D(comb9[36]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i37 (.D(comb9[37]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i38 (.D(comb9[38]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i39 (.D(comb9[39]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i40 (.D(comb9[40]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i41 (.D(comb9[41]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i42 (.D(comb9[42]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i43 (.D(comb9[43]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i44 (.D(comb9[44]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i45 (.D(comb9[45]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i46 (.D(comb9[46]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i47 (.D(comb9[47]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i48 (.D(comb9[48]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i49 (.D(comb9[49]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i50 (.D(comb9[50]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i51 (.D(comb9[51]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i52 (.D(comb9[52]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i53 (.D(comb9[53]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i54 (.D(comb9[54]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i55 (.D(comb9[55]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i56 (.D(comb9[56]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i57 (.D(comb9[57]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i58 (.D(comb9[58]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i59 (.D(comb9[59]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i60 (.D(comb9[60]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i61 (.D(comb9[61]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i62 (.D(comb9[62]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i63 (.D(comb9[63]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i64 (.D(comb9[64]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i65 (.D(comb9[65]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i66 (.D(comb9[66]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i67 (.D(comb9[67]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i68 (.D(comb9[68]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i69 (.D(comb9[69]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i70 (.D(comb9[70]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i71 (.D(comb9[71]), .SP(clk_80mhz_enable_736), .CK(clk_80mhz), 
            .Q(comb_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX comb10__i2 (.D(comb10_71__N_1739[57]), .SP(clk_80mhz_enable_736), 
            .CK(clk_80mhz), .Q(comb10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i2.GSR = "ENABLED";
    FD1P3AX comb10__i3 (.D(comb10_71__N_1739[58]), .SP(clk_80mhz_enable_736), 
            .CK(clk_80mhz), .Q(comb10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i3.GSR = "ENABLED";
    FD1P3AX comb10__i4 (.D(comb10_71__N_1739[59]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i4.GSR = "ENABLED";
    FD1P3AX comb10__i5 (.D(comb10_71__N_1739[60]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i5.GSR = "ENABLED";
    FD1P3AX comb10__i6 (.D(comb10_71__N_1739[61]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i6.GSR = "ENABLED";
    FD1P3AX comb10__i7 (.D(comb10_71__N_1739[62]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i7.GSR = "ENABLED";
    FD1P3AX comb10__i8 (.D(comb10_71__N_1739[63]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i8.GSR = "ENABLED";
    FD1P3AX comb10__i9 (.D(comb10_71__N_1739[64]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i9.GSR = "ENABLED";
    FD1P3AX comb10__i10 (.D(comb10_71__N_1739[65]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i10.GSR = "ENABLED";
    FD1P3AX comb10__i11 (.D(comb10_71__N_1739[66]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i11.GSR = "ENABLED";
    FD1P3AX comb10__i12 (.D(comb10_71__N_1739[67]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i12.GSR = "ENABLED";
    FD1P3AX comb10__i13 (.D(comb10_71__N_1739[68]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i13.GSR = "ENABLED";
    FD1P3AX comb10__i14 (.D(comb10_71__N_1739[69]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i14.GSR = "ENABLED";
    FD1P3AX comb10__i15 (.D(comb10_71__N_1739[70]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i15.GSR = "ENABLED";
    FD1P3AX comb10__i16 (.D(comb10_71__N_1739[71]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i16.GSR = "ENABLED";
    FD1P3AX data_out_i0_i1 (.D(data_out_11__N_1811[1]), .SP(clk_80mhz_enable_737), 
            .CK(clk_80mhz), .Q(mult_i_b[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i1.GSR = "ENABLED";
    FD1P3AX data_out_i0_i2 (.D(data_out_11__N_1811[2]), .SP(clk_80mhz_enable_738), 
            .CK(clk_80mhz), .Q(mult_i_b[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i2.GSR = "ENABLED";
    FD1P3AX data_out_i0_i3 (.D(data_out_11__N_1811[3]), .SP(clk_80mhz_enable_739), 
            .CK(clk_80mhz), .Q(mult_i_b[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i3.GSR = "ENABLED";
    FD1P3AX data_out_i0_i4 (.D(data_out_11__N_1811[4]), .SP(clk_80mhz_enable_740), 
            .CK(clk_80mhz), .Q(mult_i_b[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i4.GSR = "ENABLED";
    FD1P3AX data_out_i0_i5 (.D(data_out_11__N_1811[5]), .SP(clk_80mhz_enable_741), 
            .CK(clk_80mhz), .Q(mult_i_b[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i5.GSR = "ENABLED";
    FD1P3AX data_out_i0_i6 (.D(data_out_11__N_1811[6]), .SP(clk_80mhz_enable_742), 
            .CK(clk_80mhz), .Q(mult_i_b[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i6.GSR = "ENABLED";
    FD1P3AX data_out_i0_i7 (.D(data_out_11__N_1811[7]), .SP(clk_80mhz_enable_743), 
            .CK(clk_80mhz), .Q(mult_i_b[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i7.GSR = "ENABLED";
    FD1P3AX data_out_i0_i8 (.D(data_out_11__N_1811[8]), .SP(clk_80mhz_enable_744), 
            .CK(clk_80mhz), .Q(mult_i_b[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i8.GSR = "ENABLED";
    FD1P3AX data_out_i0_i9 (.D(data_out_11__N_1811[9]), .SP(clk_80mhz_enable_745), 
            .CK(clk_80mhz), .Q(mult_i_b[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i9.GSR = "ENABLED";
    FD1P3AX data_out_i0_i10 (.D(data_out_11__N_1811[10]), .SP(clk_80mhz_enable_746), 
            .CK(clk_80mhz), .Q(mult_i_b[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i10.GSR = "ENABLED";
    FD1P3AX data_out_i0_i11 (.D(data_out_11__N_1811[11]), .SP(clk_80mhz_enable_747), 
            .CK(clk_80mhz), .Q(mult_i_b[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i11.GSR = "ENABLED";
    FD1S3AX integrator1_i1 (.D(integrator1_71__N_418[1]), .CK(clk_80mhz), 
            .Q(integrator1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i1.GSR = "ENABLED";
    FD1S3AX integrator1_i2 (.D(integrator1_71__N_418[2]), .CK(clk_80mhz), 
            .Q(integrator1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i2.GSR = "ENABLED";
    FD1S3AX integrator1_i3 (.D(integrator1_71__N_418[3]), .CK(clk_80mhz), 
            .Q(integrator1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i3.GSR = "ENABLED";
    FD1S3AX integrator1_i4 (.D(integrator1_71__N_418[4]), .CK(clk_80mhz), 
            .Q(integrator1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i4.GSR = "ENABLED";
    FD1S3AX integrator1_i5 (.D(integrator1_71__N_418[5]), .CK(clk_80mhz), 
            .Q(integrator1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i5.GSR = "ENABLED";
    FD1S3AX integrator1_i6 (.D(integrator1_71__N_418[6]), .CK(clk_80mhz), 
            .Q(integrator1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i6.GSR = "ENABLED";
    FD1S3AX integrator1_i7 (.D(integrator1_71__N_418[7]), .CK(clk_80mhz), 
            .Q(integrator1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i7.GSR = "ENABLED";
    FD1S3AX integrator1_i8 (.D(integrator1_71__N_418[8]), .CK(clk_80mhz), 
            .Q(integrator1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i8.GSR = "ENABLED";
    FD1S3AX integrator1_i9 (.D(integrator1_71__N_418[9]), .CK(clk_80mhz), 
            .Q(integrator1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i9.GSR = "ENABLED";
    FD1S3AX integrator1_i10 (.D(integrator1_71__N_418[10]), .CK(clk_80mhz), 
            .Q(integrator1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i10.GSR = "ENABLED";
    FD1S3AX integrator1_i11 (.D(integrator1_71__N_418[11]), .CK(clk_80mhz), 
            .Q(integrator1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i11.GSR = "ENABLED";
    FD1S3AX integrator1_i12 (.D(integrator1_71__N_418[12]), .CK(clk_80mhz), 
            .Q(integrator1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i12.GSR = "ENABLED";
    FD1S3AX integrator1_i13 (.D(integrator1_71__N_418[13]), .CK(clk_80mhz), 
            .Q(integrator1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i13.GSR = "ENABLED";
    FD1S3AX integrator1_i14 (.D(integrator1_71__N_418[14]), .CK(clk_80mhz), 
            .Q(integrator1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i14.GSR = "ENABLED";
    FD1S3AX integrator1_i15 (.D(integrator1_71__N_418[15]), .CK(clk_80mhz), 
            .Q(integrator1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i15.GSR = "ENABLED";
    FD1S3AX integrator1_i16 (.D(integrator1_71__N_418[16]), .CK(clk_80mhz), 
            .Q(integrator1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i16.GSR = "ENABLED";
    FD1S3AX integrator1_i17 (.D(integrator1_71__N_418[17]), .CK(clk_80mhz), 
            .Q(integrator1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i17.GSR = "ENABLED";
    FD1S3AX integrator1_i18 (.D(integrator1_71__N_418[18]), .CK(clk_80mhz), 
            .Q(integrator1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i18.GSR = "ENABLED";
    FD1S3AX integrator1_i19 (.D(integrator1_71__N_418[19]), .CK(clk_80mhz), 
            .Q(integrator1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i19.GSR = "ENABLED";
    FD1S3AX integrator1_i20 (.D(integrator1_71__N_418[20]), .CK(clk_80mhz), 
            .Q(integrator1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i20.GSR = "ENABLED";
    FD1S3AX integrator1_i21 (.D(integrator1_71__N_418[21]), .CK(clk_80mhz), 
            .Q(integrator1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i21.GSR = "ENABLED";
    FD1S3AX integrator1_i22 (.D(integrator1_71__N_418[22]), .CK(clk_80mhz), 
            .Q(integrator1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i22.GSR = "ENABLED";
    FD1S3AX integrator1_i23 (.D(integrator1_71__N_418[23]), .CK(clk_80mhz), 
            .Q(integrator1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i23.GSR = "ENABLED";
    FD1S3AX integrator1_i24 (.D(integrator1_71__N_418[24]), .CK(clk_80mhz), 
            .Q(integrator1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i24.GSR = "ENABLED";
    FD1S3AX integrator1_i25 (.D(integrator1_71__N_418[25]), .CK(clk_80mhz), 
            .Q(integrator1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i25.GSR = "ENABLED";
    FD1S3AX integrator1_i26 (.D(integrator1_71__N_418[26]), .CK(clk_80mhz), 
            .Q(integrator1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i26.GSR = "ENABLED";
    FD1S3AX integrator1_i27 (.D(integrator1_71__N_418[27]), .CK(clk_80mhz), 
            .Q(integrator1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i27.GSR = "ENABLED";
    FD1S3AX integrator1_i28 (.D(integrator1_71__N_418[28]), .CK(clk_80mhz), 
            .Q(integrator1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i28.GSR = "ENABLED";
    FD1S3AX integrator1_i29 (.D(integrator1_71__N_418[29]), .CK(clk_80mhz), 
            .Q(integrator1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i29.GSR = "ENABLED";
    FD1S3AX integrator1_i30 (.D(integrator1_71__N_418[30]), .CK(clk_80mhz), 
            .Q(integrator1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i30.GSR = "ENABLED";
    FD1S3AX integrator1_i31 (.D(integrator1_71__N_418[31]), .CK(clk_80mhz), 
            .Q(integrator1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i31.GSR = "ENABLED";
    FD1S3AX integrator1_i32 (.D(integrator1_71__N_418[32]), .CK(clk_80mhz), 
            .Q(integrator1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i32.GSR = "ENABLED";
    FD1S3AX integrator1_i33 (.D(integrator1_71__N_418[33]), .CK(clk_80mhz), 
            .Q(integrator1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i33.GSR = "ENABLED";
    FD1S3AX integrator1_i34 (.D(integrator1_71__N_418[34]), .CK(clk_80mhz), 
            .Q(integrator1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i34.GSR = "ENABLED";
    FD1S3AX integrator1_i35 (.D(integrator1_71__N_418[35]), .CK(clk_80mhz), 
            .Q(integrator1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i35.GSR = "ENABLED";
    FD1S3AX integrator1_i36 (.D(integrator1_71__N_418[36]), .CK(clk_80mhz), 
            .Q(integrator1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i36.GSR = "ENABLED";
    FD1S3AX integrator1_i37 (.D(integrator1_71__N_418[37]), .CK(clk_80mhz), 
            .Q(integrator1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i37.GSR = "ENABLED";
    FD1S3AX integrator1_i38 (.D(integrator1_71__N_418[38]), .CK(clk_80mhz), 
            .Q(integrator1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i38.GSR = "ENABLED";
    FD1S3AX integrator1_i39 (.D(integrator1_71__N_418[39]), .CK(clk_80mhz), 
            .Q(integrator1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i39.GSR = "ENABLED";
    FD1S3AX integrator1_i40 (.D(integrator1_71__N_418[40]), .CK(clk_80mhz), 
            .Q(integrator1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i40.GSR = "ENABLED";
    FD1S3AX integrator1_i41 (.D(integrator1_71__N_418[41]), .CK(clk_80mhz), 
            .Q(integrator1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i41.GSR = "ENABLED";
    FD1S3AX integrator1_i42 (.D(integrator1_71__N_418[42]), .CK(clk_80mhz), 
            .Q(integrator1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i42.GSR = "ENABLED";
    FD1S3AX integrator1_i43 (.D(integrator1_71__N_418[43]), .CK(clk_80mhz), 
            .Q(integrator1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i43.GSR = "ENABLED";
    FD1S3AX integrator1_i44 (.D(integrator1_71__N_418[44]), .CK(clk_80mhz), 
            .Q(integrator1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i44.GSR = "ENABLED";
    FD1S3AX integrator1_i45 (.D(integrator1_71__N_418[45]), .CK(clk_80mhz), 
            .Q(integrator1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i45.GSR = "ENABLED";
    FD1S3AX integrator1_i46 (.D(integrator1_71__N_418[46]), .CK(clk_80mhz), 
            .Q(integrator1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i46.GSR = "ENABLED";
    FD1S3AX integrator1_i47 (.D(integrator1_71__N_418[47]), .CK(clk_80mhz), 
            .Q(integrator1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i47.GSR = "ENABLED";
    FD1S3AX integrator1_i48 (.D(integrator1_71__N_418[48]), .CK(clk_80mhz), 
            .Q(integrator1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i48.GSR = "ENABLED";
    FD1S3AX integrator1_i49 (.D(integrator1_71__N_418[49]), .CK(clk_80mhz), 
            .Q(integrator1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i49.GSR = "ENABLED";
    FD1S3AX integrator1_i50 (.D(integrator1_71__N_418[50]), .CK(clk_80mhz), 
            .Q(integrator1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i50.GSR = "ENABLED";
    FD1S3AX integrator1_i51 (.D(integrator1_71__N_418[51]), .CK(clk_80mhz), 
            .Q(integrator1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i51.GSR = "ENABLED";
    FD1S3AX integrator1_i52 (.D(integrator1_71__N_418[52]), .CK(clk_80mhz), 
            .Q(integrator1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i52.GSR = "ENABLED";
    FD1S3AX integrator1_i53 (.D(integrator1_71__N_418[53]), .CK(clk_80mhz), 
            .Q(integrator1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i53.GSR = "ENABLED";
    FD1S3AX integrator1_i54 (.D(integrator1_71__N_418[54]), .CK(clk_80mhz), 
            .Q(integrator1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i54.GSR = "ENABLED";
    FD1S3AX integrator1_i55 (.D(integrator1_71__N_418[55]), .CK(clk_80mhz), 
            .Q(integrator1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i55.GSR = "ENABLED";
    FD1S3AX integrator1_i56 (.D(integrator1_71__N_418[56]), .CK(clk_80mhz), 
            .Q(integrator1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i56.GSR = "ENABLED";
    FD1S3AX integrator1_i57 (.D(integrator1_71__N_418[57]), .CK(clk_80mhz), 
            .Q(integrator1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i57.GSR = "ENABLED";
    FD1S3AX integrator1_i58 (.D(integrator1_71__N_418[58]), .CK(clk_80mhz), 
            .Q(integrator1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i58.GSR = "ENABLED";
    FD1S3AX integrator1_i59 (.D(integrator1_71__N_418[59]), .CK(clk_80mhz), 
            .Q(integrator1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i59.GSR = "ENABLED";
    FD1S3AX integrator1_i60 (.D(integrator1_71__N_418[60]), .CK(clk_80mhz), 
            .Q(integrator1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i60.GSR = "ENABLED";
    FD1S3AX integrator1_i61 (.D(integrator1_71__N_418[61]), .CK(clk_80mhz), 
            .Q(integrator1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i61.GSR = "ENABLED";
    FD1S3AX integrator1_i62 (.D(integrator1_71__N_418[62]), .CK(clk_80mhz), 
            .Q(integrator1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i62.GSR = "ENABLED";
    FD1S3AX integrator1_i63 (.D(integrator1_71__N_418[63]), .CK(clk_80mhz), 
            .Q(integrator1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i63.GSR = "ENABLED";
    FD1S3AX integrator1_i64 (.D(integrator1_71__N_418[64]), .CK(clk_80mhz), 
            .Q(integrator1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i64.GSR = "ENABLED";
    FD1S3AX integrator1_i65 (.D(integrator1_71__N_418[65]), .CK(clk_80mhz), 
            .Q(integrator1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i65.GSR = "ENABLED";
    FD1S3AX integrator1_i66 (.D(integrator1_71__N_418[66]), .CK(clk_80mhz), 
            .Q(integrator1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i66.GSR = "ENABLED";
    FD1S3AX integrator1_i67 (.D(integrator1_71__N_418[67]), .CK(clk_80mhz), 
            .Q(integrator1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i67.GSR = "ENABLED";
    FD1S3AX integrator1_i68 (.D(integrator1_71__N_418[68]), .CK(clk_80mhz), 
            .Q(integrator1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i68.GSR = "ENABLED";
    FD1S3AX integrator1_i69 (.D(integrator1_71__N_418[69]), .CK(clk_80mhz), 
            .Q(integrator1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i69.GSR = "ENABLED";
    FD1S3AX integrator1_i70 (.D(integrator1_71__N_418[70]), .CK(clk_80mhz), 
            .Q(integrator1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i70.GSR = "ENABLED";
    FD1S3AX integrator1_i71 (.D(integrator1_71__N_418[71]), .CK(clk_80mhz), 
            .Q(integrator1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i71.GSR = "ENABLED";
    FD1S3IX count__i2 (.D(n67[2]), .CK(clk_80mhz), .CD(n11935), .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n67[3]), .CK(clk_80mhz), .CD(n11935), .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n67[4]), .CK(clk_80mhz), .CD(n11935), .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n67[5]), .CK(clk_80mhz), .CD(n11935), .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n67[6]), .CK(clk_80mhz), .CD(n11935), .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n67[7]), .CK(clk_80mhz), .CD(n11935), .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n67[8]), .CK(clk_80mhz), .CD(n11935), .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n67[9]), .CK(clk_80mhz), .CD(n11935), .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n67[10]), .CK(clk_80mhz), .CD(n11935), .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_11__N_1438[11]), .CK(clk_80mhz), .CD(decimation_clk_N_1823), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i11.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_380 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_743)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_380.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_379 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_742)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_379.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i71_1_lut (.A(comb_d7[70]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i72_1_lut (.A(comb_d7[71]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i69_1_lut (.A(comb_d7[68]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i70_1_lut (.A(comb_d7[69]), .Z(n4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i67_1_lut (.A(comb_d7[66]), .Z(n7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 i1_2_lut (.A(n73), .B(decimation_clk), .Z(n11887)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(60[32:37])
    defparam i1_2_lut.init = 16'h8888;
    FD1S3AX valid_comb_66_rep_378 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_741)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_378.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(count[11]), .B(n16525), .C(n16509), .D(n16517), 
         .Z(n73)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut.init = 16'hfffd;
    LUT4 shift_right_31_i70_rep_204_3_lut (.A(comb10[69]), .B(comb10[70]), 
         .C(\cic_gain[0] ), .Z(n16626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i70_rep_204_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_177 (.A(count[2]), .B(n16521), .C(count[5]), .D(count[9]), 
         .Z(n16525)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_177.init = 16'hfffe;
    LUT4 i1_2_lut_adj_178 (.A(count[0]), .B(count[8]), .Z(n16509)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_178.init = 16'heeee;
    LUT4 i1_2_lut_adj_179 (.A(count[6]), .B(count[3]), .Z(n16517)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_179.init = 16'heeee;
    LUT4 i1_4_lut_adj_180 (.A(count[7]), .B(count[4]), .C(count[1]), .D(count[10]), 
         .Z(n16521)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_180.init = 16'hfffe;
    LUT4 i1_2_lut_adj_181 (.A(n67[11]), .B(n73), .Z(count_11__N_1438[11])) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_181.init = 16'hbbbb;
    LUT4 sub_27_inv_0_i68_1_lut (.A(comb_d7[67]), .Z(n6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i61_rep_228_3_lut (.A(comb10[60]), .B(comb10[61]), 
         .C(\cic_gain[0] ), .Z(n16650)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i61_rep_228_3_lut.init = 16'hcaca;
    LUT4 sub_27_inv_0_i65_1_lut (.A(comb_d7[64]), .Z(n9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i66_1_lut (.A(comb_d7[65]), .Z(n8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i63_1_lut (.A(comb_d7[62]), .Z(n11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i64_1_lut (.A(comb_d7[63]), .Z(n10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i61_1_lut (.A(comb_d7[60]), .Z(n13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i62_1_lut (.A(comb_d7[61]), .Z(n12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i59_1_lut (.A(comb_d7[58]), .Z(n15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i60_1_lut (.A(comb_d7[59]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i57_1_lut (.A(comb_d7[56]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i58_1_lut (.A(comb_d7[57]), .Z(n16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i55_1_lut (.A(comb_d7[54]), .Z(n19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i56_1_lut (.A(comb_d7[55]), .Z(n18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i53_1_lut (.A(comb_d7[52]), .Z(n21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i54_1_lut (.A(comb_d7[53]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i51_1_lut (.A(comb_d7[50]), .Z(n23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i52_1_lut (.A(comb_d7[51]), .Z(n22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i49_1_lut (.A(comb_d7[48]), .Z(n25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i50_1_lut (.A(comb_d7[49]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i47_1_lut (.A(comb_d7[46]), .Z(n27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i48_1_lut (.A(comb_d7[47]), .Z(n26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i45_1_lut (.A(comb_d7[44]), .Z(n29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i46_1_lut (.A(comb_d7[45]), .Z(n28_adj_115)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i43_1_lut (.A(comb_d7[42]), .Z(n31_adj_116)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i44_1_lut (.A(comb_d7[43]), .Z(n30_adj_117)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i41_1_lut (.A(comb_d7[40]), .Z(n33_adj_118)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i42_1_lut (.A(comb_d7[41]), .Z(n32_adj_119)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i39_1_lut (.A(comb_d7[38]), .Z(n35_adj_120)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i40_1_lut (.A(comb_d7[39]), .Z(n34_adj_121)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i37_1_lut (.A(comb_d7[36]), .Z(n37_adj_122)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i38_1_lut (.A(comb_d7[37]), .Z(n36_adj_123)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i38_1_lut.init = 16'h5555;
    FD1S3AX valid_comb_66_rep_382 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_745)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_382.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_182 (.A(n67[0]), .B(n73), .Z(count_11__N_1438[0])) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_182.init = 16'hbbbb;
    LUT4 i1_4_lut_rep_399 (.A(n16569), .B(count[10]), .C(n16553), .D(count[11]), 
         .Z(n17316)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam i1_4_lut_rep_399.init = 16'h8000;
    LUT4 i1_2_lut_adj_183 (.A(n17316), .B(n73), .Z(n11935)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_183.init = 16'hbbbb;
    FD1S3AX valid_comb_66_rep_377 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_740)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_377.GSR = "ENABLED";
    LUT4 i1_4_lut_rep_400 (.A(n16569), .B(count[10]), .C(n16553), .D(count[11]), 
         .Z(clk_80mhz_enable_99)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam i1_4_lut_rep_400.init = 16'h8000;
    FD1S3AX valid_comb_66_rep_398 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_736)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_398.GSR = "ENABLED";
    LUT4 i1_4_lut_rep_401 (.A(n16569), .B(count[10]), .C(n16553), .D(count[11]), 
         .Z(clk_80mhz_enable_149)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam i1_4_lut_rep_401.init = 16'h8000;
    FD1S3AX valid_comb_66_rep_397 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_686)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_397.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_396 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_636)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_396.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_184 (.A(n16569), .B(count[10]), .C(n16553), .D(count[11]), 
         .Z(decimation_clk_N_1823)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam i1_4_lut_adj_184.init = 16'h8000;
    FD1S3AX valid_comb_66_rep_395 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_586)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_395.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_394 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_536)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_394.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_393 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_486)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_393.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_392 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_436)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_392.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_391 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_386)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_391.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_390 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_336)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_390.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_389 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_286)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_389.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_388 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_236)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_388.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_387 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_186)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_387.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_386 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1508)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_386.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_185 (.A(count[8]), .B(n16565), .C(n16551), .D(count[3]), 
         .Z(n16569)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam i1_4_lut_adj_185.init = 16'h8000;
    LUT4 i1_2_lut_adj_186 (.A(count[1]), .B(count[0]), .Z(n16553)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam i1_2_lut_adj_186.init = 16'h8888;
    LUT4 i1_4_lut_adj_187 (.A(count[4]), .B(count[5]), .C(count[2]), .D(count[7]), 
         .Z(n16565)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam i1_4_lut_adj_187.init = 16'h8000;
    LUT4 i1_2_lut_adj_188 (.A(count[9]), .B(count[6]), .Z(n16551)) /* synthesis lut_function=(A (B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam i1_2_lut_adj_188.init = 16'h8888;
    FD1S3AX valid_comb_66_rep_376 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_739)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_376.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_375 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_738)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_375.GSR = "ENABLED";
    PFUMX i5840 (.BLUT(n17206), .ALUT(n17207), .C0(\cic_gain[0] ), .Z(data_out_11__N_1811[0]));
    PFUMX i5838 (.BLUT(n17203), .ALUT(n17204), .C0(\cic_gain[0] ), .Z(data_out_11__N_1811[1]));
    PFUMX i5836 (.BLUT(n17200), .ALUT(n17201), .C0(\cic_gain[0] ), .Z(data_out_11__N_1811[9]));
    LUT4 sub_26_inv_0_i71_1_lut (.A(comb_d6[70]), .Z(n3_adj_124)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i71_1_lut.init = 16'h5555;
    FD1S3AX valid_comb_66_rep_384 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_747)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_384.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i72_1_lut (.A(comb_d6[71]), .Z(n2_adj_125)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i69_1_lut (.A(comb_d6[68]), .Z(n5_adj_126)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i70_1_lut (.A(comb_d6[69]), .Z(n4_adj_127)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i71_1_lut (.A(comb_d8[70]), .Z(n3_adj_128)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i72_1_lut (.A(comb_d8[71]), .Z(n2_adj_129)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i69_1_lut (.A(comb_d8[68]), .Z(n5_adj_130)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i70_1_lut (.A(comb_d8[69]), .Z(n4_adj_131)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i70_1_lut.init = 16'h5555;
    PFUMX i5834 (.BLUT(n17197), .ALUT(n17198), .C0(\cic_gain[0] ), .Z(data_out_11__N_1811[10]));
    LUT4 sub_28_inv_0_i67_1_lut (.A(comb_d8[66]), .Z(n7_adj_132)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i68_1_lut (.A(comb_d8[67]), .Z(n6_adj_133)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i65_1_lut (.A(comb_d8[64]), .Z(n9_adj_134)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i66_1_lut (.A(comb_d8[65]), .Z(n8_adj_135)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i63_1_lut (.A(comb_d8[62]), .Z(n11_adj_136)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i64_1_lut (.A(comb_d8[63]), .Z(n10_adj_137)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i61_1_lut (.A(comb_d8[60]), .Z(n13_adj_138)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i62_1_lut (.A(comb_d8[61]), .Z(n12_adj_139)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i59_1_lut (.A(comb_d8[58]), .Z(n15_adj_140)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i60_1_lut (.A(comb_d8[59]), .Z(n14_adj_141)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i57_1_lut (.A(comb_d8[56]), .Z(n17_adj_142)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i58_1_lut (.A(comb_d8[57]), .Z(n16_adj_143)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i55_1_lut (.A(comb_d8[54]), .Z(n19_adj_144)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i56_1_lut (.A(comb_d8[55]), .Z(n18_adj_145)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i56_1_lut.init = 16'h5555;
    PFUMX i5832 (.BLUT(n17194), .ALUT(n17195), .C0(comb10[71]), .Z(data_out_11__N_1811[11]));
    LUT4 sub_28_inv_0_i53_1_lut (.A(comb_d8[52]), .Z(n21_adj_146)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i54_1_lut (.A(comb_d8[53]), .Z(n20_adj_147)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i67_1_lut (.A(comb_d6[66]), .Z(n7_adj_148)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i68_1_lut (.A(comb_d6[67]), .Z(n6_adj_149)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i65_1_lut (.A(comb_d6[64]), .Z(n9_adj_150)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i66_1_lut (.A(comb_d6[65]), .Z(n8_adj_151)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i63_1_lut (.A(comb_d6[62]), .Z(n11_adj_152)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i64_1_lut (.A(comb_d6[63]), .Z(n10_adj_153)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i61_1_lut (.A(comb_d6[60]), .Z(n13_adj_154)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i62_1_lut (.A(comb_d6[61]), .Z(n12_adj_155)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i59_1_lut (.A(comb_d6[58]), .Z(n15_adj_156)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i60_1_lut (.A(comb_d6[59]), .Z(n14_adj_157)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i57_1_lut (.A(comb_d6[56]), .Z(n17_adj_158)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i58_1_lut (.A(comb_d6[57]), .Z(n16_adj_159)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i55_1_lut (.A(comb_d6[54]), .Z(n19_adj_160)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i55_1_lut.init = 16'h5555;
    PFUMX i5830 (.BLUT(n17191), .ALUT(n17192), .C0(\cic_gain[0] ), .Z(\data_out_11__N_1811[10] ));
    LUT4 sub_26_inv_0_i56_1_lut (.A(comb_d6[55]), .Z(n18_adj_161)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i53_1_lut (.A(comb_d6[52]), .Z(n21_adj_162)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i54_1_lut (.A(comb_d6[53]), .Z(n20_adj_163)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i51_1_lut (.A(comb_d6[50]), .Z(n23_adj_164)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i52_1_lut (.A(comb_d6[51]), .Z(n22_adj_165)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i51_1_lut (.A(comb_d8[50]), .Z(n23_adj_166)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i52_1_lut (.A(comb_d8[51]), .Z(n22_adj_167)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i49_1_lut (.A(comb_d8[48]), .Z(n25_adj_168)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i50_1_lut (.A(comb_d8[49]), .Z(n24_adj_169)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i47_1_lut (.A(comb_d8[46]), .Z(n27_adj_170)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i47_1_lut.init = 16'h5555;
    PFUMX i5828 (.BLUT(n17188), .ALUT(n17189), .C0(\cic_gain[0] ), .Z(\data_out_11__N_1811[11] ));
    LUT4 sub_28_inv_0_i48_1_lut (.A(comb_d8[47]), .Z(n26_adj_171)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i45_1_lut (.A(comb_d8[44]), .Z(n29_adj_172)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i46_1_lut (.A(comb_d8[45]), .Z(n28_adj_173)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i43_1_lut (.A(comb_d8[42]), .Z(n31_adj_174)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i44_1_lut (.A(comb_d8[43]), .Z(n30_adj_175)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i49_1_lut (.A(comb_d6[48]), .Z(n25_adj_176)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i50_1_lut (.A(comb_d6[49]), .Z(n24_adj_177)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i41_1_lut (.A(comb_d8[40]), .Z(n33_adj_178)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i42_1_lut (.A(comb_d8[41]), .Z(n32_adj_179)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i39_1_lut (.A(comb_d8[38]), .Z(n35_adj_180)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i40_1_lut (.A(comb_d8[39]), .Z(n34_adj_181)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i37_1_lut (.A(comb_d8[36]), .Z(n37_adj_182)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i38_1_lut (.A(comb_d8[37]), .Z(n36_adj_183)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i38_1_lut.init = 16'h5555;
    PFUMX i5826 (.BLUT(n17185), .ALUT(n17186), .C0(\cic_gain[1] ), .Z(data_out_11__N_1811[8]));
    LUT4 sub_26_inv_0_i47_1_lut (.A(comb_d6[46]), .Z(n27_adj_184)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i48_1_lut (.A(comb_d6[47]), .Z(n26_adj_185)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i45_1_lut (.A(comb_d6[44]), .Z(n29_adj_186)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i46_1_lut (.A(comb_d6[45]), .Z(n28_adj_187)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i43_1_lut (.A(comb_d6[42]), .Z(n31_adj_188)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i44_1_lut (.A(comb_d6[43]), .Z(n30_adj_189)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i41_1_lut (.A(comb_d6[40]), .Z(n33_adj_190)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i42_1_lut (.A(comb_d6[41]), .Z(n32_adj_191)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i39_1_lut (.A(comb_d6[38]), .Z(n35_adj_192)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i40_1_lut (.A(comb_d6[39]), .Z(n34_adj_193)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i37_1_lut (.A(comb_d6[36]), .Z(n37_adj_194)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i38_1_lut (.A(comb_d6[37]), .Z(n36_adj_195)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i38_1_lut.init = 16'h5555;
    PFUMX i5824 (.BLUT(n17182), .ALUT(n17183), .C0(\cic_gain[1] ), .Z(\data_out_11__N_1811[8] ));
    LUT4 sub_25_inv_0_i71_1_lut (.A(integrator_d_tmp[70]), .Z(n3_adj_196)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i72_1_lut (.A(integrator_d_tmp[71]), .Z(n2_adj_197)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i69_1_lut (.A(integrator_d_tmp[68]), .Z(n5_adj_198)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i69_1_lut.init = 16'h5555;
    FD1S3AX valid_comb_66_rep_383 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_746)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_383.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i70_1_lut (.A(integrator_d_tmp[69]), .Z(n4_adj_199)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i67_1_lut (.A(integrator_d_tmp[66]), .Z(n7_adj_200)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i67_1_lut.init = 16'h5555;
    PFUMX i5822 (.BLUT(n17179), .ALUT(n17180), .C0(\cic_gain[1] ), .Z(\data_out_11__N_1811[9] ));
    LUT4 sub_25_inv_0_i68_1_lut (.A(integrator_d_tmp[67]), .Z(n6_adj_201)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i68_1_lut.init = 16'h5555;
    FD1P3AX integrator_d_tmp_i0_i56 (.D(integrator_tmp[56]), .SP(clk_80mhz_enable_1508), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i56.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i65_1_lut (.A(integrator_d_tmp[64]), .Z(n9_adj_202)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i66_1_lut (.A(integrator_d_tmp[65]), .Z(n8_adj_203)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i63_1_lut (.A(integrator_d_tmp[62]), .Z(n11_adj_204)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i64_1_lut (.A(integrator_d_tmp[63]), .Z(n10_adj_205)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i61_1_lut (.A(integrator_d_tmp[60]), .Z(n13_adj_206)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i62_1_lut (.A(integrator_d_tmp[61]), .Z(n12_adj_207)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i59_1_lut (.A(integrator_d_tmp[58]), .Z(n15_adj_208)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i60_1_lut (.A(integrator_d_tmp[59]), .Z(n14_adj_209)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i57_1_lut (.A(integrator_d_tmp[56]), .Z(n17_adj_210)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i58_1_lut (.A(integrator_d_tmp[57]), .Z(n16_adj_211)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i55_1_lut (.A(integrator_d_tmp[54]), .Z(n19_adj_212)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i56_1_lut (.A(integrator_d_tmp[55]), .Z(n18_adj_213)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i53_1_lut (.A(integrator_d_tmp[52]), .Z(n21_adj_214)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i54_1_lut (.A(integrator_d_tmp[53]), .Z(n20_adj_215)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i51_1_lut (.A(integrator_d_tmp[50]), .Z(n23_adj_216)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i52_1_lut (.A(integrator_d_tmp[51]), .Z(n22_adj_217)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i49_1_lut (.A(integrator_d_tmp[48]), .Z(n25_adj_218)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i50_1_lut (.A(integrator_d_tmp[49]), .Z(n24_adj_219)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i47_1_lut (.A(integrator_d_tmp[46]), .Z(n27_adj_220)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i47_1_lut.init = 16'h5555;
    FD1S3AX valid_comb_66_rep_374 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_737)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_374.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_373 (.D(clk_80mhz_enable_99), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_38)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=155, LSE_RLINE=161 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_373.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i48_1_lut (.A(integrator_d_tmp[47]), .Z(n26_adj_221)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i45_1_lut (.A(integrator_d_tmp[44]), .Z(n29_adj_222)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i46_1_lut (.A(integrator_d_tmp[45]), .Z(n28_adj_223)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i43_1_lut (.A(integrator_d_tmp[42]), .Z(n31_adj_224)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i43_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module PWM
//

module PWM (\data_in_reg[0] , clk_80mhz, \data_in_reg_11__N_2339[0] , 
            count, \data_in_reg[1] , \data_in_reg_11__N_2339[1] , \data_in_reg[2] , 
            \data_in_reg_11__N_2339[2] , \data_in_reg[3] , \data_in_reg_11__N_2339[3] , 
            \data_in_reg[4] , \data_in_reg_11__N_2339[4] , \data_in_reg[5] , 
            \data_in_reg_11__N_2339[5] , \data_in_reg[6] , \data_in_reg_11__N_2339[6] , 
            \data_in_reg[7] , \data_in_reg_11__N_2339[7] , \data_in_reg[8] , 
            \data_in_reg_11__N_2339[8] , \data_in_reg[9] , GND_net, VCC_net, 
            \amdemod_out[9] ) /* synthesis syn_module_defined=1 */ ;
    output \data_in_reg[0] ;
    input clk_80mhz;
    input \data_in_reg_11__N_2339[0] ;
    output [9:0]count;
    output \data_in_reg[1] ;
    input \data_in_reg_11__N_2339[1] ;
    output \data_in_reg[2] ;
    input \data_in_reg_11__N_2339[2] ;
    output \data_in_reg[3] ;
    input \data_in_reg_11__N_2339[3] ;
    output \data_in_reg[4] ;
    input \data_in_reg_11__N_2339[4] ;
    output \data_in_reg[5] ;
    input \data_in_reg_11__N_2339[5] ;
    output \data_in_reg[6] ;
    input \data_in_reg_11__N_2339[6] ;
    output \data_in_reg[7] ;
    input \data_in_reg_11__N_2339[7] ;
    output \data_in_reg[8] ;
    input \data_in_reg_11__N_2339[8] ;
    output \data_in_reg[9] ;
    input GND_net;
    input VCC_net;
    input \amdemod_out[9] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(64[10:19])
    
    wire clk_80mhz_enable_1443;
    wire [9:0]n45;
    wire [11:0]n2737;
    
    wire n14824, n14823, n14822, n14821, n14820, n11, n12, n17, 
        n15;
    
    FD1P3AX data_in_reg__i1 (.D(\data_in_reg_11__N_2339[0] ), .SP(clk_80mhz_enable_1443), 
            .CK(clk_80mhz), .Q(\data_in_reg[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=198, LSE_RLINE=202 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(43[10] 58[6])
    defparam data_in_reg__i1.GSR = "ENABLED";
    FD1S3AX count_502__i0 (.D(n45[0]), .CK(clk_80mhz), .Q(count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502__i0.GSR = "ENABLED";
    FD1P3AX data_in_reg__i2 (.D(\data_in_reg_11__N_2339[1] ), .SP(clk_80mhz_enable_1443), 
            .CK(clk_80mhz), .Q(\data_in_reg[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=198, LSE_RLINE=202 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(43[10] 58[6])
    defparam data_in_reg__i2.GSR = "ENABLED";
    FD1P3AX data_in_reg__i3 (.D(\data_in_reg_11__N_2339[2] ), .SP(clk_80mhz_enable_1443), 
            .CK(clk_80mhz), .Q(\data_in_reg[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=198, LSE_RLINE=202 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(43[10] 58[6])
    defparam data_in_reg__i3.GSR = "ENABLED";
    FD1P3AX data_in_reg__i4 (.D(\data_in_reg_11__N_2339[3] ), .SP(clk_80mhz_enable_1443), 
            .CK(clk_80mhz), .Q(\data_in_reg[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=198, LSE_RLINE=202 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(43[10] 58[6])
    defparam data_in_reg__i4.GSR = "ENABLED";
    FD1P3AX data_in_reg__i5 (.D(\data_in_reg_11__N_2339[4] ), .SP(clk_80mhz_enable_1443), 
            .CK(clk_80mhz), .Q(\data_in_reg[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=198, LSE_RLINE=202 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(43[10] 58[6])
    defparam data_in_reg__i5.GSR = "ENABLED";
    FD1P3AX data_in_reg__i6 (.D(\data_in_reg_11__N_2339[5] ), .SP(clk_80mhz_enable_1443), 
            .CK(clk_80mhz), .Q(\data_in_reg[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=198, LSE_RLINE=202 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(43[10] 58[6])
    defparam data_in_reg__i6.GSR = "ENABLED";
    FD1P3AX data_in_reg__i7 (.D(\data_in_reg_11__N_2339[6] ), .SP(clk_80mhz_enable_1443), 
            .CK(clk_80mhz), .Q(\data_in_reg[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=198, LSE_RLINE=202 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(43[10] 58[6])
    defparam data_in_reg__i7.GSR = "ENABLED";
    FD1P3AX data_in_reg__i8 (.D(\data_in_reg_11__N_2339[7] ), .SP(clk_80mhz_enable_1443), 
            .CK(clk_80mhz), .Q(\data_in_reg[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=198, LSE_RLINE=202 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(43[10] 58[6])
    defparam data_in_reg__i8.GSR = "ENABLED";
    FD1P3AX data_in_reg__i9 (.D(\data_in_reg_11__N_2339[8] ), .SP(clk_80mhz_enable_1443), 
            .CK(clk_80mhz), .Q(\data_in_reg[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=198, LSE_RLINE=202 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(43[10] 58[6])
    defparam data_in_reg__i9.GSR = "ENABLED";
    FD1P3AX data_in_reg__i10 (.D(n2737[9]), .SP(clk_80mhz_enable_1443), 
            .CK(clk_80mhz), .Q(\data_in_reg[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=198, LSE_RLINE=202 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(43[10] 58[6])
    defparam data_in_reg__i10.GSR = "ENABLED";
    FD1S3AX count_502__i1 (.D(n45[1]), .CK(clk_80mhz), .Q(count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502__i1.GSR = "ENABLED";
    FD1S3AX count_502__i2 (.D(n45[2]), .CK(clk_80mhz), .Q(count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502__i2.GSR = "ENABLED";
    FD1S3AX count_502__i3 (.D(n45[3]), .CK(clk_80mhz), .Q(count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502__i3.GSR = "ENABLED";
    FD1S3AX count_502__i4 (.D(n45[4]), .CK(clk_80mhz), .Q(count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502__i4.GSR = "ENABLED";
    FD1S3AX count_502__i5 (.D(n45[5]), .CK(clk_80mhz), .Q(count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502__i5.GSR = "ENABLED";
    FD1S3AX count_502__i6 (.D(n45[6]), .CK(clk_80mhz), .Q(count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502__i6.GSR = "ENABLED";
    FD1S3AX count_502__i7 (.D(n45[7]), .CK(clk_80mhz), .Q(count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502__i7.GSR = "ENABLED";
    FD1S3AX count_502__i8 (.D(n45[8]), .CK(clk_80mhz), .Q(count[8])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502__i8.GSR = "ENABLED";
    FD1S3AX count_502__i9 (.D(n45[9]), .CK(clk_80mhz), .Q(count[9])) /* synthesis syn_use_carry_chain=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502__i9.GSR = "ENABLED";
    CCU2C count_502_add_4_11 (.A0(count[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n14824), .S0(n45[9]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502_add_4_11.INIT0 = 16'haaa0;
    defparam count_502_add_4_11.INIT1 = 16'h0000;
    defparam count_502_add_4_11.INJECT1_0 = "NO";
    defparam count_502_add_4_11.INJECT1_1 = "NO";
    CCU2C count_502_add_4_9 (.A0(count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14823), .COUT(n14824), .S0(n45[7]), .S1(n45[8]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502_add_4_9.INIT0 = 16'haaa0;
    defparam count_502_add_4_9.INIT1 = 16'haaa0;
    defparam count_502_add_4_9.INJECT1_0 = "NO";
    defparam count_502_add_4_9.INJECT1_1 = "NO";
    CCU2C count_502_add_4_7 (.A0(count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14822), .COUT(n14823), .S0(n45[5]), .S1(n45[6]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502_add_4_7.INIT0 = 16'haaa0;
    defparam count_502_add_4_7.INIT1 = 16'haaa0;
    defparam count_502_add_4_7.INJECT1_0 = "NO";
    defparam count_502_add_4_7.INJECT1_1 = "NO";
    CCU2C count_502_add_4_5 (.A0(count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14821), .COUT(n14822), .S0(n45[3]), .S1(n45[4]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502_add_4_5.INIT0 = 16'haaa0;
    defparam count_502_add_4_5.INIT1 = 16'haaa0;
    defparam count_502_add_4_5.INJECT1_0 = "NO";
    defparam count_502_add_4_5.INJECT1_1 = "NO";
    CCU2C count_502_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(count[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n14820), .COUT(n14821), .S0(n45[1]), .S1(n45[2]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502_add_4_3.INIT0 = 16'haaa0;
    defparam count_502_add_4_3.INIT1 = 16'haaa0;
    defparam count_502_add_4_3.INJECT1_0 = "NO";
    defparam count_502_add_4_3.INJECT1_1 = "NO";
    CCU2C count_502_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n14820), .S1(n45[0]));   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(45[14:26])
    defparam count_502_add_4_1.INIT0 = 16'h0000;
    defparam count_502_add_4_1.INIT1 = 16'h555f;
    defparam count_502_add_4_1.INJECT1_0 = "NO";
    defparam count_502_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(count[0]), .B(count[5]), .Z(n11)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(48[9:19])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2_2_lut (.A(count[8]), .B(count[2]), .Z(n12)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(48[9:19])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i758_1_lut (.A(\amdemod_out[9] ), .Z(n2737[9])) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(48[5] 50[8])
    defparam i758_1_lut.init = 16'h5555;
    LUT4 i5725_4_lut (.A(n17), .B(n15), .C(n11), .D(n12), .Z(clk_80mhz_enable_1443)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(48[9:19])
    defparam i5725_4_lut.init = 16'h0001;
    LUT4 i7_4_lut (.A(count[9]), .B(count[3]), .C(count[7]), .D(count[1]), 
         .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(48[9:19])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(count[6]), .B(count[4]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/PWM.v(48[9:19])
    defparam i5_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module SinCos
//

module SinCos (clk_80mhz, VCC_net, GND_net, \phase_acc[57] , \phase_acc[58] , 
            \phase_acc[59] , \phase_acc[60] , \phase_acc[61] , \phase_acc[62] , 
            \phase_acc[63] , \lo_sinewave[1] , \lo_sinewave[2] , \lo_sinewave[3] , 
            \lo_sinewave[4] , \lo_sinewave[5] , \lo_sinewave[6] , \lo_sinewave[7] , 
            \lo_sinewave[8] , \lo_sinewave[9] , \lo_sinewave[10] , \lo_sinewave[11] , 
            \lo_sinewave[12] , \lo_cosinewave[1] , \lo_cosinewave[2] , 
            \lo_cosinewave[3] , \lo_cosinewave[4] , \lo_cosinewave[5] , 
            \lo_cosinewave[6] , \lo_cosinewave[7] , \lo_cosinewave[8] , 
            \lo_cosinewave[9] , \lo_cosinewave[10] , \lo_cosinewave[11] , 
            \lo_cosinewave[12] , \phase_acc[56] ) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk_80mhz;
    input VCC_net;
    input GND_net;
    input \phase_acc[57] ;
    input \phase_acc[58] ;
    input \phase_acc[59] ;
    input \phase_acc[60] ;
    input \phase_acc[61] ;
    input \phase_acc[62] ;
    input \phase_acc[63] ;
    output \lo_sinewave[1] ;
    output \lo_sinewave[2] ;
    output \lo_sinewave[3] ;
    output \lo_sinewave[4] ;
    output \lo_sinewave[5] ;
    output \lo_sinewave[6] ;
    output \lo_sinewave[7] ;
    output \lo_sinewave[8] ;
    output \lo_sinewave[9] ;
    output \lo_sinewave[10] ;
    output \lo_sinewave[11] ;
    output \lo_sinewave[12] ;
    output \lo_cosinewave[1] ;
    output \lo_cosinewave[2] ;
    output \lo_cosinewave[3] ;
    output \lo_cosinewave[4] ;
    output \lo_cosinewave[5] ;
    output \lo_cosinewave[6] ;
    output \lo_cosinewave[7] ;
    output \lo_cosinewave[8] ;
    output \lo_cosinewave[9] ;
    output \lo_cosinewave[10] ;
    output \lo_cosinewave[11] ;
    output \lo_cosinewave[12] ;
    input \phase_acc[56] ;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(64[10:19])
    
    wire rom_addr0_r_1, rom_addr0_r_1_inv, rom_addr0_r_2, rom_addr0_r_3, 
        rom_addr0_r_4, rom_addr0_r_5, mx_ctrl_r, mx_ctrl_r_1, rom_addr0_r, 
        rom_addr0_r_n, rom_addr0_r_6, rom_dout_11, rom_dout_11_ffin, 
        rom_dout_10, rom_dout_10_ffin, rom_dout_9, rom_dout_9_ffin, 
        rom_dout_8, rom_dout_8_ffin, rom_dout_7, rom_dout_7_ffin, rom_dout_6, 
        rom_dout_6_ffin, rom_dout_5, rom_dout_5_ffin, rom_dout_4, rom_dout_4_ffin, 
        rom_dout_3, rom_dout_3_ffin, rom_dout_2, rom_dout_2_ffin, rom_dout_1, 
        rom_dout_1_ffin, rom_dout, rom_dout_ffin, rom_dout_25, rom_dout_25_ffin, 
        rom_dout_24, rom_dout_24_ffin, rom_dout_23, rom_dout_23_ffin, 
        rom_dout_22, rom_dout_22_ffin, rom_dout_21, rom_dout_21_ffin, 
        rom_dout_20, rom_dout_20_ffin, rom_dout_19, rom_dout_19_ffin, 
        rom_dout_18, rom_dout_18_ffin, rom_dout_17, rom_dout_17_ffin, 
        rom_dout_16, rom_dout_16_ffin, rom_dout_15, rom_dout_15_ffin, 
        rom_dout_14, rom_dout_14_ffin, rom_dout_13, rom_dout_13_ffin, 
        cosromoutsel_i, cosromoutsel, sinromoutsel, sinout_pre_1, sinout_pre_2, 
        sinout_pre_3, sinout_pre_4, sinout_pre_5, sinout_pre_6, sinout_pre_7, 
        sinout_pre_8, sinout_pre_9, sinout_pre_10, sinout_pre_11, sinout_pre_12, 
        cosout_pre_1, cosout_pre_2, cosout_pre_3, cosout_pre_4, cosout_pre_5, 
        cosout_pre_6, cosout_pre_7, cosout_pre_8, cosout_pre_9, cosout_pre_10, 
        cosout_pre_11, cosout_pre_12, rom_addr0_r_inv, co0, rom_addr0_r_n_1, 
        rom_addr0_r_n_2, rom_addr0_r_2_inv, co1, rom_addr0_r_n_3, rom_addr0_r_n_4, 
        rom_addr0_r_4_inv, rom_addr0_r_3_inv, co2, rom_addr0_r_n_5, 
        rom_addr0_r_5_inv, rom_dout_12_ffin, rom_addr0_r_7, rom_addr0_r_8, 
        rom_addr0_r_9, rom_addr0_r_10, rom_addr0_r_11, rom_dout_s_n_1, 
        rom_dout_s_n_2, rom_dout_2_inv, rom_dout_1_inv, co0_1, co1_1, 
        rom_dout_s_n_3, rom_dout_s_n_4, rom_dout_4_inv, rom_dout_3_inv, 
        co2_1, rom_dout_s_n_5, rom_dout_s_n_6, rom_dout_6_inv, rom_dout_5_inv, 
        co3, rom_dout_s_n_7, rom_dout_s_n_8, rom_dout_8_inv, rom_dout_7_inv, 
        co4, rom_dout_s_n_9, rom_dout_s_n_10, rom_dout_10_inv, rom_dout_9_inv, 
        co5, rom_dout_s_n_11, rom_dout_s_n_12, rom_dout_12_inv, rom_dout_11_inv, 
        rom_dout_13_inv, co0_2, rom_dout_c_n_1, rom_dout_c_n_2, rom_dout_15_inv, 
        rom_dout_14_inv, co1_2, rom_dout_c_n_3, rom_dout_c_n_4, rom_dout_17_inv, 
        rom_dout_16_inv, co2_2, rom_dout_c_n_5, rom_dout_c_n_6, rom_dout_19_inv, 
        rom_dout_18_inv, co3_1, rom_dout_c_n_7, rom_dout_c_n_8, rom_dout_21_inv, 
        rom_dout_20_inv, co4_1, rom_dout_c_n_9, rom_dout_c_n_10, rom_dout_23_inv, 
        rom_dout_22_inv, co5_1, rom_dout_c_n_11, rom_dout_c_n_12, rom_dout_25_inv, 
        rom_dout_24_inv, rom_dout_12, rom_dout_inv, func_or_inet, lx_ne0, 
        lx_ne0_inv, out_sel_i, rom_dout_s_1, rom_dout_s_2, rom_dout_s_3, 
        rom_dout_s_4, rom_dout_s_5, rom_dout_s_6, rom_dout_s_7, rom_dout_s_8, 
        rom_dout_s_9, rom_dout_s_10, rom_dout_s_11, rom_dout_s_12, rom_dout_c_1, 
        rom_dout_c_2, rom_dout_c_3, rom_dout_c_4, rom_dout_c_5, rom_dout_c_6, 
        rom_dout_c_7, rom_dout_c_8, rom_dout_c_9, rom_dout_c_10, rom_dout_c_11, 
        rom_dout_c_12, out_sel;
    
    INV INV_29 (.A(rom_addr0_r_1), .Z(rom_addr0_r_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    FD1P3DX FF_61 (.D(\phase_acc[57] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(312[13:88])
    defparam FF_61.GSR = "ENABLED";
    FD1P3DX FF_60 (.D(\phase_acc[58] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(315[13:88])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(\phase_acc[59] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(318[13:88])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(\phase_acc[60] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(321[13:88])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(\phase_acc[61] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(324[13:88])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(\phase_acc[62] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(mx_ctrl_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(327[13:84])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(\phase_acc[63] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(mx_ctrl_r_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(330[13:86])
    defparam FF_55.GSR = "ENABLED";
    MUX21 muxb_57 (.D0(rom_addr0_r), .D1(rom_addr0_r_n), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    FD1P3DX FF_53 (.D(rom_dout_11_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_11)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(355[13] 356[25])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(rom_dout_10_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_10)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(359[13] 360[25])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(rom_dout_9_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_9)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(363[13] 364[24])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(rom_dout_8_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_8)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(367[13] 368[24])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(rom_dout_7_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_7)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(371[13] 372[24])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(rom_dout_6_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_6)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(375[13] 376[24])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(rom_dout_5_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_5)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(379[13] 380[24])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(rom_dout_4_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_4)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(383[13] 384[24])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(rom_dout_3_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_3)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(387[13] 388[24])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(rom_dout_2_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_2)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(391[13] 392[24])
    defparam FF_44.GSR = "ENABLED";
    FD1P3DX FF_43 (.D(rom_dout_1_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_1)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(395[13] 396[24])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(rom_dout_ffin), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(rom_dout)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(399[13] 400[22])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(rom_dout_25_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_25)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(403[13] 404[25])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(rom_dout_24_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_24)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(407[13] 408[25])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(rom_dout_23_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_23)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(411[13] 412[25])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(rom_dout_22_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_22)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(415[13] 416[25])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(rom_dout_21_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_21)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(419[13] 420[25])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(rom_dout_20_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_20)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(423[13] 424[25])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(rom_dout_19_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_19)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(427[13] 428[25])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(rom_dout_18_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_18)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(431[13] 432[25])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(rom_dout_17_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_17)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(435[13] 436[25])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(rom_dout_16_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_16)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(439[13] 440[25])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(rom_dout_15_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_15)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(443[13] 444[25])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(rom_dout_14_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_14)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(447[13] 448[25])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(rom_dout_13_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_13)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(451[13] 452[25])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(cosromoutsel_i), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(cosromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(455[13] 456[26])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(mx_ctrl_r_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(sinromoutsel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(459[13] 460[26])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_24 (.D(sinout_pre_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_sinewave[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(599[13] 600[21])
    defparam FF_24.GSR = "ENABLED";
    FD1P3DX FF_23 (.D(sinout_pre_2), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_sinewave[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(603[13] 604[21])
    defparam FF_23.GSR = "ENABLED";
    FD1P3DX FF_22 (.D(sinout_pre_3), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_sinewave[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(607[13] 608[21])
    defparam FF_22.GSR = "ENABLED";
    FD1P3DX FF_21 (.D(sinout_pre_4), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_sinewave[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(611[13] 612[21])
    defparam FF_21.GSR = "ENABLED";
    FD1P3DX FF_20 (.D(sinout_pre_5), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_sinewave[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(615[13] 616[21])
    defparam FF_20.GSR = "ENABLED";
    FD1P3DX FF_19 (.D(sinout_pre_6), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_sinewave[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(619[13] 620[21])
    defparam FF_19.GSR = "ENABLED";
    FD1P3DX FF_18 (.D(sinout_pre_7), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_sinewave[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(623[13] 624[21])
    defparam FF_18.GSR = "ENABLED";
    FD1P3DX FF_17 (.D(sinout_pre_8), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_sinewave[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(627[13] 628[21])
    defparam FF_17.GSR = "ENABLED";
    FD1P3DX FF_16 (.D(sinout_pre_9), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_sinewave[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(631[13] 632[21])
    defparam FF_16.GSR = "ENABLED";
    FD1P3DX FF_15 (.D(sinout_pre_10), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_sinewave[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(635[13] 636[22])
    defparam FF_15.GSR = "ENABLED";
    FD1P3DX FF_14 (.D(sinout_pre_11), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_sinewave[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(639[13] 640[22])
    defparam FF_14.GSR = "ENABLED";
    FD1P3DX FF_13 (.D(sinout_pre_12), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_sinewave[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(643[13] 644[22])
    defparam FF_13.GSR = "ENABLED";
    FD1P3DX FF_11 (.D(cosout_pre_1), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_cosinewave[1] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(650[13] 651[23])
    defparam FF_11.GSR = "ENABLED";
    FD1P3DX FF_10 (.D(cosout_pre_2), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_cosinewave[2] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(654[13] 655[23])
    defparam FF_10.GSR = "ENABLED";
    FD1P3DX FF_9 (.D(cosout_pre_3), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_cosinewave[3] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(658[13] 659[23])
    defparam FF_9.GSR = "ENABLED";
    FD1P3DX FF_8 (.D(cosout_pre_4), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_cosinewave[4] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(662[13] 663[23])
    defparam FF_8.GSR = "ENABLED";
    FD1P3DX FF_7 (.D(cosout_pre_5), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_cosinewave[5] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(666[13] 667[23])
    defparam FF_7.GSR = "ENABLED";
    FD1P3DX FF_6 (.D(cosout_pre_6), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_cosinewave[6] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(670[13] 671[23])
    defparam FF_6.GSR = "ENABLED";
    FD1P3DX FF_5 (.D(cosout_pre_7), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_cosinewave[7] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(674[13] 675[23])
    defparam FF_5.GSR = "ENABLED";
    FD1P3DX FF_4 (.D(cosout_pre_8), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_cosinewave[8] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(678[13] 679[23])
    defparam FF_4.GSR = "ENABLED";
    FD1P3DX FF_3 (.D(cosout_pre_9), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_cosinewave[9] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(682[13] 683[23])
    defparam FF_3.GSR = "ENABLED";
    FD1P3DX FF_2 (.D(cosout_pre_10), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_cosinewave[10] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(686[13] 687[24])
    defparam FF_2.GSR = "ENABLED";
    FD1P3DX FF_1 (.D(cosout_pre_11), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_cosinewave[11] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(690[13] 691[24])
    defparam FF_1.GSR = "ENABLED";
    FD1P3DX FF_0 (.D(cosout_pre_12), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(\lo_cosinewave[12] )) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(694[13] 695[24])
    defparam FF_0.GSR = "ENABLED";
    CCU2C neg_rom_addr0_r_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0), .S1(rom_addr0_r_n)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(702[11] 704[71])
    defparam neg_rom_addr0_r_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_0.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_0.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_1 (.A0(rom_addr0_r_1_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_2_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0), .COUT(co1), .S0(rom_addr0_r_n_1), 
          .S1(rom_addr0_r_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(710[11] 713[42])
    defparam neg_rom_addr0_r_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_1.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_2 (.A0(rom_addr0_r_3_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_addr0_r_4_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1), .COUT(co2), .S0(rom_addr0_r_n_3), 
          .S1(rom_addr0_r_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(719[11] 722[42])
    defparam neg_rom_addr0_r_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_2.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_addr0_r_n_3 (.A0(rom_addr0_r_5_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co2), .S0(rom_addr0_r_n_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(728[11] 730[73])
    defparam neg_rom_addr0_r_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_addr0_r_n_3.INJECT1_0 = "NO";
    defparam neg_rom_addr0_r_n_3.INJECT1_1 = "NO";
    ROM64X1A triglut_1_0_25 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_12_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_25.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    CCU2C neg_rom_dout_s_n_1 (.A0(rom_dout_1_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_2_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0_1), .COUT(co1_1), .S0(rom_dout_s_n_1), 
          .S1(rom_dout_s_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(874[11] 877[43])
    defparam neg_rom_dout_s_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_1.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_2 (.A0(rom_dout_3_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_4_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1_1), .COUT(co2_1), .S0(rom_dout_s_n_3), 
          .S1(rom_dout_s_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(883[11] 886[43])
    defparam neg_rom_dout_s_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_2.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_3 (.A0(rom_dout_5_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_6_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co2_1), .COUT(co3), .S0(rom_dout_s_n_5), 
          .S1(rom_dout_s_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(892[11] 895[41])
    defparam neg_rom_dout_s_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_3.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_3.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_4 (.A0(rom_dout_7_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_8_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co3), .COUT(co4), .S0(rom_dout_s_n_7), 
          .S1(rom_dout_s_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(901[11] 904[41])
    defparam neg_rom_dout_s_n_4.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_4.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_4.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_4.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_5 (.A0(rom_dout_9_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_10_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co4), .COUT(co5), .S0(rom_dout_s_n_9), 
          .S1(rom_dout_s_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(910[11] 913[42])
    defparam neg_rom_dout_s_n_5.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_5.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_5.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_5.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_s_n_6 (.A0(rom_dout_11_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_12_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co5), .S0(rom_dout_s_n_11), .S1(rom_dout_s_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(919[11] 922[42])
    defparam neg_rom_dout_s_n_6.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_6.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_6.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_6.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_13_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(936[11] 938[72])
    defparam neg_rom_dout_c_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_0.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_0.INJECT1_1 = "NO";
    INV INV_30 (.A(rom_addr0_r_2), .Z(rom_addr0_r_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    CCU2C neg_rom_dout_c_n_1 (.A0(rom_dout_14_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_15_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0_2), .COUT(co1_2), .S0(rom_dout_c_n_1), 
          .S1(rom_dout_c_n_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(944[11] 947[43])
    defparam neg_rom_dout_c_n_1.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_1.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_1.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_1.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_2 (.A0(rom_dout_16_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_17_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co1_2), .COUT(co2_2), .S0(rom_dout_c_n_3), 
          .S1(rom_dout_c_n_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(953[11] 956[43])
    defparam neg_rom_dout_c_n_2.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_2.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_2.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_2.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_3 (.A0(rom_dout_18_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_19_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co2_2), .COUT(co3_1), .S0(rom_dout_c_n_5), 
          .S1(rom_dout_c_n_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(962[11] 965[43])
    defparam neg_rom_dout_c_n_3.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_3.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_3.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_3.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_4 (.A0(rom_dout_20_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_21_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co3_1), .COUT(co4_1), .S0(rom_dout_c_n_7), 
          .S1(rom_dout_c_n_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(971[11] 974[43])
    defparam neg_rom_dout_c_n_4.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_4.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_4.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_4.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_5 (.A0(rom_dout_22_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_23_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co4_1), .COUT(co5_1), .S0(rom_dout_c_n_9), 
          .S1(rom_dout_c_n_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(980[11] 983[44])
    defparam neg_rom_dout_c_n_5.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_5.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_5.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_5.INJECT1_1 = "NO";
    CCU2C neg_rom_dout_c_n_6 (.A0(rom_dout_24_inv), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_25_inv), .B1(GND_net), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co5_1), .S0(rom_dout_c_n_11), .S1(rom_dout_c_n_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(989[11] 992[44])
    defparam neg_rom_dout_c_n_6.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_6.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_c_n_6.INJECT1_0 = "NO";
    defparam neg_rom_dout_c_n_6.INJECT1_1 = "NO";
    INV INV_31 (.A(rom_addr0_r_3), .Z(rom_addr0_r_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_32 (.A(rom_addr0_r_4), .Z(rom_addr0_r_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_33 (.A(rom_addr0_r_5), .Z(rom_addr0_r_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_28 (.A(rom_addr0_r), .Z(rom_addr0_r_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    XOR2 XOR2_t1 (.A(mx_ctrl_r), .B(mx_ctrl_r_1), .Z(cosromoutsel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(241[10:70])
    INV INV_27 (.A(rom_dout_12), .Z(rom_dout_12_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_26 (.A(rom_dout_11), .Z(rom_dout_11_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_25 (.A(rom_dout_10), .Z(rom_dout_10_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_24 (.A(rom_dout_9), .Z(rom_dout_9_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_23 (.A(rom_dout_8), .Z(rom_dout_8_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_22 (.A(rom_dout_7), .Z(rom_dout_7_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_21 (.A(rom_dout_6), .Z(rom_dout_6_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_20 (.A(rom_dout_5), .Z(rom_dout_5_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_19 (.A(rom_dout_4), .Z(rom_dout_4_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_18 (.A(rom_dout_3), .Z(rom_dout_3_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_17 (.A(rom_dout_2), .Z(rom_dout_2_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_16 (.A(rom_dout_1), .Z(rom_dout_1_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_15 (.A(rom_dout), .Z(rom_dout_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_14 (.A(rom_dout_25), .Z(rom_dout_25_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_13 (.A(rom_dout_24), .Z(rom_dout_24_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_12 (.A(rom_dout_23), .Z(rom_dout_23_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_11 (.A(rom_dout_22), .Z(rom_dout_22_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_10 (.A(rom_dout_21), .Z(rom_dout_21_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_9 (.A(rom_dout_20), .Z(rom_dout_20_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_8 (.A(rom_dout_19), .Z(rom_dout_19_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_7 (.A(rom_dout_18), .Z(rom_dout_18_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_6 (.A(rom_dout_17), .Z(rom_dout_17_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_5 (.A(rom_dout_16), .Z(rom_dout_16_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_4 (.A(rom_dout_15), .Z(rom_dout_15_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_3 (.A(rom_dout_14), .Z(rom_dout_14_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    INV INV_2 (.A(rom_dout_13), .Z(rom_dout_13_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    ROM16X1A LUT4_1 (.AD0(rom_addr0_r_9), .AD1(rom_addr0_r_8), .AD2(rom_addr0_r_7), 
            .AD3(rom_addr0_r_6), .DO0(func_or_inet)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam LUT4_1.initval = 16'b1111111111111110;
    ROM16X1A LUT4_0 (.AD0(GND_net), .AD1(rom_addr0_r_11), .AD2(rom_addr0_r_10), 
            .AD3(func_or_inet), .DO0(lx_ne0)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam LUT4_0.initval = 16'b1111111111111110;
    INV INV_1 (.A(lx_ne0), .Z(lx_ne0_inv)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    AND2 AND2_t0 (.A(mx_ctrl_r), .B(lx_ne0_inv), .Z(out_sel_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(305[10:64])
    FD1P3DX FF_62 (.D(\phase_acc[56] ), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_addr0_r)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(309[13:86])
    defparam FF_62.GSR = "ENABLED";
    MUX21 muxb_56 (.D0(rom_addr0_r_1), .D1(rom_addr0_r_n_1), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_55 (.D0(rom_addr0_r_2), .D1(rom_addr0_r_n_2), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_54 (.D0(rom_addr0_r_3), .D1(rom_addr0_r_n_3), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_53 (.D0(rom_addr0_r_4), .D1(rom_addr0_r_n_4), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_52 (.D0(rom_addr0_r_5), .D1(rom_addr0_r_n_5), .SD(mx_ctrl_r), 
          .Z(rom_addr0_r_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    FD1P3DX FF_54 (.D(rom_dout_12_ffin), .SP(VCC_net), .CK(clk_80mhz), 
            .CD(GND_net), .Q(rom_dout_12)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(351[13] 352[25])
    defparam FF_54.GSR = "ENABLED";
    MUX21 muxb_50 (.D0(rom_dout_1), .D1(rom_dout_s_n_1), .SD(sinromoutsel), 
          .Z(rom_dout_s_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_49 (.D0(rom_dout_2), .D1(rom_dout_s_n_2), .SD(sinromoutsel), 
          .Z(rom_dout_s_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_48 (.D0(rom_dout_3), .D1(rom_dout_s_n_3), .SD(sinromoutsel), 
          .Z(rom_dout_s_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_47 (.D0(rom_dout_4), .D1(rom_dout_s_n_4), .SD(sinromoutsel), 
          .Z(rom_dout_s_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_46 (.D0(rom_dout_5), .D1(rom_dout_s_n_5), .SD(sinromoutsel), 
          .Z(rom_dout_s_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_45 (.D0(rom_dout_6), .D1(rom_dout_s_n_6), .SD(sinromoutsel), 
          .Z(rom_dout_s_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_44 (.D0(rom_dout_7), .D1(rom_dout_s_n_7), .SD(sinromoutsel), 
          .Z(rom_dout_s_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_43 (.D0(rom_dout_8), .D1(rom_dout_s_n_8), .SD(sinromoutsel), 
          .Z(rom_dout_s_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_42 (.D0(rom_dout_9), .D1(rom_dout_s_n_9), .SD(sinromoutsel), 
          .Z(rom_dout_s_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_41 (.D0(rom_dout_10), .D1(rom_dout_s_n_10), .SD(sinromoutsel), 
          .Z(rom_dout_s_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_40 (.D0(rom_dout_11), .D1(rom_dout_s_n_11), .SD(sinromoutsel), 
          .Z(rom_dout_s_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_39 (.D0(rom_dout_12), .D1(rom_dout_s_n_12), .SD(sinromoutsel), 
          .Z(rom_dout_s_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_37 (.D0(rom_dout_14), .D1(rom_dout_c_n_1), .SD(cosromoutsel), 
          .Z(rom_dout_c_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_36 (.D0(rom_dout_15), .D1(rom_dout_c_n_2), .SD(cosromoutsel), 
          .Z(rom_dout_c_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_35 (.D0(rom_dout_16), .D1(rom_dout_c_n_3), .SD(cosromoutsel), 
          .Z(rom_dout_c_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_34 (.D0(rom_dout_17), .D1(rom_dout_c_n_4), .SD(cosromoutsel), 
          .Z(rom_dout_c_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_33 (.D0(rom_dout_18), .D1(rom_dout_c_n_5), .SD(cosromoutsel), 
          .Z(rom_dout_c_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_32 (.D0(rom_dout_19), .D1(rom_dout_c_n_6), .SD(cosromoutsel), 
          .Z(rom_dout_c_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_31 (.D0(rom_dout_20), .D1(rom_dout_c_n_7), .SD(cosromoutsel), 
          .Z(rom_dout_c_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_30 (.D0(rom_dout_21), .D1(rom_dout_c_n_8), .SD(cosromoutsel), 
          .Z(rom_dout_c_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_29 (.D0(rom_dout_22), .D1(rom_dout_c_n_9), .SD(cosromoutsel), 
          .Z(rom_dout_c_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_28 (.D0(rom_dout_23), .D1(rom_dout_c_n_10), .SD(cosromoutsel), 
          .Z(rom_dout_c_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_27 (.D0(rom_dout_24), .D1(rom_dout_c_n_11), .SD(cosromoutsel), 
          .Z(rom_dout_c_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_26 (.D0(rom_dout_25), .D1(rom_dout_c_n_12), .SD(cosromoutsel), 
          .Z(rom_dout_c_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    FD1P3DX FF_26 (.D(out_sel_i), .SP(VCC_net), .CK(clk_80mhz), .CD(GND_net), 
            .Q(out_sel)) /* synthesis GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(541[13:83])
    defparam FF_26.GSR = "ENABLED";
    MUX21 muxb_24 (.D0(rom_dout_s_1), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_23 (.D0(rom_dout_s_2), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_22 (.D0(rom_dout_s_3), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_21 (.D0(rom_dout_s_4), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_20 (.D0(rom_dout_s_5), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_19 (.D0(rom_dout_s_6), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_18 (.D0(rom_dout_s_7), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_17 (.D0(rom_dout_s_8), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_16 (.D0(rom_dout_s_9), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_15 (.D0(rom_dout_s_10), .D1(GND_net), .SD(out_sel), .Z(sinout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_14 (.D0(rom_dout_s_11), .D1(VCC_net), .SD(out_sel), .Z(sinout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_13 (.D0(rom_dout_s_12), .D1(mx_ctrl_r_1), .SD(out_sel), 
          .Z(sinout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_11 (.D0(rom_dout_c_1), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_10 (.D0(rom_dout_c_2), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_2)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_9 (.D0(rom_dout_c_3), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_3)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_8 (.D0(rom_dout_c_4), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_4)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_7 (.D0(rom_dout_c_5), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_5)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_6 (.D0(rom_dout_c_6), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_6)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_5 (.D0(rom_dout_c_7), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_7)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_4 (.D0(rom_dout_c_8), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_8)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_3 (.D0(rom_dout_c_9), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_9)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_2 (.D0(rom_dout_c_10), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_10)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_1 (.D0(rom_dout_c_11), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_11)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    MUX21 muxb_0 (.D0(rom_dout_c_12), .D1(GND_net), .SD(out_sel), .Z(cosout_pre_12)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    ROM64X1A triglut_1_0_24 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_11_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_24.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_23 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_10_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_23.initval = 64'b1111111111111111111111111111111111111111110000000000000000000000;
    ROM64X1A triglut_1_0_22 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_9_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_22.initval = 64'b1111111111111111111111111111100000000000001111111111100000000000;
    ROM64X1A triglut_1_0_21 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_8_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_21.initval = 64'b1111111111111111111100000000011111110000001111110000011111000000;
    ROM64X1A triglut_1_0_20 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_7_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_20.initval = 64'b1111111111111100000011111000011110001110001110001110011100111000;
    ROM64X1A triglut_1_0_19 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_6_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_19.initval = 64'b1111111111000011100011100110011001001101101101001001011010110100;
    ROM64X1A triglut_1_0_18 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_5_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_18.initval = 64'b1111111000110011011010010101010100101001001001101100110001100110;
    ROM64X1A triglut_1_0_17 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_4_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_17.initval = 64'b1111100100101010110011000000000001110011011010110101010110101010;
    ROM64X1A triglut_1_0_16 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_3_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_16.initval = 64'b1110010110011100010101001111111101101010110011100000000011110000;
    ROM64X1A triglut_1_0_15 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_2_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_15.initval = 64'b1101000010100011001111010111110011001100010101100000000011001100;
    ROM64X1A triglut_1_0_14 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_1_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_14.initval = 64'b1111011011100010010110111011101001110011000000100111110010101010;
    ROM64X1A triglut_1_0_13 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_13.initval = 64'b1000100101001010011001010111111001010010011110001001001001111000;
    ROM64X1A triglut_1_0_12 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_25_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_12.initval = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    ROM64X1A triglut_1_0_11 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_24_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_11.initval = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    ROM64X1A triglut_1_0_10 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_23_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_10.initval = 64'b0000000000000000000001111111111111111111111111111111111111111110;
    ROM64X1A triglut_1_0_9 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_22_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_9.initval = 64'b0000000000111111111110000000000000111111111111111111111111111110;
    ROM64X1A triglut_1_0_8 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_21_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_8.initval = 64'b0000011111000001111110000001111111000000000111111111111111111110;
    ROM64X1A triglut_1_0_7 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_20_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_7.initval = 64'b0011100111001110001110001110001111000011111000000111111111111110;
    ROM64X1A triglut_1_0_6 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_19_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_6.initval = 64'b0101101011010010010110110110010011001100111000111000011111111110;
    ROM64X1A triglut_1_0_5 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_18_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_5.initval = 64'b1100110001100110110010010010100101010101001011011001100011111110;
    ROM64X1A triglut_1_0_4 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_17_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_4.initval = 64'b1010101101010101101011011001110000000000011001101010100100111110;
    ROM64X1A triglut_1_0_3 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_16_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_3.initval = 64'b0001111000000000111001101010110111111110010101000111001101001110;
    ROM64X1A triglut_1_0_2 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_15_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_2.initval = 64'b0110011000000000110101000110011001111101011110011000101000010110;
    ROM64X1A triglut_1_0_1 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_14_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_1.initval = 64'b1010101001111100100000011001110010111011101101001000111011011110;
    ROM64X1A triglut_1_0_0 (.AD0(rom_addr0_r_6), .AD1(rom_addr0_r_7), .AD2(rom_addr0_r_8), 
            .AD3(rom_addr0_r_9), .AD4(rom_addr0_r_10), .AD5(rom_addr0_r_11), 
            .DO0(rom_dout_13_ffin)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(123[12] 130[6])
    defparam triglut_1_0_0.initval = 64'b0011110010010010001111001001010011111101010011001010010100100010;
    CCU2C neg_rom_dout_s_n_0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), 
          .D0(VCC_net), .A1(rom_dout_inv), .B1(VCC_net), .C1(VCC_net), 
          .D1(VCC_net), .COUT(co0_1)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=123, LSE_RLINE=130 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/SinCos.v(866[11] 868[72])
    defparam neg_rom_dout_s_n_0.INIT0 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_0.INIT1 = 16'b0110011010101010;
    defparam neg_rom_dout_s_n_0.INJECT1_0 = "NO";
    defparam neg_rom_dout_s_n_0.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \CIC(REGISTER_WIDTH=72,DECIMATION_RATIO=4096)_U0 
//

module \CIC(REGISTER_WIDTH=72,DECIMATION_RATIO=4096)_U0  (comb_d6, n21, 
            n20, integrator_tmp, clk_80mhz, integrator5, integrator_d_tmp, 
            integrator2, integrator2_71__N_490, integrator3, integrator3_71__N_562, 
            integrator4, integrator4_71__N_634, integrator5_71__N_706, 
            comb6, comb6_71__N_1451, comb7, comb7_71__N_1523, comb_d7, 
            comb8, comb8_71__N_1595, comb_d8, comb9, comb9_71__N_1667, 
            comb_d9, n23, cic_cosine_out, integrator1, integrator1_71__N_418, 
            n22, n25, n3, n2, n5, n24, n4, n27, n26, n7, 
            n6, n9, n29, n8, n28, n31, n30, n11, count, n67, 
            n33, n10, n13, n12, n15, n32, n14, n17, n16, n19, 
            n18, n35, n21_adj_3, n20_adj_4, n23_adj_5, n34_adj_6, 
            n37_adj_7, n22_adj_8, n36, n25_adj_9, n3_adj_10, n24_adj_11, 
            n27_adj_12, \cic_gain[1] , \comb10[59] , n16607, n2_adj_13, 
            n5_adj_14, n3_adj_15, \comb10[60] , n62, n2_adj_16, n5_adj_17, 
            n26_adj_18, n29_adj_19, n4_adj_20, n28_adj_21, n4_adj_22, 
            n7_adj_23, n7_adj_24, n6_adj_25, n9_adj_26, n8_adj_27, 
            n6_adj_28, n9_adj_29, n8_adj_30, n11_adj_31, n10_adj_32, 
            n13_adj_33, n12_adj_34, n15_adj_35, n14_adj_36, n17_adj_37, 
            n16_adj_38, n19_adj_39, n18_adj_40, n31_adj_41, n21_adj_42, 
            n20_adj_43, n23_adj_44, n22_adj_45, n30_adj_46, n33_adj_47, 
            n32_adj_48, n35_adj_49, n34_adj_50, n37_adj_51, n36_adj_52, 
            n25_adj_53, n3_adj_54, n24_adj_55, n27_adj_56, n2_adj_57, 
            n26_adj_58, n29_adj_59, n5_adj_60, n28_adj_61, n4_adj_62, 
            n7_adj_63, n6_adj_64, n9_adj_65, n8_adj_66, n11_adj_67, 
            n10_adj_68, n13_adj_69, n12_adj_70, n15_adj_71, n14_adj_72, 
            n17_adj_73, n16_adj_74, n19_adj_75, n18_adj_76, n31_adj_77, 
            n11_adj_78, n10_adj_79, n13_adj_80, n12_adj_81, n15_adj_82, 
            n14_adj_83, n30_adj_84, \comb10[61] , \comb10[62] , \comb10[63] , 
            \comb10[64] , \comb10[65] , \comb10[66] , \comb10[67] , 
            \comb10[68] , \comb10[69] , \comb10[70] , \comb10[71] , 
            \data_out_11__N_1811[2] , \data_out_11__N_1811[3] , \data_out_11__N_1811[4] , 
            \data_out_11__N_1811[5] , \data_out_11__N_1811[6] , \data_out_11__N_1811[7] , 
            \data_out_11__N_1811[8] , \data_out_11__N_1811[9] , \data_out_11__N_1811[10] , 
            \data_out_11__N_1811[11] , n33_adj_85, n32_adj_86, n35_adj_87, 
            n34_adj_88, n37_adj_89, n36_adj_90, n118, n120, cout, 
            n115, n117, n112, n114, n109, n111, n106, n108, 
            n103, n105, n100, n102, n97, n99, n94, n96, n91, 
            n93, n88, n90, n85, n87, n82, n84, n79, n81, n76, 
            n78, \cic_gain[0] , n63, n64, n65, n66, n17_adj_91, 
            n16_adj_92, n19_adj_93, n18_adj_94, n21_adj_95, n20_adj_96, 
            n23_adj_97, n22_adj_98, n25_adj_99, n24_adj_100, n27_adj_101, 
            n26_adj_102, n29_adj_103, n28_adj_104, n31_adj_105, n30_adj_106, 
            n33_adj_107, n32_adj_108, n35_adj_109, n34_adj_110, n37_adj_111, 
            n36_adj_112) /* synthesis syn_module_defined=1 */ ;
    output [71:0]comb_d6;
    output n21;
    output n20;
    output [71:0]integrator_tmp;
    input clk_80mhz;
    output [71:0]integrator5;
    output [71:0]integrator_d_tmp;
    output [71:0]integrator2;
    input [71:0]integrator2_71__N_490;
    output [71:0]integrator3;
    input [71:0]integrator3_71__N_562;
    output [71:0]integrator4;
    input [71:0]integrator4_71__N_634;
    input [71:0]integrator5_71__N_706;
    output [71:0]comb6;
    input [71:0]comb6_71__N_1451;
    output [71:0]comb7;
    input [71:0]comb7_71__N_1523;
    output [71:0]comb_d7;
    output [71:0]comb8;
    input [71:0]comb8_71__N_1595;
    output [71:0]comb_d8;
    output [71:0]comb9;
    input [71:0]comb9_71__N_1667;
    output [71:0]comb_d9;
    output n23;
    output [11:0]cic_cosine_out;
    output [71:0]integrator1;
    input [71:0]integrator1_71__N_418;
    output n22;
    output n25;
    output n3;
    output n2;
    output n5;
    output n24;
    output n4;
    output n27;
    output n26;
    output n7;
    output n6;
    output n9;
    output n29;
    output n8;
    output n28;
    output n31;
    output n30;
    output n11;
    output [11:0]count;
    input [11:0]n67;
    output n33;
    output n10;
    output n13;
    output n12;
    output n15;
    output n32;
    output n14;
    output n17;
    output n16;
    output n19;
    output n18;
    output n35;
    output n21_adj_3;
    output n20_adj_4;
    output n23_adj_5;
    output n34_adj_6;
    output n37_adj_7;
    output n22_adj_8;
    output n36;
    output n25_adj_9;
    output n3_adj_10;
    output n24_adj_11;
    output n27_adj_12;
    input \cic_gain[1] ;
    output \comb10[59] ;
    output n16607;
    output n2_adj_13;
    output n5_adj_14;
    output n3_adj_15;
    output \comb10[60] ;
    output n62;
    output n2_adj_16;
    output n5_adj_17;
    output n26_adj_18;
    output n29_adj_19;
    output n4_adj_20;
    output n28_adj_21;
    output n4_adj_22;
    output n7_adj_23;
    output n7_adj_24;
    output n6_adj_25;
    output n9_adj_26;
    output n8_adj_27;
    output n6_adj_28;
    output n9_adj_29;
    output n8_adj_30;
    output n11_adj_31;
    output n10_adj_32;
    output n13_adj_33;
    output n12_adj_34;
    output n15_adj_35;
    output n14_adj_36;
    output n17_adj_37;
    output n16_adj_38;
    output n19_adj_39;
    output n18_adj_40;
    output n31_adj_41;
    output n21_adj_42;
    output n20_adj_43;
    output n23_adj_44;
    output n22_adj_45;
    output n30_adj_46;
    output n33_adj_47;
    output n32_adj_48;
    output n35_adj_49;
    output n34_adj_50;
    output n37_adj_51;
    output n36_adj_52;
    output n25_adj_53;
    output n3_adj_54;
    output n24_adj_55;
    output n27_adj_56;
    output n2_adj_57;
    output n26_adj_58;
    output n29_adj_59;
    output n5_adj_60;
    output n28_adj_61;
    output n4_adj_62;
    output n7_adj_63;
    output n6_adj_64;
    output n9_adj_65;
    output n8_adj_66;
    output n11_adj_67;
    output n10_adj_68;
    output n13_adj_69;
    output n12_adj_70;
    output n15_adj_71;
    output n14_adj_72;
    output n17_adj_73;
    output n16_adj_74;
    output n19_adj_75;
    output n18_adj_76;
    output n31_adj_77;
    output n11_adj_78;
    output n10_adj_79;
    output n13_adj_80;
    output n12_adj_81;
    output n15_adj_82;
    output n14_adj_83;
    output n30_adj_84;
    output \comb10[61] ;
    output \comb10[62] ;
    output \comb10[63] ;
    output \comb10[64] ;
    output \comb10[65] ;
    output \comb10[66] ;
    output \comb10[67] ;
    output \comb10[68] ;
    output \comb10[69] ;
    output \comb10[70] ;
    output \comb10[71] ;
    input \data_out_11__N_1811[2] ;
    input \data_out_11__N_1811[3] ;
    input \data_out_11__N_1811[4] ;
    input \data_out_11__N_1811[5] ;
    input \data_out_11__N_1811[6] ;
    input \data_out_11__N_1811[7] ;
    input \data_out_11__N_1811[8] ;
    input \data_out_11__N_1811[9] ;
    input \data_out_11__N_1811[10] ;
    input \data_out_11__N_1811[11] ;
    output n33_adj_85;
    output n32_adj_86;
    output n35_adj_87;
    output n34_adj_88;
    output n37_adj_89;
    output n36_adj_90;
    input n118;
    input n120;
    input cout;
    input n115;
    input n117;
    input n112;
    input n114;
    input n109;
    input n111;
    input n106;
    input n108;
    input n103;
    input n105;
    input n100;
    input n102;
    input n97;
    input n99;
    input n94;
    input n96;
    input n91;
    input n93;
    input n88;
    input n90;
    input n85;
    input n87;
    input n82;
    input n84;
    input n79;
    input n81;
    input n76;
    input n78;
    input \cic_gain[0] ;
    output n63;
    output n64;
    output n65;
    output n66;
    output n17_adj_91;
    output n16_adj_92;
    output n19_adj_93;
    output n18_adj_94;
    output n21_adj_95;
    output n20_adj_96;
    output n23_adj_97;
    output n22_adj_98;
    output n25_adj_99;
    output n24_adj_100;
    output n27_adj_101;
    output n26_adj_102;
    output n29_adj_103;
    output n28_adj_104;
    output n31_adj_105;
    output n30_adj_106;
    output n33_adj_107;
    output n32_adj_108;
    output n35_adj_109;
    output n34_adj_110;
    output n37_adj_111;
    output n36_adj_112;
    
    wire clk_80mhz /* synthesis SET_AS_NETWORK=clk_80mhz, is_clock=1 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/top.v(64[10:19])
    
    wire clk_80mhz_enable_794, clk_80mhz_enable_834, valid_comb;
    wire [71:0]data_out_11__N_1811;
    
    wire n11961;
    wire [11:0]count_11__N_1438;
    
    wire n23_adj_2474;
    wire [71:0]comb10;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(58[105:111])
    
    wire n17170, n17169, n17210, n17209, count_11__N_1450, clk_80mhz_enable_884, 
        clk_80mhz_enable_934, clk_80mhz_enable_984, clk_80mhz_enable_1034, 
        clk_80mhz_enable_1084, clk_80mhz_enable_1134, clk_80mhz_enable_1184, 
        clk_80mhz_enable_1234, clk_80mhz_enable_1284, clk_80mhz_enable_1334, 
        clk_80mhz_enable_1384, clk_80mhz_enable_1434;
    wire [71:0]comb10_71__N_1739;
    
    wire n16507, n16491, n16503, n16489, n17319, n16545, n16529, 
        n16537, n16541;
    
    LUT4 sub_26_inv_0_i53_1_lut (.A(comb_d6[52]), .Z(n21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i54_1_lut (.A(comb_d6[53]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i54_1_lut.init = 16'h5555;
    FD1P3AX integrator_tmp_i0_i0 (.D(integrator5[0]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i0.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i0 (.D(integrator_tmp[0]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i0.GSR = "ENABLED";
    FD1S3AX integrator2_i0 (.D(integrator2_71__N_490[0]), .CK(clk_80mhz), 
            .Q(integrator2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i0.GSR = "ENABLED";
    FD1S3AX integrator3_i0 (.D(integrator3_71__N_562[0]), .CK(clk_80mhz), 
            .Q(integrator3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i0.GSR = "ENABLED";
    FD1S3AX integrator4_i0 (.D(integrator4_71__N_634[0]), .CK(clk_80mhz), 
            .Q(integrator4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i0.GSR = "ENABLED";
    FD1S3AX integrator5_i0 (.D(integrator5_71__N_706[0]), .CK(clk_80mhz), 
            .Q(integrator5[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i0.GSR = "ENABLED";
    FD1P3AX comb6_i0_i0 (.D(comb6_71__N_1451[0]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(comb6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i0 (.D(comb6[0]), .SP(clk_80mhz_enable_834), .CK(clk_80mhz), 
            .Q(comb_d6[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i0.GSR = "ENABLED";
    FD1S3AX valid_comb_66 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), .Q(valid_comb)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66.GSR = "ENABLED";
    FD1P3AX comb7_i0_i0 (.D(comb7_71__N_1523[0]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(comb7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i0 (.D(comb7[0]), .SP(clk_80mhz_enable_834), .CK(clk_80mhz), 
            .Q(comb_d7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i0.GSR = "ENABLED";
    FD1P3AX comb8_i0_i0 (.D(comb8_71__N_1595[0]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(comb8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i0 (.D(comb8[0]), .SP(clk_80mhz_enable_834), .CK(clk_80mhz), 
            .Q(comb_d8[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i0.GSR = "ENABLED";
    FD1P3AX comb9_i0_i0 (.D(comb9_71__N_1667[0]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(comb9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i0.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i0 (.D(comb9[0]), .SP(clk_80mhz_enable_834), .CK(clk_80mhz), 
            .Q(comb_d9[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i0.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i51_1_lut (.A(comb_d6[50]), .Z(n23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i51_1_lut.init = 16'h5555;
    FD1P3AX data_out_i0_i0 (.D(data_out_11__N_1811[0]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(cic_cosine_out[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i0.GSR = "ENABLED";
    FD1S3AX integrator1_i0 (.D(integrator1_71__N_418[0]), .CK(clk_80mhz), 
            .Q(integrator1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i0.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i52_1_lut (.A(comb_d6[51]), .Z(n22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i49_1_lut (.A(comb_d6[48]), .Z(n25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i71_1_lut (.A(integrator_d_tmp[70]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i72_1_lut (.A(integrator_d_tmp[71]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i69_1_lut (.A(integrator_d_tmp[68]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i50_1_lut (.A(comb_d6[49]), .Z(n24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i70_1_lut (.A(integrator_d_tmp[69]), .Z(n4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i47_1_lut (.A(comb_d6[46]), .Z(n27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i48_1_lut (.A(comb_d6[47]), .Z(n26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i67_1_lut (.A(integrator_d_tmp[66]), .Z(n7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i68_1_lut (.A(integrator_d_tmp[67]), .Z(n6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i65_1_lut (.A(integrator_d_tmp[64]), .Z(n9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i45_1_lut (.A(comb_d6[44]), .Z(n29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i66_1_lut (.A(integrator_d_tmp[65]), .Z(n8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i46_1_lut (.A(comb_d6[45]), .Z(n28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i43_1_lut (.A(comb_d6[42]), .Z(n31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i44_1_lut (.A(comb_d6[43]), .Z(n30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i63_1_lut (.A(integrator_d_tmp[62]), .Z(n11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i63_1_lut.init = 16'h5555;
    FD1S3IX count__i1 (.D(n67[1]), .CK(clk_80mhz), .CD(n11961), .Q(count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i1.GSR = "ENABLED";
    LUT4 sub_26_inv_0_i41_1_lut (.A(comb_d6[40]), .Z(n33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i64_1_lut (.A(integrator_d_tmp[63]), .Z(n10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i61_1_lut (.A(integrator_d_tmp[60]), .Z(n13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i62_1_lut (.A(integrator_d_tmp[61]), .Z(n12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i59_1_lut (.A(integrator_d_tmp[58]), .Z(n15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i42_1_lut (.A(comb_d6[41]), .Z(n32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i60_1_lut (.A(integrator_d_tmp[59]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i57_1_lut (.A(integrator_d_tmp[56]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i58_1_lut (.A(integrator_d_tmp[57]), .Z(n16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i55_1_lut (.A(integrator_d_tmp[54]), .Z(n19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i56_1_lut (.A(integrator_d_tmp[55]), .Z(n18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i39_1_lut (.A(comb_d6[38]), .Z(n35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i53_1_lut (.A(integrator_d_tmp[52]), .Z(n21_adj_3)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i54_1_lut (.A(integrator_d_tmp[53]), .Z(n20_adj_4)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i54_1_lut.init = 16'h5555;
    FD1S3IX count__i0 (.D(count_11__N_1438[0]), .CK(clk_80mhz), .CD(clk_80mhz_enable_794), 
            .Q(count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i0.GSR = "ENABLED";
    LUT4 sub_25_inv_0_i51_1_lut (.A(integrator_d_tmp[50]), .Z(n23_adj_5)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i40_1_lut (.A(comb_d6[39]), .Z(n34_adj_6)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i37_1_lut (.A(comb_d6[36]), .Z(n37_adj_7)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i52_1_lut (.A(integrator_d_tmp[51]), .Z(n22_adj_8)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i38_1_lut (.A(comb_d6[37]), .Z(n36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 i2468_2_lut (.A(n67[11]), .B(n23_adj_2474), .Z(count_11__N_1438[11])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(82[14] 85[8])
    defparam i2468_2_lut.init = 16'hbbbb;
    LUT4 sub_25_inv_0_i49_1_lut (.A(integrator_d_tmp[48]), .Z(n25_adj_9)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i71_1_lut (.A(comb_d7[70]), .Z(n3_adj_10)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i50_1_lut (.A(integrator_d_tmp[49]), .Z(n24_adj_11)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i47_1_lut (.A(integrator_d_tmp[46]), .Z(n27_adj_12)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 i5786_then_3_lut (.A(\cic_gain[1] ), .B(\comb10[59] ), .C(comb10[57]), 
         .Z(n17170)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5786_then_3_lut.init = 16'he4e4;
    LUT4 i5786_else_3_lut (.A(n16607), .B(\cic_gain[1] ), .C(comb10[58]), 
         .Z(n17169)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5786_else_3_lut.init = 16'he2e2;
    LUT4 sub_27_inv_0_i72_1_lut (.A(comb_d7[71]), .Z(n2_adj_13)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i69_1_lut (.A(comb_d7[68]), .Z(n5_adj_14)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 i2389_2_lut (.A(n67[0]), .B(n23_adj_2474), .Z(count_11__N_1438[0])) /* synthesis lut_function=(A+!(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(82[14] 85[8])
    defparam i2389_2_lut.init = 16'hbbbb;
    LUT4 sub_28_inv_0_i71_1_lut (.A(comb_d8[70]), .Z(n3_adj_15)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 i5791_then_3_lut (.A(\cic_gain[1] ), .B(\comb10[60] ), .C(comb10[58]), 
         .Z(n17210)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i5791_then_3_lut.init = 16'he4e4;
    LUT4 i5791_else_3_lut (.A(n62), .B(\cic_gain[1] ), .C(\comb10[59] ), 
         .Z(n17209)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i5791_else_3_lut.init = 16'he2e2;
    LUT4 sub_28_inv_0_i72_1_lut (.A(comb_d8[71]), .Z(n2_adj_16)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i69_1_lut (.A(comb_d8[68]), .Z(n5_adj_17)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i48_1_lut (.A(integrator_d_tmp[47]), .Z(n26_adj_18)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i45_1_lut (.A(integrator_d_tmp[44]), .Z(n29_adj_19)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i70_1_lut (.A(comb_d7[69]), .Z(n4_adj_20)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i46_1_lut (.A(integrator_d_tmp[45]), .Z(n28_adj_21)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i70_1_lut (.A(comb_d8[69]), .Z(n4_adj_22)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i67_1_lut (.A(comb_d7[66]), .Z(n7_adj_23)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i67_1_lut (.A(comb_d8[66]), .Z(n7_adj_24)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i68_1_lut (.A(comb_d8[67]), .Z(n6_adj_25)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i65_1_lut (.A(comb_d8[64]), .Z(n9_adj_26)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i66_1_lut (.A(comb_d8[65]), .Z(n8_adj_27)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i68_1_lut (.A(comb_d7[67]), .Z(n6_adj_28)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i65_1_lut (.A(comb_d7[64]), .Z(n9_adj_29)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i66_1_lut (.A(comb_d7[65]), .Z(n8_adj_30)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i63_1_lut (.A(comb_d7[62]), .Z(n11_adj_31)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i64_1_lut (.A(comb_d7[63]), .Z(n10_adj_32)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i61_1_lut (.A(comb_d7[60]), .Z(n13_adj_33)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i62_1_lut (.A(comb_d7[61]), .Z(n12_adj_34)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i59_1_lut (.A(comb_d7[58]), .Z(n15_adj_35)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i60_1_lut (.A(comb_d7[59]), .Z(n14_adj_36)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i57_1_lut (.A(comb_d7[56]), .Z(n17_adj_37)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i58_1_lut (.A(comb_d7[57]), .Z(n16_adj_38)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i55_1_lut (.A(comb_d7[54]), .Z(n19_adj_39)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i56_1_lut (.A(comb_d7[55]), .Z(n18_adj_40)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i43_1_lut (.A(integrator_d_tmp[42]), .Z(n31_adj_41)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i53_1_lut (.A(comb_d7[52]), .Z(n21_adj_42)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i54_1_lut (.A(comb_d7[53]), .Z(n20_adj_43)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i51_1_lut (.A(comb_d7[50]), .Z(n23_adj_44)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i52_1_lut (.A(comb_d7[51]), .Z(n22_adj_45)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i44_1_lut (.A(integrator_d_tmp[43]), .Z(n30_adj_46)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i41_1_lut (.A(integrator_d_tmp[40]), .Z(n33_adj_47)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i42_1_lut (.A(integrator_d_tmp[41]), .Z(n32_adj_48)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i39_1_lut (.A(integrator_d_tmp[38]), .Z(n35_adj_49)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i40_1_lut (.A(integrator_d_tmp[39]), .Z(n34_adj_50)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i37_1_lut (.A(integrator_d_tmp[36]), .Z(n37_adj_51)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_25_inv_0_i38_1_lut (.A(integrator_d_tmp[37]), .Z(n36_adj_52)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(95[28:61])
    defparam sub_25_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i49_1_lut (.A(comb_d7[48]), .Z(n25_adj_53)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i71_1_lut (.A(comb_d6[70]), .Z(n3_adj_54)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i71_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i50_1_lut (.A(comb_d7[49]), .Z(n24_adj_55)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i47_1_lut (.A(comb_d7[46]), .Z(n27_adj_56)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i72_1_lut (.A(comb_d6[71]), .Z(n2_adj_57)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i72_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i48_1_lut (.A(comb_d7[47]), .Z(n26_adj_58)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i45_1_lut (.A(comb_d7[44]), .Z(n29_adj_59)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i69_1_lut (.A(comb_d6[68]), .Z(n5_adj_60)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i69_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i46_1_lut (.A(comb_d7[45]), .Z(n28_adj_61)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i70_1_lut (.A(comb_d6[69]), .Z(n4_adj_62)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i70_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i67_1_lut (.A(comb_d6[66]), .Z(n7_adj_63)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i67_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i68_1_lut (.A(comb_d6[67]), .Z(n6_adj_64)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i68_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i65_1_lut (.A(comb_d6[64]), .Z(n9_adj_65)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i65_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i66_1_lut (.A(comb_d6[65]), .Z(n8_adj_66)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i66_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i63_1_lut (.A(comb_d6[62]), .Z(n11_adj_67)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i64_1_lut (.A(comb_d6[63]), .Z(n10_adj_68)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i61_1_lut (.A(comb_d6[60]), .Z(n13_adj_69)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i62_1_lut (.A(comb_d6[61]), .Z(n12_adj_70)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i59_1_lut (.A(comb_d6[58]), .Z(n15_adj_71)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i60_1_lut (.A(comb_d6[59]), .Z(n14_adj_72)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i57_1_lut (.A(comb_d6[56]), .Z(n17_adj_73)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i58_1_lut (.A(comb_d6[57]), .Z(n16_adj_74)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i55_1_lut (.A(comb_d6[54]), .Z(n19_adj_75)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_26_inv_0_i56_1_lut (.A(comb_d6[55]), .Z(n18_adj_76)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(97[28:43])
    defparam sub_26_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i43_1_lut (.A(comb_d7[42]), .Z(n31_adj_77)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i63_1_lut (.A(comb_d8[62]), .Z(n11_adj_78)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i63_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i64_1_lut (.A(comb_d8[63]), .Z(n10_adj_79)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i64_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i61_1_lut (.A(comb_d8[60]), .Z(n13_adj_80)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i61_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i62_1_lut (.A(comb_d8[61]), .Z(n12_adj_81)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i62_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i59_1_lut (.A(comb_d8[58]), .Z(n15_adj_82)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i59_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i60_1_lut (.A(comb_d8[59]), .Z(n14_adj_83)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i60_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i44_1_lut (.A(comb_d7[43]), .Z(n30_adj_84)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i44_1_lut.init = 16'h5555;
    FD1P3AX integrator_tmp_i0_i1 (.D(integrator5[1]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i2 (.D(integrator5[2]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i3 (.D(integrator5[3]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i4 (.D(integrator5[4]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i5 (.D(integrator5[5]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i6 (.D(integrator5[6]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i7 (.D(integrator5[7]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i8 (.D(integrator5[8]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i9 (.D(integrator5[9]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i10 (.D(integrator5[10]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i11 (.D(integrator5[11]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i12 (.D(integrator5[12]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i13 (.D(integrator5[13]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i14 (.D(integrator5[14]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i15 (.D(integrator5[15]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i16 (.D(integrator5[16]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i17 (.D(integrator5[17]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i18 (.D(integrator5[18]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i19 (.D(integrator5[19]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i20 (.D(integrator5[20]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i21 (.D(integrator5[21]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i22 (.D(integrator5[22]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i23 (.D(integrator5[23]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i24 (.D(integrator5[24]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i25 (.D(integrator5[25]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i26 (.D(integrator5[26]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i27 (.D(integrator5[27]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i28 (.D(integrator5[28]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i29 (.D(integrator5[29]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i30 (.D(integrator5[30]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i31 (.D(integrator5[31]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i32 (.D(integrator5[32]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i33 (.D(integrator5[33]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i34 (.D(integrator5[34]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i35 (.D(integrator5[35]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i36 (.D(integrator5[36]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i37 (.D(integrator5[37]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i38 (.D(integrator5[38]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i39 (.D(integrator5[39]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i40 (.D(integrator5[40]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i41 (.D(integrator5[41]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i42 (.D(integrator5[42]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i43 (.D(integrator5[43]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i44 (.D(integrator5[44]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i45 (.D(integrator5[45]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i46 (.D(integrator5[46]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i47 (.D(integrator5[47]), .SP(clk_80mhz_enable_794), 
            .CK(clk_80mhz), .Q(integrator_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i48 (.D(integrator5[48]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i49 (.D(integrator5[49]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i50 (.D(integrator5[50]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i51 (.D(integrator5[51]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i52 (.D(integrator5[52]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i53 (.D(integrator5[53]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i54 (.D(integrator5[54]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i55 (.D(integrator5[55]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i56 (.D(integrator5[56]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i57 (.D(integrator5[57]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i58 (.D(integrator5[58]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i59 (.D(integrator5[59]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i60 (.D(integrator5[60]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i61 (.D(integrator5[61]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i62 (.D(integrator5[62]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i63 (.D(integrator5[63]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i64 (.D(integrator5[64]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i65 (.D(integrator5[65]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i66 (.D(integrator5[66]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i67 (.D(integrator5[67]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i68 (.D(integrator5[68]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i69 (.D(integrator5[69]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i70 (.D(integrator5[70]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX integrator_tmp_i0_i71 (.D(integrator5[71]), .SP(count_11__N_1450), 
            .CK(clk_80mhz), .Q(integrator_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator_tmp_i0_i71.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i1 (.D(integrator_tmp[1]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i1.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i2 (.D(integrator_tmp[2]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i2.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i3 (.D(integrator_tmp[3]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i3.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i4 (.D(integrator_tmp[4]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i4.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i5 (.D(integrator_tmp[5]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i5.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i6 (.D(integrator_tmp[6]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i6.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i7 (.D(integrator_tmp[7]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i7.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i8 (.D(integrator_tmp[8]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i8.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i9 (.D(integrator_tmp[9]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i9.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i10 (.D(integrator_tmp[10]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i10.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i11 (.D(integrator_tmp[11]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i11.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i12 (.D(integrator_tmp[12]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i12.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i13 (.D(integrator_tmp[13]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i13.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i14 (.D(integrator_tmp[14]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i14.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i15 (.D(integrator_tmp[15]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i15.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i16 (.D(integrator_tmp[16]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i16.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i17 (.D(integrator_tmp[17]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i17.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i18 (.D(integrator_tmp[18]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i18.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i19 (.D(integrator_tmp[19]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i19.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i20 (.D(integrator_tmp[20]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i20.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i21 (.D(integrator_tmp[21]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i21.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i22 (.D(integrator_tmp[22]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i22.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i23 (.D(integrator_tmp[23]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i23.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i24 (.D(integrator_tmp[24]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i24.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i25 (.D(integrator_tmp[25]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i25.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i26 (.D(integrator_tmp[26]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i26.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i27 (.D(integrator_tmp[27]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i27.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i28 (.D(integrator_tmp[28]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i28.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i29 (.D(integrator_tmp[29]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i29.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i30 (.D(integrator_tmp[30]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i30.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i31 (.D(integrator_tmp[31]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i31.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i32 (.D(integrator_tmp[32]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i32.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i33 (.D(integrator_tmp[33]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i33.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i34 (.D(integrator_tmp[34]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i34.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i35 (.D(integrator_tmp[35]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i35.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i36 (.D(integrator_tmp[36]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i36.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i37 (.D(integrator_tmp[37]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i37.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i38 (.D(integrator_tmp[38]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i38.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i39 (.D(integrator_tmp[39]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i39.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i40 (.D(integrator_tmp[40]), .SP(clk_80mhz_enable_834), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i40.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i41 (.D(integrator_tmp[41]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i41.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i42 (.D(integrator_tmp[42]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i42.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i43 (.D(integrator_tmp[43]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i43.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i44 (.D(integrator_tmp[44]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i44.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i45 (.D(integrator_tmp[45]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i45.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i46 (.D(integrator_tmp[46]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i46.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i47 (.D(integrator_tmp[47]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i47.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i48 (.D(integrator_tmp[48]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i48.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i49 (.D(integrator_tmp[49]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i49.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i50 (.D(integrator_tmp[50]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i50.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i51 (.D(integrator_tmp[51]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i51.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i52 (.D(integrator_tmp[52]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i52.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i53 (.D(integrator_tmp[53]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i53.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i54 (.D(integrator_tmp[54]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i54.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i55 (.D(integrator_tmp[55]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i55.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i56 (.D(integrator_tmp[56]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i56.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i57 (.D(integrator_tmp[57]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i57.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i58 (.D(integrator_tmp[58]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i58.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i59 (.D(integrator_tmp[59]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i59.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i60 (.D(integrator_tmp[60]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i60.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i61 (.D(integrator_tmp[61]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i61.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i62 (.D(integrator_tmp[62]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i62.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i63 (.D(integrator_tmp[63]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i63.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i64 (.D(integrator_tmp[64]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i64.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i65 (.D(integrator_tmp[65]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i65.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i66 (.D(integrator_tmp[66]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i66.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i67 (.D(integrator_tmp[67]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i67.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i68 (.D(integrator_tmp[68]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i68.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i69 (.D(integrator_tmp[69]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i69.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i70 (.D(integrator_tmp[70]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i70.GSR = "ENABLED";
    FD1P3AX integrator_d_tmp_i0_i71 (.D(integrator_tmp[71]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(integrator_d_tmp[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam integrator_d_tmp_i0_i71.GSR = "ENABLED";
    FD1S3AX integrator2_i1 (.D(integrator2_71__N_490[1]), .CK(clk_80mhz), 
            .Q(integrator2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i1.GSR = "ENABLED";
    FD1S3AX integrator2_i2 (.D(integrator2_71__N_490[2]), .CK(clk_80mhz), 
            .Q(integrator2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i2.GSR = "ENABLED";
    FD1S3AX integrator2_i3 (.D(integrator2_71__N_490[3]), .CK(clk_80mhz), 
            .Q(integrator2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i3.GSR = "ENABLED";
    FD1S3AX integrator2_i4 (.D(integrator2_71__N_490[4]), .CK(clk_80mhz), 
            .Q(integrator2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i4.GSR = "ENABLED";
    FD1S3AX integrator2_i5 (.D(integrator2_71__N_490[5]), .CK(clk_80mhz), 
            .Q(integrator2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i5.GSR = "ENABLED";
    FD1S3AX integrator2_i6 (.D(integrator2_71__N_490[6]), .CK(clk_80mhz), 
            .Q(integrator2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i6.GSR = "ENABLED";
    FD1S3AX integrator2_i7 (.D(integrator2_71__N_490[7]), .CK(clk_80mhz), 
            .Q(integrator2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i7.GSR = "ENABLED";
    FD1S3AX integrator2_i8 (.D(integrator2_71__N_490[8]), .CK(clk_80mhz), 
            .Q(integrator2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i8.GSR = "ENABLED";
    FD1S3AX integrator2_i9 (.D(integrator2_71__N_490[9]), .CK(clk_80mhz), 
            .Q(integrator2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i9.GSR = "ENABLED";
    FD1S3AX integrator2_i10 (.D(integrator2_71__N_490[10]), .CK(clk_80mhz), 
            .Q(integrator2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i10.GSR = "ENABLED";
    FD1S3AX integrator2_i11 (.D(integrator2_71__N_490[11]), .CK(clk_80mhz), 
            .Q(integrator2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i11.GSR = "ENABLED";
    FD1S3AX integrator2_i12 (.D(integrator2_71__N_490[12]), .CK(clk_80mhz), 
            .Q(integrator2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i12.GSR = "ENABLED";
    FD1S3AX integrator2_i13 (.D(integrator2_71__N_490[13]), .CK(clk_80mhz), 
            .Q(integrator2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i13.GSR = "ENABLED";
    FD1S3AX integrator2_i14 (.D(integrator2_71__N_490[14]), .CK(clk_80mhz), 
            .Q(integrator2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i14.GSR = "ENABLED";
    FD1S3AX integrator2_i15 (.D(integrator2_71__N_490[15]), .CK(clk_80mhz), 
            .Q(integrator2[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i15.GSR = "ENABLED";
    FD1S3AX integrator2_i16 (.D(integrator2_71__N_490[16]), .CK(clk_80mhz), 
            .Q(integrator2[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i16.GSR = "ENABLED";
    FD1S3AX integrator2_i17 (.D(integrator2_71__N_490[17]), .CK(clk_80mhz), 
            .Q(integrator2[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i17.GSR = "ENABLED";
    FD1S3AX integrator2_i18 (.D(integrator2_71__N_490[18]), .CK(clk_80mhz), 
            .Q(integrator2[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i18.GSR = "ENABLED";
    FD1S3AX integrator2_i19 (.D(integrator2_71__N_490[19]), .CK(clk_80mhz), 
            .Q(integrator2[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i19.GSR = "ENABLED";
    FD1S3AX integrator2_i20 (.D(integrator2_71__N_490[20]), .CK(clk_80mhz), 
            .Q(integrator2[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i20.GSR = "ENABLED";
    FD1S3AX integrator2_i21 (.D(integrator2_71__N_490[21]), .CK(clk_80mhz), 
            .Q(integrator2[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i21.GSR = "ENABLED";
    FD1S3AX integrator2_i22 (.D(integrator2_71__N_490[22]), .CK(clk_80mhz), 
            .Q(integrator2[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i22.GSR = "ENABLED";
    FD1S3AX integrator2_i23 (.D(integrator2_71__N_490[23]), .CK(clk_80mhz), 
            .Q(integrator2[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i23.GSR = "ENABLED";
    FD1S3AX integrator2_i24 (.D(integrator2_71__N_490[24]), .CK(clk_80mhz), 
            .Q(integrator2[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i24.GSR = "ENABLED";
    FD1S3AX integrator2_i25 (.D(integrator2_71__N_490[25]), .CK(clk_80mhz), 
            .Q(integrator2[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i25.GSR = "ENABLED";
    FD1S3AX integrator2_i26 (.D(integrator2_71__N_490[26]), .CK(clk_80mhz), 
            .Q(integrator2[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i26.GSR = "ENABLED";
    FD1S3AX integrator2_i27 (.D(integrator2_71__N_490[27]), .CK(clk_80mhz), 
            .Q(integrator2[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i27.GSR = "ENABLED";
    FD1S3AX integrator2_i28 (.D(integrator2_71__N_490[28]), .CK(clk_80mhz), 
            .Q(integrator2[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i28.GSR = "ENABLED";
    FD1S3AX integrator2_i29 (.D(integrator2_71__N_490[29]), .CK(clk_80mhz), 
            .Q(integrator2[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i29.GSR = "ENABLED";
    FD1S3AX integrator2_i30 (.D(integrator2_71__N_490[30]), .CK(clk_80mhz), 
            .Q(integrator2[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i30.GSR = "ENABLED";
    FD1S3AX integrator2_i31 (.D(integrator2_71__N_490[31]), .CK(clk_80mhz), 
            .Q(integrator2[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i31.GSR = "ENABLED";
    FD1S3AX integrator2_i32 (.D(integrator2_71__N_490[32]), .CK(clk_80mhz), 
            .Q(integrator2[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i32.GSR = "ENABLED";
    FD1S3AX integrator2_i33 (.D(integrator2_71__N_490[33]), .CK(clk_80mhz), 
            .Q(integrator2[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i33.GSR = "ENABLED";
    FD1S3AX integrator2_i34 (.D(integrator2_71__N_490[34]), .CK(clk_80mhz), 
            .Q(integrator2[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i34.GSR = "ENABLED";
    FD1S3AX integrator2_i35 (.D(integrator2_71__N_490[35]), .CK(clk_80mhz), 
            .Q(integrator2[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i35.GSR = "ENABLED";
    FD1S3AX integrator2_i36 (.D(integrator2_71__N_490[36]), .CK(clk_80mhz), 
            .Q(integrator2[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i36.GSR = "ENABLED";
    FD1S3AX integrator2_i37 (.D(integrator2_71__N_490[37]), .CK(clk_80mhz), 
            .Q(integrator2[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i37.GSR = "ENABLED";
    FD1S3AX integrator2_i38 (.D(integrator2_71__N_490[38]), .CK(clk_80mhz), 
            .Q(integrator2[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i38.GSR = "ENABLED";
    FD1S3AX integrator2_i39 (.D(integrator2_71__N_490[39]), .CK(clk_80mhz), 
            .Q(integrator2[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i39.GSR = "ENABLED";
    FD1S3AX integrator2_i40 (.D(integrator2_71__N_490[40]), .CK(clk_80mhz), 
            .Q(integrator2[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i40.GSR = "ENABLED";
    FD1S3AX integrator2_i41 (.D(integrator2_71__N_490[41]), .CK(clk_80mhz), 
            .Q(integrator2[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i41.GSR = "ENABLED";
    FD1S3AX integrator2_i42 (.D(integrator2_71__N_490[42]), .CK(clk_80mhz), 
            .Q(integrator2[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i42.GSR = "ENABLED";
    FD1S3AX integrator2_i43 (.D(integrator2_71__N_490[43]), .CK(clk_80mhz), 
            .Q(integrator2[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i43.GSR = "ENABLED";
    FD1S3AX integrator2_i44 (.D(integrator2_71__N_490[44]), .CK(clk_80mhz), 
            .Q(integrator2[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i44.GSR = "ENABLED";
    FD1S3AX integrator2_i45 (.D(integrator2_71__N_490[45]), .CK(clk_80mhz), 
            .Q(integrator2[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i45.GSR = "ENABLED";
    FD1S3AX integrator2_i46 (.D(integrator2_71__N_490[46]), .CK(clk_80mhz), 
            .Q(integrator2[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i46.GSR = "ENABLED";
    FD1S3AX integrator2_i47 (.D(integrator2_71__N_490[47]), .CK(clk_80mhz), 
            .Q(integrator2[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i47.GSR = "ENABLED";
    FD1S3AX integrator2_i48 (.D(integrator2_71__N_490[48]), .CK(clk_80mhz), 
            .Q(integrator2[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i48.GSR = "ENABLED";
    FD1S3AX integrator2_i49 (.D(integrator2_71__N_490[49]), .CK(clk_80mhz), 
            .Q(integrator2[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i49.GSR = "ENABLED";
    FD1S3AX integrator2_i50 (.D(integrator2_71__N_490[50]), .CK(clk_80mhz), 
            .Q(integrator2[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i50.GSR = "ENABLED";
    FD1S3AX integrator2_i51 (.D(integrator2_71__N_490[51]), .CK(clk_80mhz), 
            .Q(integrator2[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i51.GSR = "ENABLED";
    FD1S3AX integrator2_i52 (.D(integrator2_71__N_490[52]), .CK(clk_80mhz), 
            .Q(integrator2[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i52.GSR = "ENABLED";
    FD1S3AX integrator2_i53 (.D(integrator2_71__N_490[53]), .CK(clk_80mhz), 
            .Q(integrator2[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i53.GSR = "ENABLED";
    FD1S3AX integrator2_i54 (.D(integrator2_71__N_490[54]), .CK(clk_80mhz), 
            .Q(integrator2[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i54.GSR = "ENABLED";
    FD1S3AX integrator2_i55 (.D(integrator2_71__N_490[55]), .CK(clk_80mhz), 
            .Q(integrator2[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i55.GSR = "ENABLED";
    FD1S3AX integrator2_i56 (.D(integrator2_71__N_490[56]), .CK(clk_80mhz), 
            .Q(integrator2[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i56.GSR = "ENABLED";
    FD1S3AX integrator2_i57 (.D(integrator2_71__N_490[57]), .CK(clk_80mhz), 
            .Q(integrator2[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i57.GSR = "ENABLED";
    FD1S3AX integrator2_i58 (.D(integrator2_71__N_490[58]), .CK(clk_80mhz), 
            .Q(integrator2[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i58.GSR = "ENABLED";
    FD1S3AX integrator2_i59 (.D(integrator2_71__N_490[59]), .CK(clk_80mhz), 
            .Q(integrator2[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i59.GSR = "ENABLED";
    FD1S3AX integrator2_i60 (.D(integrator2_71__N_490[60]), .CK(clk_80mhz), 
            .Q(integrator2[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i60.GSR = "ENABLED";
    FD1S3AX integrator2_i61 (.D(integrator2_71__N_490[61]), .CK(clk_80mhz), 
            .Q(integrator2[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i61.GSR = "ENABLED";
    FD1S3AX integrator2_i62 (.D(integrator2_71__N_490[62]), .CK(clk_80mhz), 
            .Q(integrator2[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i62.GSR = "ENABLED";
    FD1S3AX integrator2_i63 (.D(integrator2_71__N_490[63]), .CK(clk_80mhz), 
            .Q(integrator2[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i63.GSR = "ENABLED";
    FD1S3AX integrator2_i64 (.D(integrator2_71__N_490[64]), .CK(clk_80mhz), 
            .Q(integrator2[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i64.GSR = "ENABLED";
    FD1S3AX integrator2_i65 (.D(integrator2_71__N_490[65]), .CK(clk_80mhz), 
            .Q(integrator2[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i65.GSR = "ENABLED";
    FD1S3AX integrator2_i66 (.D(integrator2_71__N_490[66]), .CK(clk_80mhz), 
            .Q(integrator2[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i66.GSR = "ENABLED";
    FD1S3AX integrator2_i67 (.D(integrator2_71__N_490[67]), .CK(clk_80mhz), 
            .Q(integrator2[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i67.GSR = "ENABLED";
    FD1S3AX integrator2_i68 (.D(integrator2_71__N_490[68]), .CK(clk_80mhz), 
            .Q(integrator2[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i68.GSR = "ENABLED";
    FD1S3AX integrator2_i69 (.D(integrator2_71__N_490[69]), .CK(clk_80mhz), 
            .Q(integrator2[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i69.GSR = "ENABLED";
    FD1S3AX integrator2_i70 (.D(integrator2_71__N_490[70]), .CK(clk_80mhz), 
            .Q(integrator2[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i70.GSR = "ENABLED";
    FD1S3AX integrator2_i71 (.D(integrator2_71__N_490[71]), .CK(clk_80mhz), 
            .Q(integrator2[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator2_i71.GSR = "ENABLED";
    FD1S3AX integrator3_i1 (.D(integrator3_71__N_562[1]), .CK(clk_80mhz), 
            .Q(integrator3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i1.GSR = "ENABLED";
    FD1S3AX integrator3_i2 (.D(integrator3_71__N_562[2]), .CK(clk_80mhz), 
            .Q(integrator3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i2.GSR = "ENABLED";
    FD1S3AX integrator3_i3 (.D(integrator3_71__N_562[3]), .CK(clk_80mhz), 
            .Q(integrator3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i3.GSR = "ENABLED";
    FD1S3AX integrator3_i4 (.D(integrator3_71__N_562[4]), .CK(clk_80mhz), 
            .Q(integrator3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i4.GSR = "ENABLED";
    FD1S3AX integrator3_i5 (.D(integrator3_71__N_562[5]), .CK(clk_80mhz), 
            .Q(integrator3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i5.GSR = "ENABLED";
    FD1S3AX integrator3_i6 (.D(integrator3_71__N_562[6]), .CK(clk_80mhz), 
            .Q(integrator3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i6.GSR = "ENABLED";
    FD1S3AX integrator3_i7 (.D(integrator3_71__N_562[7]), .CK(clk_80mhz), 
            .Q(integrator3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i7.GSR = "ENABLED";
    FD1S3AX integrator3_i8 (.D(integrator3_71__N_562[8]), .CK(clk_80mhz), 
            .Q(integrator3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i8.GSR = "ENABLED";
    FD1S3AX integrator3_i9 (.D(integrator3_71__N_562[9]), .CK(clk_80mhz), 
            .Q(integrator3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i9.GSR = "ENABLED";
    FD1S3AX integrator3_i10 (.D(integrator3_71__N_562[10]), .CK(clk_80mhz), 
            .Q(integrator3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i10.GSR = "ENABLED";
    FD1S3AX integrator3_i11 (.D(integrator3_71__N_562[11]), .CK(clk_80mhz), 
            .Q(integrator3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i11.GSR = "ENABLED";
    FD1S3AX integrator3_i12 (.D(integrator3_71__N_562[12]), .CK(clk_80mhz), 
            .Q(integrator3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i12.GSR = "ENABLED";
    FD1S3AX integrator3_i13 (.D(integrator3_71__N_562[13]), .CK(clk_80mhz), 
            .Q(integrator3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i13.GSR = "ENABLED";
    FD1S3AX integrator3_i14 (.D(integrator3_71__N_562[14]), .CK(clk_80mhz), 
            .Q(integrator3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i14.GSR = "ENABLED";
    FD1S3AX integrator3_i15 (.D(integrator3_71__N_562[15]), .CK(clk_80mhz), 
            .Q(integrator3[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i15.GSR = "ENABLED";
    FD1S3AX integrator3_i16 (.D(integrator3_71__N_562[16]), .CK(clk_80mhz), 
            .Q(integrator3[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i16.GSR = "ENABLED";
    FD1S3AX integrator3_i17 (.D(integrator3_71__N_562[17]), .CK(clk_80mhz), 
            .Q(integrator3[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i17.GSR = "ENABLED";
    FD1S3AX integrator3_i18 (.D(integrator3_71__N_562[18]), .CK(clk_80mhz), 
            .Q(integrator3[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i18.GSR = "ENABLED";
    FD1S3AX integrator3_i19 (.D(integrator3_71__N_562[19]), .CK(clk_80mhz), 
            .Q(integrator3[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i19.GSR = "ENABLED";
    FD1S3AX integrator3_i20 (.D(integrator3_71__N_562[20]), .CK(clk_80mhz), 
            .Q(integrator3[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i20.GSR = "ENABLED";
    FD1S3AX integrator3_i21 (.D(integrator3_71__N_562[21]), .CK(clk_80mhz), 
            .Q(integrator3[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i21.GSR = "ENABLED";
    FD1S3AX integrator3_i22 (.D(integrator3_71__N_562[22]), .CK(clk_80mhz), 
            .Q(integrator3[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i22.GSR = "ENABLED";
    FD1S3AX integrator3_i23 (.D(integrator3_71__N_562[23]), .CK(clk_80mhz), 
            .Q(integrator3[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i23.GSR = "ENABLED";
    FD1S3AX integrator3_i24 (.D(integrator3_71__N_562[24]), .CK(clk_80mhz), 
            .Q(integrator3[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i24.GSR = "ENABLED";
    FD1S3AX integrator3_i25 (.D(integrator3_71__N_562[25]), .CK(clk_80mhz), 
            .Q(integrator3[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i25.GSR = "ENABLED";
    FD1S3AX integrator3_i26 (.D(integrator3_71__N_562[26]), .CK(clk_80mhz), 
            .Q(integrator3[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i26.GSR = "ENABLED";
    FD1S3AX integrator3_i27 (.D(integrator3_71__N_562[27]), .CK(clk_80mhz), 
            .Q(integrator3[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i27.GSR = "ENABLED";
    FD1S3AX integrator3_i28 (.D(integrator3_71__N_562[28]), .CK(clk_80mhz), 
            .Q(integrator3[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i28.GSR = "ENABLED";
    FD1S3AX integrator3_i29 (.D(integrator3_71__N_562[29]), .CK(clk_80mhz), 
            .Q(integrator3[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i29.GSR = "ENABLED";
    FD1S3AX integrator3_i30 (.D(integrator3_71__N_562[30]), .CK(clk_80mhz), 
            .Q(integrator3[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i30.GSR = "ENABLED";
    FD1S3AX integrator3_i31 (.D(integrator3_71__N_562[31]), .CK(clk_80mhz), 
            .Q(integrator3[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i31.GSR = "ENABLED";
    FD1S3AX integrator3_i32 (.D(integrator3_71__N_562[32]), .CK(clk_80mhz), 
            .Q(integrator3[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i32.GSR = "ENABLED";
    FD1S3AX integrator3_i33 (.D(integrator3_71__N_562[33]), .CK(clk_80mhz), 
            .Q(integrator3[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i33.GSR = "ENABLED";
    FD1S3AX integrator3_i34 (.D(integrator3_71__N_562[34]), .CK(clk_80mhz), 
            .Q(integrator3[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i34.GSR = "ENABLED";
    FD1S3AX integrator3_i35 (.D(integrator3_71__N_562[35]), .CK(clk_80mhz), 
            .Q(integrator3[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i35.GSR = "ENABLED";
    FD1S3AX integrator3_i36 (.D(integrator3_71__N_562[36]), .CK(clk_80mhz), 
            .Q(integrator3[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i36.GSR = "ENABLED";
    FD1S3AX integrator3_i37 (.D(integrator3_71__N_562[37]), .CK(clk_80mhz), 
            .Q(integrator3[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i37.GSR = "ENABLED";
    FD1S3AX integrator3_i38 (.D(integrator3_71__N_562[38]), .CK(clk_80mhz), 
            .Q(integrator3[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i38.GSR = "ENABLED";
    FD1S3AX integrator3_i39 (.D(integrator3_71__N_562[39]), .CK(clk_80mhz), 
            .Q(integrator3[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i39.GSR = "ENABLED";
    FD1S3AX integrator3_i40 (.D(integrator3_71__N_562[40]), .CK(clk_80mhz), 
            .Q(integrator3[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i40.GSR = "ENABLED";
    FD1S3AX integrator3_i41 (.D(integrator3_71__N_562[41]), .CK(clk_80mhz), 
            .Q(integrator3[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i41.GSR = "ENABLED";
    FD1S3AX integrator3_i42 (.D(integrator3_71__N_562[42]), .CK(clk_80mhz), 
            .Q(integrator3[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i42.GSR = "ENABLED";
    FD1S3AX integrator3_i43 (.D(integrator3_71__N_562[43]), .CK(clk_80mhz), 
            .Q(integrator3[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i43.GSR = "ENABLED";
    FD1S3AX integrator3_i44 (.D(integrator3_71__N_562[44]), .CK(clk_80mhz), 
            .Q(integrator3[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i44.GSR = "ENABLED";
    FD1S3AX integrator3_i45 (.D(integrator3_71__N_562[45]), .CK(clk_80mhz), 
            .Q(integrator3[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i45.GSR = "ENABLED";
    FD1S3AX integrator3_i46 (.D(integrator3_71__N_562[46]), .CK(clk_80mhz), 
            .Q(integrator3[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i46.GSR = "ENABLED";
    FD1S3AX integrator3_i47 (.D(integrator3_71__N_562[47]), .CK(clk_80mhz), 
            .Q(integrator3[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i47.GSR = "ENABLED";
    FD1S3AX integrator3_i48 (.D(integrator3_71__N_562[48]), .CK(clk_80mhz), 
            .Q(integrator3[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i48.GSR = "ENABLED";
    FD1S3AX integrator3_i49 (.D(integrator3_71__N_562[49]), .CK(clk_80mhz), 
            .Q(integrator3[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i49.GSR = "ENABLED";
    FD1S3AX integrator3_i50 (.D(integrator3_71__N_562[50]), .CK(clk_80mhz), 
            .Q(integrator3[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i50.GSR = "ENABLED";
    FD1S3AX integrator3_i51 (.D(integrator3_71__N_562[51]), .CK(clk_80mhz), 
            .Q(integrator3[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i51.GSR = "ENABLED";
    FD1S3AX integrator3_i52 (.D(integrator3_71__N_562[52]), .CK(clk_80mhz), 
            .Q(integrator3[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i52.GSR = "ENABLED";
    FD1S3AX integrator3_i53 (.D(integrator3_71__N_562[53]), .CK(clk_80mhz), 
            .Q(integrator3[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i53.GSR = "ENABLED";
    FD1S3AX integrator3_i54 (.D(integrator3_71__N_562[54]), .CK(clk_80mhz), 
            .Q(integrator3[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i54.GSR = "ENABLED";
    FD1S3AX integrator3_i55 (.D(integrator3_71__N_562[55]), .CK(clk_80mhz), 
            .Q(integrator3[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i55.GSR = "ENABLED";
    FD1S3AX integrator3_i56 (.D(integrator3_71__N_562[56]), .CK(clk_80mhz), 
            .Q(integrator3[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i56.GSR = "ENABLED";
    FD1S3AX integrator3_i57 (.D(integrator3_71__N_562[57]), .CK(clk_80mhz), 
            .Q(integrator3[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i57.GSR = "ENABLED";
    FD1S3AX integrator3_i58 (.D(integrator3_71__N_562[58]), .CK(clk_80mhz), 
            .Q(integrator3[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i58.GSR = "ENABLED";
    FD1S3AX integrator3_i59 (.D(integrator3_71__N_562[59]), .CK(clk_80mhz), 
            .Q(integrator3[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i59.GSR = "ENABLED";
    FD1S3AX integrator3_i60 (.D(integrator3_71__N_562[60]), .CK(clk_80mhz), 
            .Q(integrator3[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i60.GSR = "ENABLED";
    FD1S3AX integrator3_i61 (.D(integrator3_71__N_562[61]), .CK(clk_80mhz), 
            .Q(integrator3[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i61.GSR = "ENABLED";
    FD1S3AX integrator3_i62 (.D(integrator3_71__N_562[62]), .CK(clk_80mhz), 
            .Q(integrator3[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i62.GSR = "ENABLED";
    FD1S3AX integrator3_i63 (.D(integrator3_71__N_562[63]), .CK(clk_80mhz), 
            .Q(integrator3[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i63.GSR = "ENABLED";
    FD1S3AX integrator3_i64 (.D(integrator3_71__N_562[64]), .CK(clk_80mhz), 
            .Q(integrator3[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i64.GSR = "ENABLED";
    FD1S3AX integrator3_i65 (.D(integrator3_71__N_562[65]), .CK(clk_80mhz), 
            .Q(integrator3[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i65.GSR = "ENABLED";
    FD1S3AX integrator3_i66 (.D(integrator3_71__N_562[66]), .CK(clk_80mhz), 
            .Q(integrator3[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i66.GSR = "ENABLED";
    FD1S3AX integrator3_i67 (.D(integrator3_71__N_562[67]), .CK(clk_80mhz), 
            .Q(integrator3[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i67.GSR = "ENABLED";
    FD1S3AX integrator3_i68 (.D(integrator3_71__N_562[68]), .CK(clk_80mhz), 
            .Q(integrator3[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i68.GSR = "ENABLED";
    FD1S3AX integrator3_i69 (.D(integrator3_71__N_562[69]), .CK(clk_80mhz), 
            .Q(integrator3[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i69.GSR = "ENABLED";
    FD1S3AX integrator3_i70 (.D(integrator3_71__N_562[70]), .CK(clk_80mhz), 
            .Q(integrator3[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i70.GSR = "ENABLED";
    FD1S3AX integrator3_i71 (.D(integrator3_71__N_562[71]), .CK(clk_80mhz), 
            .Q(integrator3[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator3_i71.GSR = "ENABLED";
    FD1S3AX integrator4_i1 (.D(integrator4_71__N_634[1]), .CK(clk_80mhz), 
            .Q(integrator4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i1.GSR = "ENABLED";
    FD1S3AX integrator4_i2 (.D(integrator4_71__N_634[2]), .CK(clk_80mhz), 
            .Q(integrator4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i2.GSR = "ENABLED";
    FD1S3AX integrator4_i3 (.D(integrator4_71__N_634[3]), .CK(clk_80mhz), 
            .Q(integrator4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i3.GSR = "ENABLED";
    FD1S3AX integrator4_i4 (.D(integrator4_71__N_634[4]), .CK(clk_80mhz), 
            .Q(integrator4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i4.GSR = "ENABLED";
    FD1S3AX integrator4_i5 (.D(integrator4_71__N_634[5]), .CK(clk_80mhz), 
            .Q(integrator4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i5.GSR = "ENABLED";
    FD1S3AX integrator4_i6 (.D(integrator4_71__N_634[6]), .CK(clk_80mhz), 
            .Q(integrator4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i6.GSR = "ENABLED";
    FD1S3AX integrator4_i7 (.D(integrator4_71__N_634[7]), .CK(clk_80mhz), 
            .Q(integrator4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i7.GSR = "ENABLED";
    FD1S3AX integrator4_i8 (.D(integrator4_71__N_634[8]), .CK(clk_80mhz), 
            .Q(integrator4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i8.GSR = "ENABLED";
    FD1S3AX integrator4_i9 (.D(integrator4_71__N_634[9]), .CK(clk_80mhz), 
            .Q(integrator4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i9.GSR = "ENABLED";
    FD1S3AX integrator4_i10 (.D(integrator4_71__N_634[10]), .CK(clk_80mhz), 
            .Q(integrator4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i10.GSR = "ENABLED";
    FD1S3AX integrator4_i11 (.D(integrator4_71__N_634[11]), .CK(clk_80mhz), 
            .Q(integrator4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i11.GSR = "ENABLED";
    FD1S3AX integrator4_i12 (.D(integrator4_71__N_634[12]), .CK(clk_80mhz), 
            .Q(integrator4[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i12.GSR = "ENABLED";
    FD1S3AX integrator4_i13 (.D(integrator4_71__N_634[13]), .CK(clk_80mhz), 
            .Q(integrator4[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i13.GSR = "ENABLED";
    FD1S3AX integrator4_i14 (.D(integrator4_71__N_634[14]), .CK(clk_80mhz), 
            .Q(integrator4[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i14.GSR = "ENABLED";
    FD1S3AX integrator4_i15 (.D(integrator4_71__N_634[15]), .CK(clk_80mhz), 
            .Q(integrator4[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i15.GSR = "ENABLED";
    FD1S3AX integrator4_i16 (.D(integrator4_71__N_634[16]), .CK(clk_80mhz), 
            .Q(integrator4[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i16.GSR = "ENABLED";
    FD1S3AX integrator4_i17 (.D(integrator4_71__N_634[17]), .CK(clk_80mhz), 
            .Q(integrator4[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i17.GSR = "ENABLED";
    FD1S3AX integrator4_i18 (.D(integrator4_71__N_634[18]), .CK(clk_80mhz), 
            .Q(integrator4[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i18.GSR = "ENABLED";
    FD1S3AX integrator4_i19 (.D(integrator4_71__N_634[19]), .CK(clk_80mhz), 
            .Q(integrator4[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i19.GSR = "ENABLED";
    FD1S3AX integrator4_i20 (.D(integrator4_71__N_634[20]), .CK(clk_80mhz), 
            .Q(integrator4[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i20.GSR = "ENABLED";
    FD1S3AX integrator4_i21 (.D(integrator4_71__N_634[21]), .CK(clk_80mhz), 
            .Q(integrator4[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i21.GSR = "ENABLED";
    FD1S3AX integrator4_i22 (.D(integrator4_71__N_634[22]), .CK(clk_80mhz), 
            .Q(integrator4[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i22.GSR = "ENABLED";
    FD1S3AX integrator4_i23 (.D(integrator4_71__N_634[23]), .CK(clk_80mhz), 
            .Q(integrator4[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i23.GSR = "ENABLED";
    FD1S3AX integrator4_i24 (.D(integrator4_71__N_634[24]), .CK(clk_80mhz), 
            .Q(integrator4[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i24.GSR = "ENABLED";
    FD1S3AX integrator4_i25 (.D(integrator4_71__N_634[25]), .CK(clk_80mhz), 
            .Q(integrator4[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i25.GSR = "ENABLED";
    FD1S3AX integrator4_i26 (.D(integrator4_71__N_634[26]), .CK(clk_80mhz), 
            .Q(integrator4[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i26.GSR = "ENABLED";
    FD1S3AX integrator4_i27 (.D(integrator4_71__N_634[27]), .CK(clk_80mhz), 
            .Q(integrator4[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i27.GSR = "ENABLED";
    FD1S3AX integrator4_i28 (.D(integrator4_71__N_634[28]), .CK(clk_80mhz), 
            .Q(integrator4[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i28.GSR = "ENABLED";
    FD1S3AX integrator4_i29 (.D(integrator4_71__N_634[29]), .CK(clk_80mhz), 
            .Q(integrator4[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i29.GSR = "ENABLED";
    FD1S3AX integrator4_i30 (.D(integrator4_71__N_634[30]), .CK(clk_80mhz), 
            .Q(integrator4[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i30.GSR = "ENABLED";
    FD1S3AX integrator4_i31 (.D(integrator4_71__N_634[31]), .CK(clk_80mhz), 
            .Q(integrator4[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i31.GSR = "ENABLED";
    FD1S3AX integrator4_i32 (.D(integrator4_71__N_634[32]), .CK(clk_80mhz), 
            .Q(integrator4[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i32.GSR = "ENABLED";
    FD1S3AX integrator4_i33 (.D(integrator4_71__N_634[33]), .CK(clk_80mhz), 
            .Q(integrator4[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i33.GSR = "ENABLED";
    FD1S3AX integrator4_i34 (.D(integrator4_71__N_634[34]), .CK(clk_80mhz), 
            .Q(integrator4[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i34.GSR = "ENABLED";
    FD1S3AX integrator4_i35 (.D(integrator4_71__N_634[35]), .CK(clk_80mhz), 
            .Q(integrator4[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i35.GSR = "ENABLED";
    FD1S3AX integrator4_i36 (.D(integrator4_71__N_634[36]), .CK(clk_80mhz), 
            .Q(integrator4[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i36.GSR = "ENABLED";
    FD1S3AX integrator4_i37 (.D(integrator4_71__N_634[37]), .CK(clk_80mhz), 
            .Q(integrator4[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i37.GSR = "ENABLED";
    FD1S3AX integrator4_i38 (.D(integrator4_71__N_634[38]), .CK(clk_80mhz), 
            .Q(integrator4[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i38.GSR = "ENABLED";
    FD1S3AX integrator4_i39 (.D(integrator4_71__N_634[39]), .CK(clk_80mhz), 
            .Q(integrator4[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i39.GSR = "ENABLED";
    FD1S3AX integrator4_i40 (.D(integrator4_71__N_634[40]), .CK(clk_80mhz), 
            .Q(integrator4[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i40.GSR = "ENABLED";
    FD1S3AX integrator4_i41 (.D(integrator4_71__N_634[41]), .CK(clk_80mhz), 
            .Q(integrator4[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i41.GSR = "ENABLED";
    FD1S3AX integrator4_i42 (.D(integrator4_71__N_634[42]), .CK(clk_80mhz), 
            .Q(integrator4[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i42.GSR = "ENABLED";
    FD1S3AX integrator4_i43 (.D(integrator4_71__N_634[43]), .CK(clk_80mhz), 
            .Q(integrator4[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i43.GSR = "ENABLED";
    FD1S3AX integrator4_i44 (.D(integrator4_71__N_634[44]), .CK(clk_80mhz), 
            .Q(integrator4[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i44.GSR = "ENABLED";
    FD1S3AX integrator4_i45 (.D(integrator4_71__N_634[45]), .CK(clk_80mhz), 
            .Q(integrator4[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i45.GSR = "ENABLED";
    FD1S3AX integrator4_i46 (.D(integrator4_71__N_634[46]), .CK(clk_80mhz), 
            .Q(integrator4[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i46.GSR = "ENABLED";
    FD1S3AX integrator4_i47 (.D(integrator4_71__N_634[47]), .CK(clk_80mhz), 
            .Q(integrator4[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i47.GSR = "ENABLED";
    FD1S3AX integrator4_i48 (.D(integrator4_71__N_634[48]), .CK(clk_80mhz), 
            .Q(integrator4[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i48.GSR = "ENABLED";
    FD1S3AX integrator4_i49 (.D(integrator4_71__N_634[49]), .CK(clk_80mhz), 
            .Q(integrator4[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i49.GSR = "ENABLED";
    FD1S3AX integrator4_i50 (.D(integrator4_71__N_634[50]), .CK(clk_80mhz), 
            .Q(integrator4[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i50.GSR = "ENABLED";
    FD1S3AX integrator4_i51 (.D(integrator4_71__N_634[51]), .CK(clk_80mhz), 
            .Q(integrator4[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i51.GSR = "ENABLED";
    FD1S3AX integrator4_i52 (.D(integrator4_71__N_634[52]), .CK(clk_80mhz), 
            .Q(integrator4[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i52.GSR = "ENABLED";
    FD1S3AX integrator4_i53 (.D(integrator4_71__N_634[53]), .CK(clk_80mhz), 
            .Q(integrator4[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i53.GSR = "ENABLED";
    FD1S3AX integrator4_i54 (.D(integrator4_71__N_634[54]), .CK(clk_80mhz), 
            .Q(integrator4[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i54.GSR = "ENABLED";
    FD1S3AX integrator4_i55 (.D(integrator4_71__N_634[55]), .CK(clk_80mhz), 
            .Q(integrator4[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i55.GSR = "ENABLED";
    FD1S3AX integrator4_i56 (.D(integrator4_71__N_634[56]), .CK(clk_80mhz), 
            .Q(integrator4[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i56.GSR = "ENABLED";
    FD1S3AX integrator4_i57 (.D(integrator4_71__N_634[57]), .CK(clk_80mhz), 
            .Q(integrator4[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i57.GSR = "ENABLED";
    FD1S3AX integrator4_i58 (.D(integrator4_71__N_634[58]), .CK(clk_80mhz), 
            .Q(integrator4[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i58.GSR = "ENABLED";
    FD1S3AX integrator4_i59 (.D(integrator4_71__N_634[59]), .CK(clk_80mhz), 
            .Q(integrator4[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i59.GSR = "ENABLED";
    FD1S3AX integrator4_i60 (.D(integrator4_71__N_634[60]), .CK(clk_80mhz), 
            .Q(integrator4[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i60.GSR = "ENABLED";
    FD1S3AX integrator4_i61 (.D(integrator4_71__N_634[61]), .CK(clk_80mhz), 
            .Q(integrator4[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i61.GSR = "ENABLED";
    FD1S3AX integrator4_i62 (.D(integrator4_71__N_634[62]), .CK(clk_80mhz), 
            .Q(integrator4[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i62.GSR = "ENABLED";
    FD1S3AX integrator4_i63 (.D(integrator4_71__N_634[63]), .CK(clk_80mhz), 
            .Q(integrator4[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i63.GSR = "ENABLED";
    FD1S3AX integrator4_i64 (.D(integrator4_71__N_634[64]), .CK(clk_80mhz), 
            .Q(integrator4[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i64.GSR = "ENABLED";
    FD1S3AX integrator4_i65 (.D(integrator4_71__N_634[65]), .CK(clk_80mhz), 
            .Q(integrator4[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i65.GSR = "ENABLED";
    FD1S3AX integrator4_i66 (.D(integrator4_71__N_634[66]), .CK(clk_80mhz), 
            .Q(integrator4[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i66.GSR = "ENABLED";
    FD1S3AX integrator4_i67 (.D(integrator4_71__N_634[67]), .CK(clk_80mhz), 
            .Q(integrator4[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i67.GSR = "ENABLED";
    FD1S3AX integrator4_i68 (.D(integrator4_71__N_634[68]), .CK(clk_80mhz), 
            .Q(integrator4[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i68.GSR = "ENABLED";
    FD1S3AX integrator4_i69 (.D(integrator4_71__N_634[69]), .CK(clk_80mhz), 
            .Q(integrator4[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i69.GSR = "ENABLED";
    FD1S3AX integrator4_i70 (.D(integrator4_71__N_634[70]), .CK(clk_80mhz), 
            .Q(integrator4[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i70.GSR = "ENABLED";
    FD1S3AX integrator4_i71 (.D(integrator4_71__N_634[71]), .CK(clk_80mhz), 
            .Q(integrator4[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator4_i71.GSR = "ENABLED";
    FD1S3AX integrator5_i1 (.D(integrator5_71__N_706[1]), .CK(clk_80mhz), 
            .Q(integrator5[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i1.GSR = "ENABLED";
    FD1S3AX integrator5_i2 (.D(integrator5_71__N_706[2]), .CK(clk_80mhz), 
            .Q(integrator5[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i2.GSR = "ENABLED";
    FD1S3AX integrator5_i3 (.D(integrator5_71__N_706[3]), .CK(clk_80mhz), 
            .Q(integrator5[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i3.GSR = "ENABLED";
    FD1S3AX integrator5_i4 (.D(integrator5_71__N_706[4]), .CK(clk_80mhz), 
            .Q(integrator5[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i4.GSR = "ENABLED";
    FD1S3AX integrator5_i5 (.D(integrator5_71__N_706[5]), .CK(clk_80mhz), 
            .Q(integrator5[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i5.GSR = "ENABLED";
    FD1S3AX integrator5_i6 (.D(integrator5_71__N_706[6]), .CK(clk_80mhz), 
            .Q(integrator5[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i6.GSR = "ENABLED";
    FD1S3AX integrator5_i7 (.D(integrator5_71__N_706[7]), .CK(clk_80mhz), 
            .Q(integrator5[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i7.GSR = "ENABLED";
    FD1S3AX integrator5_i8 (.D(integrator5_71__N_706[8]), .CK(clk_80mhz), 
            .Q(integrator5[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i8.GSR = "ENABLED";
    FD1S3AX integrator5_i9 (.D(integrator5_71__N_706[9]), .CK(clk_80mhz), 
            .Q(integrator5[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i9.GSR = "ENABLED";
    FD1S3AX integrator5_i10 (.D(integrator5_71__N_706[10]), .CK(clk_80mhz), 
            .Q(integrator5[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i10.GSR = "ENABLED";
    FD1S3AX integrator5_i11 (.D(integrator5_71__N_706[11]), .CK(clk_80mhz), 
            .Q(integrator5[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i11.GSR = "ENABLED";
    FD1S3AX integrator5_i12 (.D(integrator5_71__N_706[12]), .CK(clk_80mhz), 
            .Q(integrator5[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i12.GSR = "ENABLED";
    FD1S3AX integrator5_i13 (.D(integrator5_71__N_706[13]), .CK(clk_80mhz), 
            .Q(integrator5[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i13.GSR = "ENABLED";
    FD1S3AX integrator5_i14 (.D(integrator5_71__N_706[14]), .CK(clk_80mhz), 
            .Q(integrator5[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i14.GSR = "ENABLED";
    FD1S3AX integrator5_i15 (.D(integrator5_71__N_706[15]), .CK(clk_80mhz), 
            .Q(integrator5[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i15.GSR = "ENABLED";
    FD1S3AX integrator5_i16 (.D(integrator5_71__N_706[16]), .CK(clk_80mhz), 
            .Q(integrator5[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i16.GSR = "ENABLED";
    FD1S3AX integrator5_i17 (.D(integrator5_71__N_706[17]), .CK(clk_80mhz), 
            .Q(integrator5[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i17.GSR = "ENABLED";
    FD1S3AX integrator5_i18 (.D(integrator5_71__N_706[18]), .CK(clk_80mhz), 
            .Q(integrator5[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i18.GSR = "ENABLED";
    FD1S3AX integrator5_i19 (.D(integrator5_71__N_706[19]), .CK(clk_80mhz), 
            .Q(integrator5[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i19.GSR = "ENABLED";
    FD1S3AX integrator5_i20 (.D(integrator5_71__N_706[20]), .CK(clk_80mhz), 
            .Q(integrator5[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i20.GSR = "ENABLED";
    FD1S3AX integrator5_i21 (.D(integrator5_71__N_706[21]), .CK(clk_80mhz), 
            .Q(integrator5[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i21.GSR = "ENABLED";
    FD1S3AX integrator5_i22 (.D(integrator5_71__N_706[22]), .CK(clk_80mhz), 
            .Q(integrator5[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i22.GSR = "ENABLED";
    FD1S3AX integrator5_i23 (.D(integrator5_71__N_706[23]), .CK(clk_80mhz), 
            .Q(integrator5[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i23.GSR = "ENABLED";
    FD1S3AX integrator5_i24 (.D(integrator5_71__N_706[24]), .CK(clk_80mhz), 
            .Q(integrator5[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i24.GSR = "ENABLED";
    FD1S3AX integrator5_i25 (.D(integrator5_71__N_706[25]), .CK(clk_80mhz), 
            .Q(integrator5[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i25.GSR = "ENABLED";
    FD1S3AX integrator5_i26 (.D(integrator5_71__N_706[26]), .CK(clk_80mhz), 
            .Q(integrator5[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i26.GSR = "ENABLED";
    FD1S3AX integrator5_i27 (.D(integrator5_71__N_706[27]), .CK(clk_80mhz), 
            .Q(integrator5[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i27.GSR = "ENABLED";
    FD1S3AX integrator5_i28 (.D(integrator5_71__N_706[28]), .CK(clk_80mhz), 
            .Q(integrator5[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i28.GSR = "ENABLED";
    FD1S3AX integrator5_i29 (.D(integrator5_71__N_706[29]), .CK(clk_80mhz), 
            .Q(integrator5[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i29.GSR = "ENABLED";
    FD1S3AX integrator5_i30 (.D(integrator5_71__N_706[30]), .CK(clk_80mhz), 
            .Q(integrator5[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i30.GSR = "ENABLED";
    FD1S3AX integrator5_i31 (.D(integrator5_71__N_706[31]), .CK(clk_80mhz), 
            .Q(integrator5[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i31.GSR = "ENABLED";
    FD1S3AX integrator5_i32 (.D(integrator5_71__N_706[32]), .CK(clk_80mhz), 
            .Q(integrator5[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i32.GSR = "ENABLED";
    FD1S3AX integrator5_i33 (.D(integrator5_71__N_706[33]), .CK(clk_80mhz), 
            .Q(integrator5[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i33.GSR = "ENABLED";
    FD1S3AX integrator5_i34 (.D(integrator5_71__N_706[34]), .CK(clk_80mhz), 
            .Q(integrator5[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i34.GSR = "ENABLED";
    FD1S3AX integrator5_i35 (.D(integrator5_71__N_706[35]), .CK(clk_80mhz), 
            .Q(integrator5[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i35.GSR = "ENABLED";
    FD1S3AX integrator5_i36 (.D(integrator5_71__N_706[36]), .CK(clk_80mhz), 
            .Q(integrator5[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i36.GSR = "ENABLED";
    FD1S3AX integrator5_i37 (.D(integrator5_71__N_706[37]), .CK(clk_80mhz), 
            .Q(integrator5[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i37.GSR = "ENABLED";
    FD1S3AX integrator5_i38 (.D(integrator5_71__N_706[38]), .CK(clk_80mhz), 
            .Q(integrator5[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i38.GSR = "ENABLED";
    FD1S3AX integrator5_i39 (.D(integrator5_71__N_706[39]), .CK(clk_80mhz), 
            .Q(integrator5[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i39.GSR = "ENABLED";
    FD1S3AX integrator5_i40 (.D(integrator5_71__N_706[40]), .CK(clk_80mhz), 
            .Q(integrator5[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i40.GSR = "ENABLED";
    FD1S3AX integrator5_i41 (.D(integrator5_71__N_706[41]), .CK(clk_80mhz), 
            .Q(integrator5[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i41.GSR = "ENABLED";
    FD1S3AX integrator5_i42 (.D(integrator5_71__N_706[42]), .CK(clk_80mhz), 
            .Q(integrator5[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i42.GSR = "ENABLED";
    FD1S3AX integrator5_i43 (.D(integrator5_71__N_706[43]), .CK(clk_80mhz), 
            .Q(integrator5[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i43.GSR = "ENABLED";
    FD1S3AX integrator5_i44 (.D(integrator5_71__N_706[44]), .CK(clk_80mhz), 
            .Q(integrator5[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i44.GSR = "ENABLED";
    FD1S3AX integrator5_i45 (.D(integrator5_71__N_706[45]), .CK(clk_80mhz), 
            .Q(integrator5[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i45.GSR = "ENABLED";
    FD1S3AX integrator5_i46 (.D(integrator5_71__N_706[46]), .CK(clk_80mhz), 
            .Q(integrator5[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i46.GSR = "ENABLED";
    FD1S3AX integrator5_i47 (.D(integrator5_71__N_706[47]), .CK(clk_80mhz), 
            .Q(integrator5[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i47.GSR = "ENABLED";
    FD1S3AX integrator5_i48 (.D(integrator5_71__N_706[48]), .CK(clk_80mhz), 
            .Q(integrator5[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i48.GSR = "ENABLED";
    FD1S3AX integrator5_i49 (.D(integrator5_71__N_706[49]), .CK(clk_80mhz), 
            .Q(integrator5[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i49.GSR = "ENABLED";
    FD1S3AX integrator5_i50 (.D(integrator5_71__N_706[50]), .CK(clk_80mhz), 
            .Q(integrator5[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i50.GSR = "ENABLED";
    FD1S3AX integrator5_i51 (.D(integrator5_71__N_706[51]), .CK(clk_80mhz), 
            .Q(integrator5[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i51.GSR = "ENABLED";
    FD1S3AX integrator5_i52 (.D(integrator5_71__N_706[52]), .CK(clk_80mhz), 
            .Q(integrator5[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i52.GSR = "ENABLED";
    FD1S3AX integrator5_i53 (.D(integrator5_71__N_706[53]), .CK(clk_80mhz), 
            .Q(integrator5[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i53.GSR = "ENABLED";
    FD1S3AX integrator5_i54 (.D(integrator5_71__N_706[54]), .CK(clk_80mhz), 
            .Q(integrator5[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i54.GSR = "ENABLED";
    FD1S3AX integrator5_i55 (.D(integrator5_71__N_706[55]), .CK(clk_80mhz), 
            .Q(integrator5[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i55.GSR = "ENABLED";
    FD1S3AX integrator5_i56 (.D(integrator5_71__N_706[56]), .CK(clk_80mhz), 
            .Q(integrator5[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i56.GSR = "ENABLED";
    FD1S3AX integrator5_i57 (.D(integrator5_71__N_706[57]), .CK(clk_80mhz), 
            .Q(integrator5[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i57.GSR = "ENABLED";
    FD1S3AX integrator5_i58 (.D(integrator5_71__N_706[58]), .CK(clk_80mhz), 
            .Q(integrator5[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i58.GSR = "ENABLED";
    FD1S3AX integrator5_i59 (.D(integrator5_71__N_706[59]), .CK(clk_80mhz), 
            .Q(integrator5[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i59.GSR = "ENABLED";
    FD1S3AX integrator5_i60 (.D(integrator5_71__N_706[60]), .CK(clk_80mhz), 
            .Q(integrator5[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i60.GSR = "ENABLED";
    FD1S3AX integrator5_i61 (.D(integrator5_71__N_706[61]), .CK(clk_80mhz), 
            .Q(integrator5[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i61.GSR = "ENABLED";
    FD1S3AX integrator5_i62 (.D(integrator5_71__N_706[62]), .CK(clk_80mhz), 
            .Q(integrator5[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i62.GSR = "ENABLED";
    FD1S3AX integrator5_i63 (.D(integrator5_71__N_706[63]), .CK(clk_80mhz), 
            .Q(integrator5[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i63.GSR = "ENABLED";
    FD1S3AX integrator5_i64 (.D(integrator5_71__N_706[64]), .CK(clk_80mhz), 
            .Q(integrator5[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i64.GSR = "ENABLED";
    FD1S3AX integrator5_i65 (.D(integrator5_71__N_706[65]), .CK(clk_80mhz), 
            .Q(integrator5[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i65.GSR = "ENABLED";
    FD1S3AX integrator5_i66 (.D(integrator5_71__N_706[66]), .CK(clk_80mhz), 
            .Q(integrator5[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i66.GSR = "ENABLED";
    FD1S3AX integrator5_i67 (.D(integrator5_71__N_706[67]), .CK(clk_80mhz), 
            .Q(integrator5[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i67.GSR = "ENABLED";
    FD1S3AX integrator5_i68 (.D(integrator5_71__N_706[68]), .CK(clk_80mhz), 
            .Q(integrator5[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i68.GSR = "ENABLED";
    FD1S3AX integrator5_i69 (.D(integrator5_71__N_706[69]), .CK(clk_80mhz), 
            .Q(integrator5[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i69.GSR = "ENABLED";
    FD1S3AX integrator5_i70 (.D(integrator5_71__N_706[70]), .CK(clk_80mhz), 
            .Q(integrator5[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i70.GSR = "ENABLED";
    FD1S3AX integrator5_i71 (.D(integrator5_71__N_706[71]), .CK(clk_80mhz), 
            .Q(integrator5[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator5_i71.GSR = "ENABLED";
    FD1P3AX comb6_i0_i1 (.D(comb6_71__N_1451[1]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i1.GSR = "ENABLED";
    FD1P3AX comb6_i0_i2 (.D(comb6_71__N_1451[2]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i2.GSR = "ENABLED";
    FD1P3AX comb6_i0_i3 (.D(comb6_71__N_1451[3]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i3.GSR = "ENABLED";
    FD1P3AX comb6_i0_i4 (.D(comb6_71__N_1451[4]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i4.GSR = "ENABLED";
    FD1P3AX comb6_i0_i5 (.D(comb6_71__N_1451[5]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i5.GSR = "ENABLED";
    FD1P3AX comb6_i0_i6 (.D(comb6_71__N_1451[6]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i6.GSR = "ENABLED";
    FD1P3AX comb6_i0_i7 (.D(comb6_71__N_1451[7]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i7.GSR = "ENABLED";
    FD1P3AX comb6_i0_i8 (.D(comb6_71__N_1451[8]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i8.GSR = "ENABLED";
    FD1P3AX comb6_i0_i9 (.D(comb6_71__N_1451[9]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i9.GSR = "ENABLED";
    FD1P3AX comb6_i0_i10 (.D(comb6_71__N_1451[10]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i10.GSR = "ENABLED";
    FD1P3AX comb6_i0_i11 (.D(comb6_71__N_1451[11]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i11.GSR = "ENABLED";
    FD1P3AX comb6_i0_i12 (.D(comb6_71__N_1451[12]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i12.GSR = "ENABLED";
    FD1P3AX comb6_i0_i13 (.D(comb6_71__N_1451[13]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i13.GSR = "ENABLED";
    FD1P3AX comb6_i0_i14 (.D(comb6_71__N_1451[14]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i14.GSR = "ENABLED";
    FD1P3AX comb6_i0_i15 (.D(comb6_71__N_1451[15]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i15.GSR = "ENABLED";
    FD1P3AX comb6_i0_i16 (.D(comb6_71__N_1451[16]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i16.GSR = "ENABLED";
    FD1P3AX comb6_i0_i17 (.D(comb6_71__N_1451[17]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i17.GSR = "ENABLED";
    FD1P3AX comb6_i0_i18 (.D(comb6_71__N_1451[18]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i18.GSR = "ENABLED";
    FD1P3AX comb6_i0_i19 (.D(comb6_71__N_1451[19]), .SP(clk_80mhz_enable_884), 
            .CK(clk_80mhz), .Q(comb6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i19.GSR = "ENABLED";
    FD1P3AX comb6_i0_i20 (.D(comb6_71__N_1451[20]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i20.GSR = "ENABLED";
    FD1P3AX comb6_i0_i21 (.D(comb6_71__N_1451[21]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i21.GSR = "ENABLED";
    FD1P3AX comb6_i0_i22 (.D(comb6_71__N_1451[22]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i22.GSR = "ENABLED";
    FD1P3AX comb6_i0_i23 (.D(comb6_71__N_1451[23]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i23.GSR = "ENABLED";
    FD1P3AX comb6_i0_i24 (.D(comb6_71__N_1451[24]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i24.GSR = "ENABLED";
    FD1P3AX comb6_i0_i25 (.D(comb6_71__N_1451[25]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i25.GSR = "ENABLED";
    FD1P3AX comb6_i0_i26 (.D(comb6_71__N_1451[26]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i26.GSR = "ENABLED";
    FD1P3AX comb6_i0_i27 (.D(comb6_71__N_1451[27]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i27.GSR = "ENABLED";
    FD1P3AX comb6_i0_i28 (.D(comb6_71__N_1451[28]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i28.GSR = "ENABLED";
    FD1P3AX comb6_i0_i29 (.D(comb6_71__N_1451[29]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i29.GSR = "ENABLED";
    FD1P3AX comb6_i0_i30 (.D(comb6_71__N_1451[30]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i30.GSR = "ENABLED";
    FD1P3AX comb6_i0_i31 (.D(comb6_71__N_1451[31]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i31.GSR = "ENABLED";
    FD1P3AX comb6_i0_i32 (.D(comb6_71__N_1451[32]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i32.GSR = "ENABLED";
    FD1P3AX comb6_i0_i33 (.D(comb6_71__N_1451[33]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i33.GSR = "ENABLED";
    FD1P3AX comb6_i0_i34 (.D(comb6_71__N_1451[34]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i34.GSR = "ENABLED";
    FD1P3AX comb6_i0_i35 (.D(comb6_71__N_1451[35]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i35.GSR = "ENABLED";
    FD1P3AX comb6_i0_i36 (.D(comb6_71__N_1451[36]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i36.GSR = "ENABLED";
    FD1P3AX comb6_i0_i37 (.D(comb6_71__N_1451[37]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i37.GSR = "ENABLED";
    FD1P3AX comb6_i0_i38 (.D(comb6_71__N_1451[38]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i38.GSR = "ENABLED";
    FD1P3AX comb6_i0_i39 (.D(comb6_71__N_1451[39]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i39.GSR = "ENABLED";
    FD1P3AX comb6_i0_i40 (.D(comb6_71__N_1451[40]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i40.GSR = "ENABLED";
    FD1P3AX comb6_i0_i41 (.D(comb6_71__N_1451[41]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i41.GSR = "ENABLED";
    FD1P3AX comb6_i0_i42 (.D(comb6_71__N_1451[42]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i42.GSR = "ENABLED";
    FD1P3AX comb6_i0_i43 (.D(comb6_71__N_1451[43]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i43.GSR = "ENABLED";
    FD1P3AX comb6_i0_i44 (.D(comb6_71__N_1451[44]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i44.GSR = "ENABLED";
    FD1P3AX comb6_i0_i45 (.D(comb6_71__N_1451[45]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i45.GSR = "ENABLED";
    FD1P3AX comb6_i0_i46 (.D(comb6_71__N_1451[46]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i46.GSR = "ENABLED";
    FD1P3AX comb6_i0_i47 (.D(comb6_71__N_1451[47]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i47.GSR = "ENABLED";
    FD1P3AX comb6_i0_i48 (.D(comb6_71__N_1451[48]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i48.GSR = "ENABLED";
    FD1P3AX comb6_i0_i49 (.D(comb6_71__N_1451[49]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i49.GSR = "ENABLED";
    FD1P3AX comb6_i0_i50 (.D(comb6_71__N_1451[50]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i50.GSR = "ENABLED";
    FD1P3AX comb6_i0_i51 (.D(comb6_71__N_1451[51]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i51.GSR = "ENABLED";
    FD1P3AX comb6_i0_i52 (.D(comb6_71__N_1451[52]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i52.GSR = "ENABLED";
    FD1P3AX comb6_i0_i53 (.D(comb6_71__N_1451[53]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i53.GSR = "ENABLED";
    FD1P3AX comb6_i0_i54 (.D(comb6_71__N_1451[54]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i54.GSR = "ENABLED";
    FD1P3AX comb6_i0_i55 (.D(comb6_71__N_1451[55]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i55.GSR = "ENABLED";
    FD1P3AX comb6_i0_i56 (.D(comb6_71__N_1451[56]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i56.GSR = "ENABLED";
    FD1P3AX comb6_i0_i57 (.D(comb6_71__N_1451[57]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i57.GSR = "ENABLED";
    FD1P3AX comb6_i0_i58 (.D(comb6_71__N_1451[58]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i58.GSR = "ENABLED";
    FD1P3AX comb6_i0_i59 (.D(comb6_71__N_1451[59]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i59.GSR = "ENABLED";
    FD1P3AX comb6_i0_i60 (.D(comb6_71__N_1451[60]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i60.GSR = "ENABLED";
    FD1P3AX comb6_i0_i61 (.D(comb6_71__N_1451[61]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i61.GSR = "ENABLED";
    FD1P3AX comb6_i0_i62 (.D(comb6_71__N_1451[62]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i62.GSR = "ENABLED";
    FD1P3AX comb6_i0_i63 (.D(comb6_71__N_1451[63]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i63.GSR = "ENABLED";
    FD1P3AX comb6_i0_i64 (.D(comb6_71__N_1451[64]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i64.GSR = "ENABLED";
    FD1P3AX comb6_i0_i65 (.D(comb6_71__N_1451[65]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i65.GSR = "ENABLED";
    FD1P3AX comb6_i0_i66 (.D(comb6_71__N_1451[66]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i66.GSR = "ENABLED";
    FD1P3AX comb6_i0_i67 (.D(comb6_71__N_1451[67]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i67.GSR = "ENABLED";
    FD1P3AX comb6_i0_i68 (.D(comb6_71__N_1451[68]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i68.GSR = "ENABLED";
    FD1P3AX comb6_i0_i69 (.D(comb6_71__N_1451[69]), .SP(clk_80mhz_enable_934), 
            .CK(clk_80mhz), .Q(comb6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i69.GSR = "ENABLED";
    FD1P3AX comb6_i0_i70 (.D(comb6_71__N_1451[70]), .SP(clk_80mhz_enable_984), 
            .CK(clk_80mhz), .Q(comb6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i70.GSR = "ENABLED";
    FD1P3AX comb6_i0_i71 (.D(comb6_71__N_1451[71]), .SP(clk_80mhz_enable_984), 
            .CK(clk_80mhz), .Q(comb6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb6_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i1 (.D(comb6[1]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i2 (.D(comb6[2]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i3 (.D(comb6[3]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i4 (.D(comb6[4]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i5 (.D(comb6[5]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i6 (.D(comb6[6]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i7 (.D(comb6[7]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i8 (.D(comb6[8]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i9 (.D(comb6[9]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i10 (.D(comb6[10]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i11 (.D(comb6[11]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i12 (.D(comb6[12]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i13 (.D(comb6[13]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i14 (.D(comb6[14]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i15 (.D(comb6[15]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i16 (.D(comb6[16]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i17 (.D(comb6[17]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i18 (.D(comb6[18]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i19 (.D(comb6[19]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i20 (.D(comb6[20]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i21 (.D(comb6[21]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i22 (.D(comb6[22]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i23 (.D(comb6[23]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i24 (.D(comb6[24]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i25 (.D(comb6[25]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i26 (.D(comb6[26]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i27 (.D(comb6[27]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i28 (.D(comb6[28]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i29 (.D(comb6[29]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i30 (.D(comb6[30]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i31 (.D(comb6[31]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i32 (.D(comb6[32]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i33 (.D(comb6[33]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i34 (.D(comb6[34]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i35 (.D(comb6[35]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i36 (.D(comb6[36]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i37 (.D(comb6[37]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i38 (.D(comb6[38]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i39 (.D(comb6[39]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i40 (.D(comb6[40]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i41 (.D(comb6[41]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i42 (.D(comb6[42]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i43 (.D(comb6[43]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i44 (.D(comb6[44]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i45 (.D(comb6[45]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i46 (.D(comb6[46]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i47 (.D(comb6[47]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i48 (.D(comb6[48]), .SP(clk_80mhz_enable_984), .CK(clk_80mhz), 
            .Q(comb_d6[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i49 (.D(comb6[49]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i50 (.D(comb6[50]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i51 (.D(comb6[51]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i52 (.D(comb6[52]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i53 (.D(comb6[53]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i54 (.D(comb6[54]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i55 (.D(comb6[55]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i56 (.D(comb6[56]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i57 (.D(comb6[57]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i58 (.D(comb6[58]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i59 (.D(comb6[59]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i60 (.D(comb6[60]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i61 (.D(comb6[61]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i62 (.D(comb6[62]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i63 (.D(comb6[63]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i64 (.D(comb6[64]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i65 (.D(comb6[65]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i66 (.D(comb6[66]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i67 (.D(comb6[67]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i68 (.D(comb6[68]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i69 (.D(comb6[69]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i70 (.D(comb6[70]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d6_i0_i71 (.D(comb6[71]), .SP(clk_80mhz_enable_1034), .CK(clk_80mhz), 
            .Q(comb_d6[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d6_i0_i71.GSR = "ENABLED";
    FD1P3AX comb7_i0_i1 (.D(comb7_71__N_1523[1]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i1.GSR = "ENABLED";
    FD1P3AX comb7_i0_i2 (.D(comb7_71__N_1523[2]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i2.GSR = "ENABLED";
    FD1P3AX comb7_i0_i3 (.D(comb7_71__N_1523[3]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i3.GSR = "ENABLED";
    FD1P3AX comb7_i0_i4 (.D(comb7_71__N_1523[4]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i4.GSR = "ENABLED";
    FD1P3AX comb7_i0_i5 (.D(comb7_71__N_1523[5]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i5.GSR = "ENABLED";
    FD1P3AX comb7_i0_i6 (.D(comb7_71__N_1523[6]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i6.GSR = "ENABLED";
    FD1P3AX comb7_i0_i7 (.D(comb7_71__N_1523[7]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i7.GSR = "ENABLED";
    FD1P3AX comb7_i0_i8 (.D(comb7_71__N_1523[8]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i8.GSR = "ENABLED";
    FD1P3AX comb7_i0_i9 (.D(comb7_71__N_1523[9]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i9.GSR = "ENABLED";
    FD1P3AX comb7_i0_i10 (.D(comb7_71__N_1523[10]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i10.GSR = "ENABLED";
    FD1P3AX comb7_i0_i11 (.D(comb7_71__N_1523[11]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i11.GSR = "ENABLED";
    FD1P3AX comb7_i0_i12 (.D(comb7_71__N_1523[12]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i12.GSR = "ENABLED";
    FD1P3AX comb7_i0_i13 (.D(comb7_71__N_1523[13]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i13.GSR = "ENABLED";
    FD1P3AX comb7_i0_i14 (.D(comb7_71__N_1523[14]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i14.GSR = "ENABLED";
    FD1P3AX comb7_i0_i15 (.D(comb7_71__N_1523[15]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i15.GSR = "ENABLED";
    FD1P3AX comb7_i0_i16 (.D(comb7_71__N_1523[16]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i16.GSR = "ENABLED";
    FD1P3AX comb7_i0_i17 (.D(comb7_71__N_1523[17]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i17.GSR = "ENABLED";
    FD1P3AX comb7_i0_i18 (.D(comb7_71__N_1523[18]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i18.GSR = "ENABLED";
    FD1P3AX comb7_i0_i19 (.D(comb7_71__N_1523[19]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i19.GSR = "ENABLED";
    FD1P3AX comb7_i0_i20 (.D(comb7_71__N_1523[20]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i20.GSR = "ENABLED";
    FD1P3AX comb7_i0_i21 (.D(comb7_71__N_1523[21]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i21.GSR = "ENABLED";
    FD1P3AX comb7_i0_i22 (.D(comb7_71__N_1523[22]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i22.GSR = "ENABLED";
    FD1P3AX comb7_i0_i23 (.D(comb7_71__N_1523[23]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i23.GSR = "ENABLED";
    FD1P3AX comb7_i0_i24 (.D(comb7_71__N_1523[24]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i24.GSR = "ENABLED";
    FD1P3AX comb7_i0_i25 (.D(comb7_71__N_1523[25]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i25.GSR = "ENABLED";
    FD1P3AX comb7_i0_i26 (.D(comb7_71__N_1523[26]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i26.GSR = "ENABLED";
    FD1P3AX comb7_i0_i27 (.D(comb7_71__N_1523[27]), .SP(clk_80mhz_enable_1034), 
            .CK(clk_80mhz), .Q(comb7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i27.GSR = "ENABLED";
    FD1P3AX comb7_i0_i28 (.D(comb7_71__N_1523[28]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i28.GSR = "ENABLED";
    FD1P3AX comb7_i0_i29 (.D(comb7_71__N_1523[29]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i29.GSR = "ENABLED";
    FD1P3AX comb7_i0_i30 (.D(comb7_71__N_1523[30]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i30.GSR = "ENABLED";
    FD1P3AX comb7_i0_i31 (.D(comb7_71__N_1523[31]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i31.GSR = "ENABLED";
    FD1P3AX comb7_i0_i32 (.D(comb7_71__N_1523[32]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i32.GSR = "ENABLED";
    FD1P3AX comb7_i0_i33 (.D(comb7_71__N_1523[33]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i33.GSR = "ENABLED";
    FD1P3AX comb7_i0_i34 (.D(comb7_71__N_1523[34]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i34.GSR = "ENABLED";
    FD1P3AX comb7_i0_i35 (.D(comb7_71__N_1523[35]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i35.GSR = "ENABLED";
    FD1P3AX comb7_i0_i36 (.D(comb7_71__N_1523[36]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i36.GSR = "ENABLED";
    FD1P3AX comb7_i0_i37 (.D(comb7_71__N_1523[37]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i37.GSR = "ENABLED";
    FD1P3AX comb7_i0_i38 (.D(comb7_71__N_1523[38]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i38.GSR = "ENABLED";
    FD1P3AX comb7_i0_i39 (.D(comb7_71__N_1523[39]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i39.GSR = "ENABLED";
    FD1P3AX comb7_i0_i40 (.D(comb7_71__N_1523[40]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i40.GSR = "ENABLED";
    FD1P3AX comb7_i0_i41 (.D(comb7_71__N_1523[41]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i41.GSR = "ENABLED";
    FD1P3AX comb7_i0_i42 (.D(comb7_71__N_1523[42]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i42.GSR = "ENABLED";
    FD1P3AX comb7_i0_i43 (.D(comb7_71__N_1523[43]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i43.GSR = "ENABLED";
    FD1P3AX comb7_i0_i44 (.D(comb7_71__N_1523[44]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i44.GSR = "ENABLED";
    FD1P3AX comb7_i0_i45 (.D(comb7_71__N_1523[45]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i45.GSR = "ENABLED";
    FD1P3AX comb7_i0_i46 (.D(comb7_71__N_1523[46]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i46.GSR = "ENABLED";
    FD1P3AX comb7_i0_i47 (.D(comb7_71__N_1523[47]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i47.GSR = "ENABLED";
    FD1P3AX comb7_i0_i48 (.D(comb7_71__N_1523[48]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i48.GSR = "ENABLED";
    FD1P3AX comb7_i0_i49 (.D(comb7_71__N_1523[49]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i49.GSR = "ENABLED";
    FD1P3AX comb7_i0_i50 (.D(comb7_71__N_1523[50]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i50.GSR = "ENABLED";
    FD1P3AX comb7_i0_i51 (.D(comb7_71__N_1523[51]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i51.GSR = "ENABLED";
    FD1P3AX comb7_i0_i52 (.D(comb7_71__N_1523[52]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i52.GSR = "ENABLED";
    FD1P3AX comb7_i0_i53 (.D(comb7_71__N_1523[53]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i53.GSR = "ENABLED";
    FD1P3AX comb7_i0_i54 (.D(comb7_71__N_1523[54]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i54.GSR = "ENABLED";
    FD1P3AX comb7_i0_i55 (.D(comb7_71__N_1523[55]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i55.GSR = "ENABLED";
    FD1P3AX comb7_i0_i56 (.D(comb7_71__N_1523[56]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i56.GSR = "ENABLED";
    FD1P3AX comb7_i0_i57 (.D(comb7_71__N_1523[57]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i57.GSR = "ENABLED";
    FD1P3AX comb7_i0_i58 (.D(comb7_71__N_1523[58]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i58.GSR = "ENABLED";
    FD1P3AX comb7_i0_i59 (.D(comb7_71__N_1523[59]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i59.GSR = "ENABLED";
    FD1P3AX comb7_i0_i60 (.D(comb7_71__N_1523[60]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i60.GSR = "ENABLED";
    FD1P3AX comb7_i0_i61 (.D(comb7_71__N_1523[61]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i61.GSR = "ENABLED";
    FD1P3AX comb7_i0_i62 (.D(comb7_71__N_1523[62]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i62.GSR = "ENABLED";
    FD1P3AX comb7_i0_i63 (.D(comb7_71__N_1523[63]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i63.GSR = "ENABLED";
    FD1P3AX comb7_i0_i64 (.D(comb7_71__N_1523[64]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i64.GSR = "ENABLED";
    FD1P3AX comb7_i0_i65 (.D(comb7_71__N_1523[65]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i65.GSR = "ENABLED";
    FD1P3AX comb7_i0_i66 (.D(comb7_71__N_1523[66]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i66.GSR = "ENABLED";
    FD1P3AX comb7_i0_i67 (.D(comb7_71__N_1523[67]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i67.GSR = "ENABLED";
    FD1P3AX comb7_i0_i68 (.D(comb7_71__N_1523[68]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i68.GSR = "ENABLED";
    FD1P3AX comb7_i0_i69 (.D(comb7_71__N_1523[69]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i69.GSR = "ENABLED";
    FD1P3AX comb7_i0_i70 (.D(comb7_71__N_1523[70]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i70.GSR = "ENABLED";
    FD1P3AX comb7_i0_i71 (.D(comb7_71__N_1523[71]), .SP(clk_80mhz_enable_1084), 
            .CK(clk_80mhz), .Q(comb7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb7_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i1 (.D(comb7[1]), .SP(clk_80mhz_enable_1084), .CK(clk_80mhz), 
            .Q(comb_d7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i2 (.D(comb7[2]), .SP(clk_80mhz_enable_1084), .CK(clk_80mhz), 
            .Q(comb_d7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i3 (.D(comb7[3]), .SP(clk_80mhz_enable_1084), .CK(clk_80mhz), 
            .Q(comb_d7[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i4 (.D(comb7[4]), .SP(clk_80mhz_enable_1084), .CK(clk_80mhz), 
            .Q(comb_d7[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i5 (.D(comb7[5]), .SP(clk_80mhz_enable_1084), .CK(clk_80mhz), 
            .Q(comb_d7[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i6 (.D(comb7[6]), .SP(clk_80mhz_enable_1084), .CK(clk_80mhz), 
            .Q(comb_d7[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i7 (.D(comb7[7]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i8 (.D(comb7[8]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i9 (.D(comb7[9]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i10 (.D(comb7[10]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i11 (.D(comb7[11]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i12 (.D(comb7[12]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i13 (.D(comb7[13]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i14 (.D(comb7[14]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i15 (.D(comb7[15]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i16 (.D(comb7[16]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i17 (.D(comb7[17]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i18 (.D(comb7[18]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i19 (.D(comb7[19]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i20 (.D(comb7[20]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i21 (.D(comb7[21]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i22 (.D(comb7[22]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i23 (.D(comb7[23]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i24 (.D(comb7[24]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i25 (.D(comb7[25]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i26 (.D(comb7[26]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i27 (.D(comb7[27]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i28 (.D(comb7[28]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i29 (.D(comb7[29]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i30 (.D(comb7[30]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i31 (.D(comb7[31]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i32 (.D(comb7[32]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i33 (.D(comb7[33]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i34 (.D(comb7[34]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i35 (.D(comb7[35]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i36 (.D(comb7[36]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i37 (.D(comb7[37]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i38 (.D(comb7[38]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i39 (.D(comb7[39]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i40 (.D(comb7[40]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i41 (.D(comb7[41]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i42 (.D(comb7[42]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i43 (.D(comb7[43]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i44 (.D(comb7[44]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i45 (.D(comb7[45]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i46 (.D(comb7[46]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i47 (.D(comb7[47]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i48 (.D(comb7[48]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i49 (.D(comb7[49]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i50 (.D(comb7[50]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i51 (.D(comb7[51]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i52 (.D(comb7[52]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i53 (.D(comb7[53]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i54 (.D(comb7[54]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i55 (.D(comb7[55]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i56 (.D(comb7[56]), .SP(clk_80mhz_enable_1134), .CK(clk_80mhz), 
            .Q(comb_d7[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i57 (.D(comb7[57]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i58 (.D(comb7[58]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i59 (.D(comb7[59]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i60 (.D(comb7[60]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i61 (.D(comb7[61]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i62 (.D(comb7[62]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i63 (.D(comb7[63]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i64 (.D(comb7[64]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i65 (.D(comb7[65]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i66 (.D(comb7[66]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i67 (.D(comb7[67]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i68 (.D(comb7[68]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i69 (.D(comb7[69]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i70 (.D(comb7[70]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d7_i0_i71 (.D(comb7[71]), .SP(clk_80mhz_enable_1184), .CK(clk_80mhz), 
            .Q(comb_d7[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d7_i0_i71.GSR = "ENABLED";
    FD1P3AX comb8_i0_i1 (.D(comb8_71__N_1595[1]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i1.GSR = "ENABLED";
    FD1P3AX comb8_i0_i2 (.D(comb8_71__N_1595[2]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i2.GSR = "ENABLED";
    FD1P3AX comb8_i0_i3 (.D(comb8_71__N_1595[3]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i3.GSR = "ENABLED";
    FD1P3AX comb8_i0_i4 (.D(comb8_71__N_1595[4]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i4.GSR = "ENABLED";
    FD1P3AX comb8_i0_i5 (.D(comb8_71__N_1595[5]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i5.GSR = "ENABLED";
    FD1P3AX comb8_i0_i6 (.D(comb8_71__N_1595[6]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i6.GSR = "ENABLED";
    FD1P3AX comb8_i0_i7 (.D(comb8_71__N_1595[7]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i7.GSR = "ENABLED";
    FD1P3AX comb8_i0_i8 (.D(comb8_71__N_1595[8]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i8.GSR = "ENABLED";
    FD1P3AX comb8_i0_i9 (.D(comb8_71__N_1595[9]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i9.GSR = "ENABLED";
    FD1P3AX comb8_i0_i10 (.D(comb8_71__N_1595[10]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i10.GSR = "ENABLED";
    FD1P3AX comb8_i0_i11 (.D(comb8_71__N_1595[11]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i11.GSR = "ENABLED";
    FD1P3AX comb8_i0_i12 (.D(comb8_71__N_1595[12]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i12.GSR = "ENABLED";
    FD1P3AX comb8_i0_i13 (.D(comb8_71__N_1595[13]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i13.GSR = "ENABLED";
    FD1P3AX comb8_i0_i14 (.D(comb8_71__N_1595[14]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i14.GSR = "ENABLED";
    FD1P3AX comb8_i0_i15 (.D(comb8_71__N_1595[15]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i15.GSR = "ENABLED";
    FD1P3AX comb8_i0_i16 (.D(comb8_71__N_1595[16]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i16.GSR = "ENABLED";
    FD1P3AX comb8_i0_i17 (.D(comb8_71__N_1595[17]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i17.GSR = "ENABLED";
    FD1P3AX comb8_i0_i18 (.D(comb8_71__N_1595[18]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i18.GSR = "ENABLED";
    FD1P3AX comb8_i0_i19 (.D(comb8_71__N_1595[19]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i19.GSR = "ENABLED";
    FD1P3AX comb8_i0_i20 (.D(comb8_71__N_1595[20]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i20.GSR = "ENABLED";
    FD1P3AX comb8_i0_i21 (.D(comb8_71__N_1595[21]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i21.GSR = "ENABLED";
    FD1P3AX comb8_i0_i22 (.D(comb8_71__N_1595[22]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i22.GSR = "ENABLED";
    FD1P3AX comb8_i0_i23 (.D(comb8_71__N_1595[23]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i23.GSR = "ENABLED";
    FD1P3AX comb8_i0_i24 (.D(comb8_71__N_1595[24]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i24.GSR = "ENABLED";
    FD1P3AX comb8_i0_i25 (.D(comb8_71__N_1595[25]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i25.GSR = "ENABLED";
    FD1P3AX comb8_i0_i26 (.D(comb8_71__N_1595[26]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i26.GSR = "ENABLED";
    FD1P3AX comb8_i0_i27 (.D(comb8_71__N_1595[27]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i27.GSR = "ENABLED";
    FD1P3AX comb8_i0_i28 (.D(comb8_71__N_1595[28]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i28.GSR = "ENABLED";
    FD1P3AX comb8_i0_i29 (.D(comb8_71__N_1595[29]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i29.GSR = "ENABLED";
    FD1P3AX comb8_i0_i30 (.D(comb8_71__N_1595[30]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i30.GSR = "ENABLED";
    FD1P3AX comb8_i0_i31 (.D(comb8_71__N_1595[31]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i31.GSR = "ENABLED";
    FD1P3AX comb8_i0_i32 (.D(comb8_71__N_1595[32]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i32.GSR = "ENABLED";
    FD1P3AX comb8_i0_i33 (.D(comb8_71__N_1595[33]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i33.GSR = "ENABLED";
    FD1P3AX comb8_i0_i34 (.D(comb8_71__N_1595[34]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i34.GSR = "ENABLED";
    FD1P3AX comb8_i0_i35 (.D(comb8_71__N_1595[35]), .SP(clk_80mhz_enable_1184), 
            .CK(clk_80mhz), .Q(comb8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i35.GSR = "ENABLED";
    FD1P3AX comb8_i0_i36 (.D(comb8_71__N_1595[36]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i36.GSR = "ENABLED";
    FD1P3AX comb8_i0_i37 (.D(comb8_71__N_1595[37]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i37.GSR = "ENABLED";
    FD1P3AX comb8_i0_i38 (.D(comb8_71__N_1595[38]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i38.GSR = "ENABLED";
    FD1P3AX comb8_i0_i39 (.D(comb8_71__N_1595[39]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i39.GSR = "ENABLED";
    FD1P3AX comb8_i0_i40 (.D(comb8_71__N_1595[40]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i40.GSR = "ENABLED";
    FD1P3AX comb8_i0_i41 (.D(comb8_71__N_1595[41]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i41.GSR = "ENABLED";
    FD1P3AX comb8_i0_i42 (.D(comb8_71__N_1595[42]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i42.GSR = "ENABLED";
    FD1P3AX comb8_i0_i43 (.D(comb8_71__N_1595[43]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i43.GSR = "ENABLED";
    FD1P3AX comb8_i0_i44 (.D(comb8_71__N_1595[44]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i44.GSR = "ENABLED";
    FD1P3AX comb8_i0_i45 (.D(comb8_71__N_1595[45]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i45.GSR = "ENABLED";
    FD1P3AX comb8_i0_i46 (.D(comb8_71__N_1595[46]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i46.GSR = "ENABLED";
    FD1P3AX comb8_i0_i47 (.D(comb8_71__N_1595[47]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i47.GSR = "ENABLED";
    FD1P3AX comb8_i0_i48 (.D(comb8_71__N_1595[48]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i48.GSR = "ENABLED";
    FD1P3AX comb8_i0_i49 (.D(comb8_71__N_1595[49]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i49.GSR = "ENABLED";
    FD1P3AX comb8_i0_i50 (.D(comb8_71__N_1595[50]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i50.GSR = "ENABLED";
    FD1P3AX comb8_i0_i51 (.D(comb8_71__N_1595[51]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i51.GSR = "ENABLED";
    FD1P3AX comb8_i0_i52 (.D(comb8_71__N_1595[52]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i52.GSR = "ENABLED";
    FD1P3AX comb8_i0_i53 (.D(comb8_71__N_1595[53]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i53.GSR = "ENABLED";
    FD1P3AX comb8_i0_i54 (.D(comb8_71__N_1595[54]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i54.GSR = "ENABLED";
    FD1P3AX comb8_i0_i55 (.D(comb8_71__N_1595[55]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i55.GSR = "ENABLED";
    FD1P3AX comb8_i0_i56 (.D(comb8_71__N_1595[56]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i56.GSR = "ENABLED";
    FD1P3AX comb8_i0_i57 (.D(comb8_71__N_1595[57]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i57.GSR = "ENABLED";
    FD1P3AX comb8_i0_i58 (.D(comb8_71__N_1595[58]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i58.GSR = "ENABLED";
    FD1P3AX comb8_i0_i59 (.D(comb8_71__N_1595[59]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i59.GSR = "ENABLED";
    FD1P3AX comb8_i0_i60 (.D(comb8_71__N_1595[60]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i60.GSR = "ENABLED";
    FD1P3AX comb8_i0_i61 (.D(comb8_71__N_1595[61]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i61.GSR = "ENABLED";
    FD1P3AX comb8_i0_i62 (.D(comb8_71__N_1595[62]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i62.GSR = "ENABLED";
    FD1P3AX comb8_i0_i63 (.D(comb8_71__N_1595[63]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i63.GSR = "ENABLED";
    FD1P3AX comb8_i0_i64 (.D(comb8_71__N_1595[64]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i64.GSR = "ENABLED";
    FD1P3AX comb8_i0_i65 (.D(comb8_71__N_1595[65]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i65.GSR = "ENABLED";
    FD1P3AX comb8_i0_i66 (.D(comb8_71__N_1595[66]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i66.GSR = "ENABLED";
    FD1P3AX comb8_i0_i67 (.D(comb8_71__N_1595[67]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i67.GSR = "ENABLED";
    FD1P3AX comb8_i0_i68 (.D(comb8_71__N_1595[68]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i68.GSR = "ENABLED";
    FD1P3AX comb8_i0_i69 (.D(comb8_71__N_1595[69]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i69.GSR = "ENABLED";
    FD1P3AX comb8_i0_i70 (.D(comb8_71__N_1595[70]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i70.GSR = "ENABLED";
    FD1P3AX comb8_i0_i71 (.D(comb8_71__N_1595[71]), .SP(clk_80mhz_enable_1234), 
            .CK(clk_80mhz), .Q(comb8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb8_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i1 (.D(comb8[1]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i2 (.D(comb8[2]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i3 (.D(comb8[3]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i4 (.D(comb8[4]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i5 (.D(comb8[5]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i6 (.D(comb8[6]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i7 (.D(comb8[7]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i8 (.D(comb8[8]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i9 (.D(comb8[9]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i10 (.D(comb8[10]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i11 (.D(comb8[11]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i12 (.D(comb8[12]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i13 (.D(comb8[13]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i14 (.D(comb8[14]), .SP(clk_80mhz_enable_1234), .CK(clk_80mhz), 
            .Q(comb_d8[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i15 (.D(comb8[15]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i16 (.D(comb8[16]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i17 (.D(comb8[17]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i18 (.D(comb8[18]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i19 (.D(comb8[19]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i20 (.D(comb8[20]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i21 (.D(comb8[21]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i22 (.D(comb8[22]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i23 (.D(comb8[23]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i24 (.D(comb8[24]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i25 (.D(comb8[25]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i26 (.D(comb8[26]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i27 (.D(comb8[27]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i28 (.D(comb8[28]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i29 (.D(comb8[29]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i30 (.D(comb8[30]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i31 (.D(comb8[31]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i32 (.D(comb8[32]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i33 (.D(comb8[33]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i34 (.D(comb8[34]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i35 (.D(comb8[35]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i36 (.D(comb8[36]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i37 (.D(comb8[37]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i38 (.D(comb8[38]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i39 (.D(comb8[39]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i40 (.D(comb8[40]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i41 (.D(comb8[41]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i42 (.D(comb8[42]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i43 (.D(comb8[43]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i44 (.D(comb8[44]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i45 (.D(comb8[45]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i46 (.D(comb8[46]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i47 (.D(comb8[47]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i48 (.D(comb8[48]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i49 (.D(comb8[49]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i50 (.D(comb8[50]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i51 (.D(comb8[51]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i52 (.D(comb8[52]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i53 (.D(comb8[53]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i54 (.D(comb8[54]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i55 (.D(comb8[55]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i56 (.D(comb8[56]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i57 (.D(comb8[57]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i58 (.D(comb8[58]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i59 (.D(comb8[59]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i60 (.D(comb8[60]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i61 (.D(comb8[61]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i62 (.D(comb8[62]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i63 (.D(comb8[63]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i64 (.D(comb8[64]), .SP(clk_80mhz_enable_1284), .CK(clk_80mhz), 
            .Q(comb_d8[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i65 (.D(comb8[65]), .SP(clk_80mhz_enable_1334), .CK(clk_80mhz), 
            .Q(comb_d8[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i66 (.D(comb8[66]), .SP(clk_80mhz_enable_1334), .CK(clk_80mhz), 
            .Q(comb_d8[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i67 (.D(comb8[67]), .SP(clk_80mhz_enable_1334), .CK(clk_80mhz), 
            .Q(comb_d8[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i68 (.D(comb8[68]), .SP(clk_80mhz_enable_1334), .CK(clk_80mhz), 
            .Q(comb_d8[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i69 (.D(comb8[69]), .SP(clk_80mhz_enable_1334), .CK(clk_80mhz), 
            .Q(comb_d8[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i70 (.D(comb8[70]), .SP(clk_80mhz_enable_1334), .CK(clk_80mhz), 
            .Q(comb_d8[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d8_i0_i71 (.D(comb8[71]), .SP(clk_80mhz_enable_1334), .CK(clk_80mhz), 
            .Q(comb_d8[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d8_i0_i71.GSR = "ENABLED";
    FD1P3AX comb9_i0_i1 (.D(comb9_71__N_1667[1]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i1.GSR = "ENABLED";
    FD1P3AX comb9_i0_i2 (.D(comb9_71__N_1667[2]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i2.GSR = "ENABLED";
    FD1P3AX comb9_i0_i3 (.D(comb9_71__N_1667[3]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i3.GSR = "ENABLED";
    FD1P3AX comb9_i0_i4 (.D(comb9_71__N_1667[4]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i4.GSR = "ENABLED";
    FD1P3AX comb9_i0_i5 (.D(comb9_71__N_1667[5]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i5.GSR = "ENABLED";
    FD1P3AX comb9_i0_i6 (.D(comb9_71__N_1667[6]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i6.GSR = "ENABLED";
    FD1P3AX comb9_i0_i7 (.D(comb9_71__N_1667[7]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i7.GSR = "ENABLED";
    FD1P3AX comb9_i0_i8 (.D(comb9_71__N_1667[8]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i8.GSR = "ENABLED";
    FD1P3AX comb9_i0_i9 (.D(comb9_71__N_1667[9]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i9.GSR = "ENABLED";
    FD1P3AX comb9_i0_i10 (.D(comb9_71__N_1667[10]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i10.GSR = "ENABLED";
    FD1P3AX comb9_i0_i11 (.D(comb9_71__N_1667[11]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i11.GSR = "ENABLED";
    FD1P3AX comb9_i0_i12 (.D(comb9_71__N_1667[12]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i12.GSR = "ENABLED";
    FD1P3AX comb9_i0_i13 (.D(comb9_71__N_1667[13]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i13.GSR = "ENABLED";
    FD1P3AX comb9_i0_i14 (.D(comb9_71__N_1667[14]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i14.GSR = "ENABLED";
    FD1P3AX comb9_i0_i15 (.D(comb9_71__N_1667[15]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i15.GSR = "ENABLED";
    FD1P3AX comb9_i0_i16 (.D(comb9_71__N_1667[16]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i16.GSR = "ENABLED";
    FD1P3AX comb9_i0_i17 (.D(comb9_71__N_1667[17]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i17.GSR = "ENABLED";
    FD1P3AX comb9_i0_i18 (.D(comb9_71__N_1667[18]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i18.GSR = "ENABLED";
    FD1P3AX comb9_i0_i19 (.D(comb9_71__N_1667[19]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i19.GSR = "ENABLED";
    FD1P3AX comb9_i0_i20 (.D(comb9_71__N_1667[20]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i20.GSR = "ENABLED";
    FD1P3AX comb9_i0_i21 (.D(comb9_71__N_1667[21]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i21.GSR = "ENABLED";
    FD1P3AX comb9_i0_i22 (.D(comb9_71__N_1667[22]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i22.GSR = "ENABLED";
    FD1P3AX comb9_i0_i23 (.D(comb9_71__N_1667[23]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i23.GSR = "ENABLED";
    FD1P3AX comb9_i0_i24 (.D(comb9_71__N_1667[24]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i24.GSR = "ENABLED";
    FD1P3AX comb9_i0_i25 (.D(comb9_71__N_1667[25]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i25.GSR = "ENABLED";
    FD1P3AX comb9_i0_i26 (.D(comb9_71__N_1667[26]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i26.GSR = "ENABLED";
    FD1P3AX comb9_i0_i27 (.D(comb9_71__N_1667[27]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i27.GSR = "ENABLED";
    FD1P3AX comb9_i0_i28 (.D(comb9_71__N_1667[28]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i28.GSR = "ENABLED";
    FD1P3AX comb9_i0_i29 (.D(comb9_71__N_1667[29]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i29.GSR = "ENABLED";
    FD1P3AX comb9_i0_i30 (.D(comb9_71__N_1667[30]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i30.GSR = "ENABLED";
    FD1P3AX comb9_i0_i31 (.D(comb9_71__N_1667[31]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i31.GSR = "ENABLED";
    FD1P3AX comb9_i0_i32 (.D(comb9_71__N_1667[32]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i32.GSR = "ENABLED";
    FD1P3AX comb9_i0_i33 (.D(comb9_71__N_1667[33]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i33.GSR = "ENABLED";
    FD1P3AX comb9_i0_i34 (.D(comb9_71__N_1667[34]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i34.GSR = "ENABLED";
    FD1P3AX comb9_i0_i35 (.D(comb9_71__N_1667[35]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i35.GSR = "ENABLED";
    FD1P3AX comb9_i0_i36 (.D(comb9_71__N_1667[36]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i36.GSR = "ENABLED";
    FD1P3AX comb9_i0_i37 (.D(comb9_71__N_1667[37]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i37.GSR = "ENABLED";
    FD1P3AX comb9_i0_i38 (.D(comb9_71__N_1667[38]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i38.GSR = "ENABLED";
    FD1P3AX comb9_i0_i39 (.D(comb9_71__N_1667[39]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i39.GSR = "ENABLED";
    FD1P3AX comb9_i0_i40 (.D(comb9_71__N_1667[40]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i40.GSR = "ENABLED";
    FD1P3AX comb9_i0_i41 (.D(comb9_71__N_1667[41]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i41.GSR = "ENABLED";
    FD1P3AX comb9_i0_i42 (.D(comb9_71__N_1667[42]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i42.GSR = "ENABLED";
    FD1P3AX comb9_i0_i43 (.D(comb9_71__N_1667[43]), .SP(clk_80mhz_enable_1334), 
            .CK(clk_80mhz), .Q(comb9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i43.GSR = "ENABLED";
    FD1P3AX comb9_i0_i44 (.D(comb9_71__N_1667[44]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i44.GSR = "ENABLED";
    FD1P3AX comb9_i0_i45 (.D(comb9_71__N_1667[45]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i45.GSR = "ENABLED";
    FD1P3AX comb9_i0_i46 (.D(comb9_71__N_1667[46]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i46.GSR = "ENABLED";
    FD1P3AX comb9_i0_i47 (.D(comb9_71__N_1667[47]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i47.GSR = "ENABLED";
    FD1P3AX comb9_i0_i48 (.D(comb9_71__N_1667[48]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i48.GSR = "ENABLED";
    FD1P3AX comb9_i0_i49 (.D(comb9_71__N_1667[49]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i49.GSR = "ENABLED";
    FD1P3AX comb9_i0_i50 (.D(comb9_71__N_1667[50]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i50.GSR = "ENABLED";
    FD1P3AX comb9_i0_i51 (.D(comb9_71__N_1667[51]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i51.GSR = "ENABLED";
    FD1P3AX comb9_i0_i52 (.D(comb9_71__N_1667[52]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i52.GSR = "ENABLED";
    FD1P3AX comb9_i0_i53 (.D(comb9_71__N_1667[53]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i53.GSR = "ENABLED";
    FD1P3AX comb9_i0_i54 (.D(comb9_71__N_1667[54]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i54.GSR = "ENABLED";
    FD1P3AX comb9_i0_i55 (.D(comb9_71__N_1667[55]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i55.GSR = "ENABLED";
    FD1P3AX comb9_i0_i56 (.D(comb9_71__N_1667[56]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i56.GSR = "ENABLED";
    FD1P3AX comb9_i0_i57 (.D(comb9_71__N_1667[57]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i57.GSR = "ENABLED";
    FD1P3AX comb9_i0_i58 (.D(comb9_71__N_1667[58]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i58.GSR = "ENABLED";
    FD1P3AX comb9_i0_i59 (.D(comb9_71__N_1667[59]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i59.GSR = "ENABLED";
    FD1P3AX comb9_i0_i60 (.D(comb9_71__N_1667[60]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i60.GSR = "ENABLED";
    FD1P3AX comb9_i0_i61 (.D(comb9_71__N_1667[61]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i61.GSR = "ENABLED";
    FD1P3AX comb9_i0_i62 (.D(comb9_71__N_1667[62]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i62.GSR = "ENABLED";
    FD1P3AX comb9_i0_i63 (.D(comb9_71__N_1667[63]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i63.GSR = "ENABLED";
    FD1P3AX comb9_i0_i64 (.D(comb9_71__N_1667[64]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i64.GSR = "ENABLED";
    FD1P3AX comb9_i0_i65 (.D(comb9_71__N_1667[65]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i65.GSR = "ENABLED";
    FD1P3AX comb9_i0_i66 (.D(comb9_71__N_1667[66]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i66.GSR = "ENABLED";
    FD1P3AX comb9_i0_i67 (.D(comb9_71__N_1667[67]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i67.GSR = "ENABLED";
    FD1P3AX comb9_i0_i68 (.D(comb9_71__N_1667[68]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i68.GSR = "ENABLED";
    FD1P3AX comb9_i0_i69 (.D(comb9_71__N_1667[69]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i69.GSR = "ENABLED";
    FD1P3AX comb9_i0_i70 (.D(comb9_71__N_1667[70]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i70.GSR = "ENABLED";
    FD1P3AX comb9_i0_i71 (.D(comb9_71__N_1667[71]), .SP(clk_80mhz_enable_1384), 
            .CK(clk_80mhz), .Q(comb9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb9_i0_i71.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i1 (.D(comb9[1]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i1.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i2 (.D(comb9[2]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i2.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i3 (.D(comb9[3]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i3.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i4 (.D(comb9[4]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i4.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i5 (.D(comb9[5]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i5.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i6 (.D(comb9[6]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i6.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i7 (.D(comb9[7]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i7.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i8 (.D(comb9[8]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i8.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i9 (.D(comb9[9]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i9.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i10 (.D(comb9[10]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i10.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i11 (.D(comb9[11]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i11.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i12 (.D(comb9[12]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i12.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i13 (.D(comb9[13]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i13.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i14 (.D(comb9[14]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i14.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i15 (.D(comb9[15]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i15.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i16 (.D(comb9[16]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i16.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i17 (.D(comb9[17]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i17.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i18 (.D(comb9[18]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i18.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i19 (.D(comb9[19]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i19.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i20 (.D(comb9[20]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i20.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i21 (.D(comb9[21]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i21.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i22 (.D(comb9[22]), .SP(clk_80mhz_enable_1384), .CK(clk_80mhz), 
            .Q(comb_d9[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i22.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i23 (.D(comb9[23]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i23.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i24 (.D(comb9[24]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i24.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i25 (.D(comb9[25]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i25.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i26 (.D(comb9[26]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i26.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i27 (.D(comb9[27]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i27.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i28 (.D(comb9[28]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i28.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i29 (.D(comb9[29]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i29.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i30 (.D(comb9[30]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i30.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i31 (.D(comb9[31]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i31.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i32 (.D(comb9[32]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i32.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i33 (.D(comb9[33]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i33.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i34 (.D(comb9[34]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i34.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i35 (.D(comb9[35]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i35.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i36 (.D(comb9[36]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i36.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i37 (.D(comb9[37]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i37.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i38 (.D(comb9[38]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i38.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i39 (.D(comb9[39]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i39.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i40 (.D(comb9[40]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i40.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i41 (.D(comb9[41]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i41.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i42 (.D(comb9[42]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i42.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i43 (.D(comb9[43]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i43.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i44 (.D(comb9[44]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i44.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i45 (.D(comb9[45]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i45.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i46 (.D(comb9[46]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i46.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i47 (.D(comb9[47]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i47.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i48 (.D(comb9[48]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i48.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i49 (.D(comb9[49]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i49.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i50 (.D(comb9[50]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i50.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i51 (.D(comb9[51]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i51.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i52 (.D(comb9[52]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i52.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i53 (.D(comb9[53]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i53.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i54 (.D(comb9[54]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i54.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i55 (.D(comb9[55]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i55.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i56 (.D(comb9[56]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i56.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i57 (.D(comb9[57]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i57.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i58 (.D(comb9[58]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i58.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i59 (.D(comb9[59]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i59.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i60 (.D(comb9[60]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i60.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i61 (.D(comb9[61]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i61.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i62 (.D(comb9[62]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i62.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i63 (.D(comb9[63]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i63.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i64 (.D(comb9[64]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i64.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i65 (.D(comb9[65]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i65.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i66 (.D(comb9[66]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i66.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i67 (.D(comb9[67]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i67.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i68 (.D(comb9[68]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i68.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i69 (.D(comb9[69]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i69.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i70 (.D(comb9[70]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i70.GSR = "ENABLED";
    FD1P3AX comb_d9_i0_i71 (.D(comb9[71]), .SP(clk_80mhz_enable_1434), .CK(clk_80mhz), 
            .Q(comb_d9[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb_d9_i0_i71.GSR = "ENABLED";
    FD1P3AX comb10__i2 (.D(comb10_71__N_1739[57]), .SP(clk_80mhz_enable_1434), 
            .CK(clk_80mhz), .Q(comb10[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i2.GSR = "ENABLED";
    FD1P3AX comb10__i3 (.D(comb10_71__N_1739[58]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(comb10[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i3.GSR = "ENABLED";
    FD1P3AX comb10__i4 (.D(comb10_71__N_1739[59]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i4.GSR = "ENABLED";
    FD1P3AX comb10__i5 (.D(comb10_71__N_1739[60]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i5.GSR = "ENABLED";
    FD1P3AX comb10__i6 (.D(comb10_71__N_1739[61]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[61] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i6.GSR = "ENABLED";
    FD1P3AX comb10__i7 (.D(comb10_71__N_1739[62]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[62] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i7.GSR = "ENABLED";
    FD1P3AX comb10__i8 (.D(comb10_71__N_1739[63]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[63] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i8.GSR = "ENABLED";
    FD1P3AX comb10__i9 (.D(comb10_71__N_1739[64]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[64] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i9.GSR = "ENABLED";
    FD1P3AX comb10__i10 (.D(comb10_71__N_1739[65]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[65] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i10.GSR = "ENABLED";
    FD1P3AX comb10__i11 (.D(comb10_71__N_1739[66]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[66] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i11.GSR = "ENABLED";
    FD1P3AX comb10__i12 (.D(comb10_71__N_1739[67]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[67] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i12.GSR = "ENABLED";
    FD1P3AX comb10__i13 (.D(comb10_71__N_1739[68]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[68] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i13.GSR = "ENABLED";
    FD1P3AX comb10__i14 (.D(comb10_71__N_1739[69]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[69] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i14.GSR = "ENABLED";
    FD1P3AX comb10__i15 (.D(comb10_71__N_1739[70]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[70] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i15.GSR = "ENABLED";
    FD1P3AX comb10__i16 (.D(comb10_71__N_1739[71]), .SP(valid_comb), .CK(clk_80mhz), 
            .Q(\comb10[71] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam comb10__i16.GSR = "ENABLED";
    FD1P3AX data_out_i0_i1 (.D(data_out_11__N_1811[1]), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(cic_cosine_out[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i1.GSR = "ENABLED";
    FD1P3AX data_out_i0_i2 (.D(\data_out_11__N_1811[2] ), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(cic_cosine_out[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i2.GSR = "ENABLED";
    FD1P3AX data_out_i0_i3 (.D(\data_out_11__N_1811[3] ), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(cic_cosine_out[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i3.GSR = "ENABLED";
    FD1P3AX data_out_i0_i4 (.D(\data_out_11__N_1811[4] ), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(cic_cosine_out[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i4.GSR = "ENABLED";
    FD1P3AX data_out_i0_i5 (.D(\data_out_11__N_1811[5] ), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(cic_cosine_out[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i5.GSR = "ENABLED";
    FD1P3AX data_out_i0_i6 (.D(\data_out_11__N_1811[6] ), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(cic_cosine_out[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i6.GSR = "ENABLED";
    FD1P3AX data_out_i0_i7 (.D(\data_out_11__N_1811[7] ), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(cic_cosine_out[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i7.GSR = "ENABLED";
    FD1P3AX data_out_i0_i8 (.D(\data_out_11__N_1811[8] ), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(cic_cosine_out[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i8.GSR = "ENABLED";
    FD1P3AX data_out_i0_i9 (.D(\data_out_11__N_1811[9] ), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(cic_cosine_out[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i9.GSR = "ENABLED";
    FD1P3AX data_out_i0_i10 (.D(\data_out_11__N_1811[10] ), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(cic_cosine_out[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i10.GSR = "ENABLED";
    FD1P3AX data_out_i0_i11 (.D(\data_out_11__N_1811[11] ), .SP(valid_comb), 
            .CK(clk_80mhz), .Q(cic_cosine_out[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(89[10] 108[6])
    defparam data_out_i0_i11.GSR = "ENABLED";
    FD1S3AX integrator1_i1 (.D(integrator1_71__N_418[1]), .CK(clk_80mhz), 
            .Q(integrator1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i1.GSR = "ENABLED";
    FD1S3AX integrator1_i2 (.D(integrator1_71__N_418[2]), .CK(clk_80mhz), 
            .Q(integrator1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i2.GSR = "ENABLED";
    FD1S3AX integrator1_i3 (.D(integrator1_71__N_418[3]), .CK(clk_80mhz), 
            .Q(integrator1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i3.GSR = "ENABLED";
    FD1S3AX integrator1_i4 (.D(integrator1_71__N_418[4]), .CK(clk_80mhz), 
            .Q(integrator1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i4.GSR = "ENABLED";
    FD1S3AX integrator1_i5 (.D(integrator1_71__N_418[5]), .CK(clk_80mhz), 
            .Q(integrator1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i5.GSR = "ENABLED";
    FD1S3AX integrator1_i6 (.D(integrator1_71__N_418[6]), .CK(clk_80mhz), 
            .Q(integrator1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i6.GSR = "ENABLED";
    FD1S3AX integrator1_i7 (.D(integrator1_71__N_418[7]), .CK(clk_80mhz), 
            .Q(integrator1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i7.GSR = "ENABLED";
    FD1S3AX integrator1_i8 (.D(integrator1_71__N_418[8]), .CK(clk_80mhz), 
            .Q(integrator1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i8.GSR = "ENABLED";
    FD1S3AX integrator1_i9 (.D(integrator1_71__N_418[9]), .CK(clk_80mhz), 
            .Q(integrator1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i9.GSR = "ENABLED";
    FD1S3AX integrator1_i10 (.D(integrator1_71__N_418[10]), .CK(clk_80mhz), 
            .Q(integrator1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i10.GSR = "ENABLED";
    FD1S3AX integrator1_i11 (.D(integrator1_71__N_418[11]), .CK(clk_80mhz), 
            .Q(integrator1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i11.GSR = "ENABLED";
    FD1S3AX integrator1_i12 (.D(integrator1_71__N_418[12]), .CK(clk_80mhz), 
            .Q(integrator1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i12.GSR = "ENABLED";
    FD1S3AX integrator1_i13 (.D(integrator1_71__N_418[13]), .CK(clk_80mhz), 
            .Q(integrator1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i13.GSR = "ENABLED";
    FD1S3AX integrator1_i14 (.D(integrator1_71__N_418[14]), .CK(clk_80mhz), 
            .Q(integrator1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i14.GSR = "ENABLED";
    FD1S3AX integrator1_i15 (.D(integrator1_71__N_418[15]), .CK(clk_80mhz), 
            .Q(integrator1[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i15.GSR = "ENABLED";
    FD1S3AX integrator1_i16 (.D(integrator1_71__N_418[16]), .CK(clk_80mhz), 
            .Q(integrator1[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i16.GSR = "ENABLED";
    FD1S3AX integrator1_i17 (.D(integrator1_71__N_418[17]), .CK(clk_80mhz), 
            .Q(integrator1[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i17.GSR = "ENABLED";
    FD1S3AX integrator1_i18 (.D(integrator1_71__N_418[18]), .CK(clk_80mhz), 
            .Q(integrator1[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i18.GSR = "ENABLED";
    FD1S3AX integrator1_i19 (.D(integrator1_71__N_418[19]), .CK(clk_80mhz), 
            .Q(integrator1[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i19.GSR = "ENABLED";
    FD1S3AX integrator1_i20 (.D(integrator1_71__N_418[20]), .CK(clk_80mhz), 
            .Q(integrator1[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i20.GSR = "ENABLED";
    FD1S3AX integrator1_i21 (.D(integrator1_71__N_418[21]), .CK(clk_80mhz), 
            .Q(integrator1[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i21.GSR = "ENABLED";
    FD1S3AX integrator1_i22 (.D(integrator1_71__N_418[22]), .CK(clk_80mhz), 
            .Q(integrator1[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i22.GSR = "ENABLED";
    FD1S3AX integrator1_i23 (.D(integrator1_71__N_418[23]), .CK(clk_80mhz), 
            .Q(integrator1[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i23.GSR = "ENABLED";
    FD1S3AX integrator1_i24 (.D(integrator1_71__N_418[24]), .CK(clk_80mhz), 
            .Q(integrator1[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i24.GSR = "ENABLED";
    FD1S3AX integrator1_i25 (.D(integrator1_71__N_418[25]), .CK(clk_80mhz), 
            .Q(integrator1[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i25.GSR = "ENABLED";
    FD1S3AX integrator1_i26 (.D(integrator1_71__N_418[26]), .CK(clk_80mhz), 
            .Q(integrator1[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i26.GSR = "ENABLED";
    FD1S3AX integrator1_i27 (.D(integrator1_71__N_418[27]), .CK(clk_80mhz), 
            .Q(integrator1[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i27.GSR = "ENABLED";
    FD1S3AX integrator1_i28 (.D(integrator1_71__N_418[28]), .CK(clk_80mhz), 
            .Q(integrator1[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i28.GSR = "ENABLED";
    FD1S3AX integrator1_i29 (.D(integrator1_71__N_418[29]), .CK(clk_80mhz), 
            .Q(integrator1[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i29.GSR = "ENABLED";
    FD1S3AX integrator1_i30 (.D(integrator1_71__N_418[30]), .CK(clk_80mhz), 
            .Q(integrator1[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i30.GSR = "ENABLED";
    FD1S3AX integrator1_i31 (.D(integrator1_71__N_418[31]), .CK(clk_80mhz), 
            .Q(integrator1[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i31.GSR = "ENABLED";
    FD1S3AX integrator1_i32 (.D(integrator1_71__N_418[32]), .CK(clk_80mhz), 
            .Q(integrator1[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i32.GSR = "ENABLED";
    FD1S3AX integrator1_i33 (.D(integrator1_71__N_418[33]), .CK(clk_80mhz), 
            .Q(integrator1[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i33.GSR = "ENABLED";
    FD1S3AX integrator1_i34 (.D(integrator1_71__N_418[34]), .CK(clk_80mhz), 
            .Q(integrator1[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i34.GSR = "ENABLED";
    FD1S3AX integrator1_i35 (.D(integrator1_71__N_418[35]), .CK(clk_80mhz), 
            .Q(integrator1[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i35.GSR = "ENABLED";
    FD1S3AX integrator1_i36 (.D(integrator1_71__N_418[36]), .CK(clk_80mhz), 
            .Q(integrator1[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i36.GSR = "ENABLED";
    FD1S3AX integrator1_i37 (.D(integrator1_71__N_418[37]), .CK(clk_80mhz), 
            .Q(integrator1[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i37.GSR = "ENABLED";
    FD1S3AX integrator1_i38 (.D(integrator1_71__N_418[38]), .CK(clk_80mhz), 
            .Q(integrator1[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i38.GSR = "ENABLED";
    FD1S3AX integrator1_i39 (.D(integrator1_71__N_418[39]), .CK(clk_80mhz), 
            .Q(integrator1[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i39.GSR = "ENABLED";
    FD1S3AX integrator1_i40 (.D(integrator1_71__N_418[40]), .CK(clk_80mhz), 
            .Q(integrator1[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i40.GSR = "ENABLED";
    FD1S3AX integrator1_i41 (.D(integrator1_71__N_418[41]), .CK(clk_80mhz), 
            .Q(integrator1[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i41.GSR = "ENABLED";
    FD1S3AX integrator1_i42 (.D(integrator1_71__N_418[42]), .CK(clk_80mhz), 
            .Q(integrator1[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i42.GSR = "ENABLED";
    FD1S3AX integrator1_i43 (.D(integrator1_71__N_418[43]), .CK(clk_80mhz), 
            .Q(integrator1[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i43.GSR = "ENABLED";
    FD1S3AX integrator1_i44 (.D(integrator1_71__N_418[44]), .CK(clk_80mhz), 
            .Q(integrator1[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i44.GSR = "ENABLED";
    FD1S3AX integrator1_i45 (.D(integrator1_71__N_418[45]), .CK(clk_80mhz), 
            .Q(integrator1[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i45.GSR = "ENABLED";
    FD1S3AX integrator1_i46 (.D(integrator1_71__N_418[46]), .CK(clk_80mhz), 
            .Q(integrator1[46])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i46.GSR = "ENABLED";
    FD1S3AX integrator1_i47 (.D(integrator1_71__N_418[47]), .CK(clk_80mhz), 
            .Q(integrator1[47])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i47.GSR = "ENABLED";
    FD1S3AX integrator1_i48 (.D(integrator1_71__N_418[48]), .CK(clk_80mhz), 
            .Q(integrator1[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i48.GSR = "ENABLED";
    FD1S3AX integrator1_i49 (.D(integrator1_71__N_418[49]), .CK(clk_80mhz), 
            .Q(integrator1[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i49.GSR = "ENABLED";
    FD1S3AX integrator1_i50 (.D(integrator1_71__N_418[50]), .CK(clk_80mhz), 
            .Q(integrator1[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i50.GSR = "ENABLED";
    FD1S3AX integrator1_i51 (.D(integrator1_71__N_418[51]), .CK(clk_80mhz), 
            .Q(integrator1[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i51.GSR = "ENABLED";
    FD1S3AX integrator1_i52 (.D(integrator1_71__N_418[52]), .CK(clk_80mhz), 
            .Q(integrator1[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i52.GSR = "ENABLED";
    FD1S3AX integrator1_i53 (.D(integrator1_71__N_418[53]), .CK(clk_80mhz), 
            .Q(integrator1[53])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i53.GSR = "ENABLED";
    FD1S3AX integrator1_i54 (.D(integrator1_71__N_418[54]), .CK(clk_80mhz), 
            .Q(integrator1[54])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i54.GSR = "ENABLED";
    FD1S3AX integrator1_i55 (.D(integrator1_71__N_418[55]), .CK(clk_80mhz), 
            .Q(integrator1[55])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i55.GSR = "ENABLED";
    FD1S3AX integrator1_i56 (.D(integrator1_71__N_418[56]), .CK(clk_80mhz), 
            .Q(integrator1[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i56.GSR = "ENABLED";
    FD1S3AX integrator1_i57 (.D(integrator1_71__N_418[57]), .CK(clk_80mhz), 
            .Q(integrator1[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i57.GSR = "ENABLED";
    FD1S3AX integrator1_i58 (.D(integrator1_71__N_418[58]), .CK(clk_80mhz), 
            .Q(integrator1[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i58.GSR = "ENABLED";
    FD1S3AX integrator1_i59 (.D(integrator1_71__N_418[59]), .CK(clk_80mhz), 
            .Q(integrator1[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i59.GSR = "ENABLED";
    FD1S3AX integrator1_i60 (.D(integrator1_71__N_418[60]), .CK(clk_80mhz), 
            .Q(integrator1[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i60.GSR = "ENABLED";
    FD1S3AX integrator1_i61 (.D(integrator1_71__N_418[61]), .CK(clk_80mhz), 
            .Q(integrator1[61])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i61.GSR = "ENABLED";
    FD1S3AX integrator1_i62 (.D(integrator1_71__N_418[62]), .CK(clk_80mhz), 
            .Q(integrator1[62])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i62.GSR = "ENABLED";
    FD1S3AX integrator1_i63 (.D(integrator1_71__N_418[63]), .CK(clk_80mhz), 
            .Q(integrator1[63])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i63.GSR = "ENABLED";
    FD1S3AX integrator1_i64 (.D(integrator1_71__N_418[64]), .CK(clk_80mhz), 
            .Q(integrator1[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i64.GSR = "ENABLED";
    FD1S3AX integrator1_i65 (.D(integrator1_71__N_418[65]), .CK(clk_80mhz), 
            .Q(integrator1[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i65.GSR = "ENABLED";
    FD1S3AX integrator1_i66 (.D(integrator1_71__N_418[66]), .CK(clk_80mhz), 
            .Q(integrator1[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i66.GSR = "ENABLED";
    FD1S3AX integrator1_i67 (.D(integrator1_71__N_418[67]), .CK(clk_80mhz), 
            .Q(integrator1[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i67.GSR = "ENABLED";
    FD1S3AX integrator1_i68 (.D(integrator1_71__N_418[68]), .CK(clk_80mhz), 
            .Q(integrator1[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i68.GSR = "ENABLED";
    FD1S3AX integrator1_i69 (.D(integrator1_71__N_418[69]), .CK(clk_80mhz), 
            .Q(integrator1[69])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i69.GSR = "ENABLED";
    FD1S3AX integrator1_i70 (.D(integrator1_71__N_418[70]), .CK(clk_80mhz), 
            .Q(integrator1[70])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i70.GSR = "ENABLED";
    FD1S3AX integrator1_i71 (.D(integrator1_71__N_418[71]), .CK(clk_80mhz), 
            .Q(integrator1[71])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam integrator1_i71.GSR = "ENABLED";
    LUT4 sub_27_inv_0_i41_1_lut (.A(comb_d7[40]), .Z(n33_adj_85)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i42_1_lut (.A(comb_d7[41]), .Z(n32_adj_86)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i39_1_lut (.A(comb_d7[38]), .Z(n35_adj_87)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i40_1_lut (.A(comb_d7[39]), .Z(n34_adj_88)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i37_1_lut (.A(comb_d7[36]), .Z(n37_adj_89)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_27_inv_0_i38_1_lut (.A(comb_d7[37]), .Z(n36_adj_90)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(99[28:43])
    defparam sub_27_inv_0_i38_1_lut.init = 16'h5555;
    LUT4 mux_874_i2_3_lut (.A(n118), .B(n120), .C(cout), .Z(comb10_71__N_1739[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i2_3_lut.init = 16'hcaca;
    LUT4 mux_874_i3_3_lut (.A(n115), .B(n117), .C(cout), .Z(comb10_71__N_1739[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i3_3_lut.init = 16'hcaca;
    LUT4 mux_874_i4_3_lut (.A(n112), .B(n114), .C(cout), .Z(comb10_71__N_1739[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i4_3_lut.init = 16'hcaca;
    LUT4 mux_874_i5_3_lut (.A(n109), .B(n111), .C(cout), .Z(comb10_71__N_1739[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i5_3_lut.init = 16'hcaca;
    LUT4 mux_874_i6_3_lut (.A(n106), .B(n108), .C(cout), .Z(comb10_71__N_1739[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i6_3_lut.init = 16'hcaca;
    LUT4 mux_874_i7_3_lut (.A(n103), .B(n105), .C(cout), .Z(comb10_71__N_1739[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i7_3_lut.init = 16'hcaca;
    LUT4 mux_874_i8_3_lut (.A(n100), .B(n102), .C(cout), .Z(comb10_71__N_1739[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i8_3_lut.init = 16'hcaca;
    LUT4 mux_874_i9_3_lut (.A(n97), .B(n99), .C(cout), .Z(comb10_71__N_1739[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i9_3_lut.init = 16'hcaca;
    LUT4 mux_874_i10_3_lut (.A(n94), .B(n96), .C(cout), .Z(comb10_71__N_1739[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i10_3_lut.init = 16'hcaca;
    FD1S3IX count__i2 (.D(n67[2]), .CK(clk_80mhz), .CD(n11961), .Q(count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i2.GSR = "ENABLED";
    FD1S3IX count__i3 (.D(n67[3]), .CK(clk_80mhz), .CD(n11961), .Q(count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i3.GSR = "ENABLED";
    FD1S3IX count__i4 (.D(n67[4]), .CK(clk_80mhz), .CD(n11961), .Q(count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i4.GSR = "ENABLED";
    FD1S3IX count__i5 (.D(n67[5]), .CK(clk_80mhz), .CD(n11961), .Q(count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i5.GSR = "ENABLED";
    FD1S3IX count__i6 (.D(n67[6]), .CK(clk_80mhz), .CD(n11961), .Q(count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i6.GSR = "ENABLED";
    FD1S3IX count__i7 (.D(n67[7]), .CK(clk_80mhz), .CD(n11961), .Q(count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i7.GSR = "ENABLED";
    FD1S3IX count__i8 (.D(n67[8]), .CK(clk_80mhz), .CD(n11961), .Q(count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i8.GSR = "ENABLED";
    FD1S3IX count__i9 (.D(n67[9]), .CK(clk_80mhz), .CD(n11961), .Q(count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i9.GSR = "ENABLED";
    FD1S3IX count__i10 (.D(n67[10]), .CK(clk_80mhz), .CD(n11961), .Q(count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i10.GSR = "ENABLED";
    FD1S3IX count__i11 (.D(count_11__N_1438[11]), .CK(clk_80mhz), .CD(count_11__N_1450), 
            .Q(count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam count__i11.GSR = "ENABLED";
    LUT4 mux_874_i11_3_lut (.A(n91), .B(n93), .C(cout), .Z(comb10_71__N_1739[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i11_3_lut.init = 16'hcaca;
    LUT4 mux_874_i12_3_lut (.A(n88), .B(n90), .C(cout), .Z(comb10_71__N_1739[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i12_3_lut.init = 16'hcaca;
    LUT4 mux_874_i13_3_lut (.A(n85), .B(n87), .C(cout), .Z(comb10_71__N_1739[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i13_3_lut.init = 16'hcaca;
    LUT4 mux_874_i14_3_lut (.A(n82), .B(n84), .C(cout), .Z(comb10_71__N_1739[69])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i14_3_lut.init = 16'hcaca;
    LUT4 mux_874_i15_3_lut (.A(n79), .B(n81), .C(cout), .Z(comb10_71__N_1739[70])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i15_3_lut.init = 16'hcaca;
    LUT4 mux_874_i16_3_lut (.A(n76), .B(n78), .C(cout), .Z(comb10_71__N_1739[71])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(103[28:43])
    defparam mux_874_i16_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n16507), .B(count[6]), .C(n16491), .D(count[8]), 
         .Z(count_11__N_1450)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_153 (.A(count[2]), .B(n16503), .C(n16489), .D(count[4]), 
         .Z(n16507)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_153.init = 16'h8000;
    LUT4 i1_2_lut (.A(count[11]), .B(count[9]), .Z(n16491)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_154 (.A(count[1]), .B(count[3]), .C(count[0]), .D(count[10]), 
         .Z(n16503)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_154.init = 16'h8000;
    LUT4 i1_2_lut_adj_155 (.A(count[7]), .B(count[5]), .Z(n16489)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_155.init = 16'h8888;
    LUT4 shift_right_31_i62_3_lut (.A(\comb10[61] ), .B(\comb10[62] ), .C(\cic_gain[0] ), 
         .Z(n62)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i62_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i63_3_lut (.A(\comb10[62] ), .B(\comb10[63] ), .C(\cic_gain[0] ), 
         .Z(n63)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i63_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i64_3_lut (.A(\comb10[63] ), .B(\comb10[64] ), .C(\cic_gain[0] ), 
         .Z(n64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i64_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i65_3_lut (.A(\comb10[64] ), .B(\comb10[65] ), .C(\cic_gain[0] ), 
         .Z(n65)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i65_3_lut.init = 16'hcaca;
    LUT4 shift_right_31_i66_3_lut (.A(\comb10[65] ), .B(\comb10[66] ), .C(\cic_gain[0] ), 
         .Z(n66)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i66_3_lut.init = 16'hcaca;
    LUT4 i5751_2_lut (.A(n23_adj_2474), .B(n17319), .Z(n11961)) /* synthesis lut_function=((B)+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam i5751_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_adj_156 (.A(count[11]), .B(n16545), .C(n16529), .D(n16537), 
         .Z(n23_adj_2474)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(78[18:48])
    defparam i1_4_lut_adj_156.init = 16'hfffd;
    LUT4 i1_4_lut_adj_157 (.A(count[6]), .B(n16541), .C(count[7]), .D(count[4]), 
         .Z(n16545)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(78[18:48])
    defparam i1_4_lut_adj_157.init = 16'hfffe;
    LUT4 i1_2_lut_adj_158 (.A(count[2]), .B(count[5]), .Z(n16529)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(78[18:48])
    defparam i1_2_lut_adj_158.init = 16'heeee;
    LUT4 i1_2_lut_adj_159 (.A(count[9]), .B(count[10]), .Z(n16537)) /* synthesis lut_function=(A+(B)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(78[18:48])
    defparam i1_2_lut_adj_159.init = 16'heeee;
    LUT4 i1_4_lut_adj_160 (.A(count[1]), .B(count[3]), .C(count[0]), .D(count[8]), 
         .Z(n16541)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(78[18:48])
    defparam i1_4_lut_adj_160.init = 16'hfffe;
    LUT4 i1_4_lut_rep_402 (.A(n16507), .B(count[6]), .C(n16491), .D(count[8]), 
         .Z(n17319)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_rep_402.init = 16'h8000;
    LUT4 sub_28_inv_0_i57_1_lut (.A(comb_d8[56]), .Z(n17_adj_91)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i57_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i58_1_lut (.A(comb_d8[57]), .Z(n16_adj_92)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i58_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i55_1_lut (.A(comb_d8[54]), .Z(n19_adj_93)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i55_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i56_1_lut (.A(comb_d8[55]), .Z(n18_adj_94)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i56_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i53_1_lut (.A(comb_d8[52]), .Z(n21_adj_95)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i53_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i54_1_lut (.A(comb_d8[53]), .Z(n20_adj_96)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i54_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i51_1_lut (.A(comb_d8[50]), .Z(n23_adj_97)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i51_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i52_1_lut (.A(comb_d8[51]), .Z(n22_adj_98)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i52_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i49_1_lut (.A(comb_d8[48]), .Z(n25_adj_99)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i49_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i50_1_lut (.A(comb_d8[49]), .Z(n24_adj_100)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i50_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i47_1_lut (.A(comb_d8[46]), .Z(n27_adj_101)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i47_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i48_1_lut (.A(comb_d8[47]), .Z(n26_adj_102)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i48_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i45_1_lut (.A(comb_d8[44]), .Z(n29_adj_103)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i45_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i46_1_lut (.A(comb_d8[45]), .Z(n28_adj_104)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i46_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i43_1_lut (.A(comb_d8[42]), .Z(n31_adj_105)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i43_1_lut.init = 16'h5555;
    LUT4 shift_right_31_i61_rep_185_3_lut (.A(\comb10[60] ), .B(\comb10[61] ), 
         .C(\cic_gain[0] ), .Z(n16607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(106[28:76])
    defparam shift_right_31_i61_rep_185_3_lut.init = 16'hcaca;
    LUT4 sub_28_inv_0_i44_1_lut (.A(comb_d8[43]), .Z(n30_adj_106)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i44_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i41_1_lut (.A(comb_d8[40]), .Z(n33_adj_107)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i41_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i42_1_lut (.A(comb_d8[41]), .Z(n32_adj_108)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i42_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i39_1_lut (.A(comb_d8[38]), .Z(n35_adj_109)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i39_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i40_1_lut (.A(comb_d8[39]), .Z(n34_adj_110)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i40_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i37_1_lut (.A(comb_d8[36]), .Z(n37_adj_111)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i37_1_lut.init = 16'h5555;
    LUT4 sub_28_inv_0_i38_1_lut (.A(comb_d8[37]), .Z(n36_adj_112)) /* synthesis lut_function=(!(A)) */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(101[28:43])
    defparam sub_28_inv_0_i38_1_lut.init = 16'h5555;
    PFUMX i5842 (.BLUT(n17209), .ALUT(n17210), .C0(\cic_gain[0] ), .Z(data_out_11__N_1811[1]));
    LUT4 i1_4_lut_rep_403 (.A(n16507), .B(count[6]), .C(n16491), .D(count[8]), 
         .Z(clk_80mhz_enable_794)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_rep_403.init = 16'h8000;
    FD1S3AX valid_comb_66_rep_417 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1434)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_417.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_416 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1384)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_416.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_415 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1334)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_415.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_414 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1284)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_414.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_413 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1234)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_413.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_412 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1184)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_412.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_411 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1134)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_411.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_410 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1084)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_410.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_409 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_1034)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_409.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_408 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_984)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_408.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_407 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_934)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_407.GSR = "ENABLED";
    FD1S3AX valid_comb_66_rep_406 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_884)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_406.GSR = "ENABLED";
    PFUMX i5816 (.BLUT(n17169), .ALUT(n17170), .C0(\cic_gain[0] ), .Z(data_out_11__N_1811[0]));
    FD1S3AX valid_comb_66_rep_405 (.D(clk_80mhz_enable_794), .CK(clk_80mhz), 
            .Q(clk_80mhz_enable_834)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=171, LSE_RLINE=177 */ ;   // /home/user/SDR-HLS/1.RTLImplementation/3.lattice/Version2/impl1/source/CIC.v(65[10] 86[6])
    defparam valid_comb_66_rep_405.GSR = "ENABLED";
    
endmodule
