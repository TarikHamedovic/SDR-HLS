module simpleSineO(
    clk,
    rst,
    sample_clock_ce,
    phase_inc_carrGen,
    sinewave
);

input clk;
input wire rst;
input wire sample_clock_ce;
input reg signed [63:0] phase_inc_carrGen;
output reg signed[11:0] sinewave;

reg [63:0]	phase = 0;

always @(posedge clk or posedge rst) begin
    if (rst)
        phase <= 0;
    else if (sample_clock_ce)
        phase <= phase + phase_inc_carrGen;
end

always @(posedge clk) begin
	if (sample_clock_ce) begin
        case(phase[63:56])
        8'h00: sinewave <= 12'h019;
        8'h01: sinewave <= 12'h04B;
        8'h02: sinewave <= 12'h07D;
        8'h03: sinewave <= 12'h0AF;
        8'h04: sinewave <= 12'h0E1;
        8'h05: sinewave <= 12'h113;
        8'h06: sinewave <= 12'h145;
        8'h07: sinewave <= 12'h176;
        8'h08: sinewave <= 12'h1A7;
        8'h09: sinewave <= 12'h1D8;
        8'h0A: sinewave <= 12'h209;
        8'h0B: sinewave <= 12'h23A;
        8'h0C: sinewave <= 12'h26A;
        8'h0D: sinewave <= 12'h299;
        8'h0E: sinewave <= 12'h2C9;
        8'h0F: sinewave <= 12'h2F8;
        8'h10: sinewave <= 12'h326;
        8'h11: sinewave <= 12'h354;
        8'h12: sinewave <= 12'h381;
        8'h13: sinewave <= 12'h3AE;
        8'h14: sinewave <= 12'h3DB;
        8'h15: sinewave <= 12'h406;
        8'h16: sinewave <= 12'h431;
        8'h17: sinewave <= 12'h45C;
        8'h18: sinewave <= 12'h486;
        8'h19: sinewave <= 12'h4AF;
        8'h1A: sinewave <= 12'h4D7;
        8'h1B: sinewave <= 12'h4FF;
        8'h1C: sinewave <= 12'h525;
        8'h1D: sinewave <= 12'h54B;
        8'h1E: sinewave <= 12'h571;
        8'h1F: sinewave <= 12'h595;
        8'h20: sinewave <= 12'h5B9;
        8'h21: sinewave <= 12'h5DB;
        8'h22: sinewave <= 12'h5FD;
        8'h23: sinewave <= 12'h61E;
        8'h24: sinewave <= 12'h63E;
        8'h25: sinewave <= 12'h65D;
        8'h26: sinewave <= 12'h67B;
        8'h27: sinewave <= 12'h697;
        8'h28: sinewave <= 12'h6B3;
        8'h29: sinewave <= 12'h6CE;
        8'h2A: sinewave <= 12'h6E8;
        8'h2B: sinewave <= 12'h701;
        8'h2C: sinewave <= 12'h718;
        8'h2D: sinewave <= 12'h72F;
        8'h2E: sinewave <= 12'h745;
        8'h2F: sinewave <= 12'h759;
        8'h30: sinewave <= 12'h76C;
        8'h31: sinewave <= 12'h77E;
        8'h32: sinewave <= 12'h78F;
        8'h33: sinewave <= 12'h79F;
        8'h34: sinewave <= 12'h7AE;
        8'h35: sinewave <= 12'h7BB;
        8'h36: sinewave <= 12'h7C7;
        8'h37: sinewave <= 12'h7D2;
        8'h38: sinewave <= 12'h7DC;
        8'h39: sinewave <= 12'h7E5;
        8'h3A: sinewave <= 12'h7EC;
        8'h3B: sinewave <= 12'h7F2;
        8'h3C: sinewave <= 12'h7F7;
        8'h3D: sinewave <= 12'h7FB;
        8'h3E: sinewave <= 12'h7FD;
        8'h3F: sinewave <= 12'h7FE;
        8'h40: sinewave <= 12'h7FE;
        8'h41: sinewave <= 12'h7FD;
        8'h42: sinewave <= 12'h7FB;
        8'h43: sinewave <= 12'h7F7;
        8'h44: sinewave <= 12'h7F2;
        8'h45: sinewave <= 12'h7EC;
        8'h46: sinewave <= 12'h7E5;
        8'h47: sinewave <= 12'h7DC;
        8'h48: sinewave <= 12'h7D2;
        8'h49: sinewave <= 12'h7C7;
        8'h4A: sinewave <= 12'h7BB;
        8'h4B: sinewave <= 12'h7AE;
        8'h4C: sinewave <= 12'h79F;
        8'h4D: sinewave <= 12'h78F;
        8'h4E: sinewave <= 12'h77E;
        8'h4F: sinewave <= 12'h76C;
        8'h50: sinewave <= 12'h759;
        8'h51: sinewave <= 12'h745;
        8'h52: sinewave <= 12'h72F;
        8'h53: sinewave <= 12'h718;
        8'h54: sinewave <= 12'h701;
        8'h55: sinewave <= 12'h6E8;
        8'h56: sinewave <= 12'h6CE;
        8'h57: sinewave <= 12'h6B3;
        8'h58: sinewave <= 12'h697;
        8'h59: sinewave <= 12'h67B;
        8'h5A: sinewave <= 12'h65D;
        8'h5B: sinewave <= 12'h63E;
        8'h5C: sinewave <= 12'h61E;
        8'h5D: sinewave <= 12'h5FD;
        8'h5E: sinewave <= 12'h5DB;
        8'h5F: sinewave <= 12'h5B9;
        8'h60: sinewave <= 12'h595;
        8'h61: sinewave <= 12'h571;
        8'h62: sinewave <= 12'h54B;
        8'h63: sinewave <= 12'h525;
        8'h64: sinewave <= 12'h4FF;
        8'h65: sinewave <= 12'h4D7;
        8'h66: sinewave <= 12'h4AF;
        8'h67: sinewave <= 12'h486;
        8'h68: sinewave <= 12'h45C;
        8'h69: sinewave <= 12'h431;
        8'h6A: sinewave <= 12'h406;
        8'h6B: sinewave <= 12'h3DB;
        8'h6C: sinewave <= 12'h3AE;
        8'h6D: sinewave <= 12'h381;
        8'h6E: sinewave <= 12'h354;
        8'h6F: sinewave <= 12'h326;
        8'h70: sinewave <= 12'h2F8;
        8'h71: sinewave <= 12'h2C9;
        8'h72: sinewave <= 12'h299;
        8'h73: sinewave <= 12'h26A;
        8'h74: sinewave <= 12'h23A;
        8'h75: sinewave <= 12'h209;
        8'h76: sinewave <= 12'h1D8;
        8'h77: sinewave <= 12'h1A7;
        8'h78: sinewave <= 12'h176;
        8'h79: sinewave <= 12'h145;
        8'h7A: sinewave <= 12'h113;
        8'h7B: sinewave <= 12'h0E1;
        8'h7C: sinewave <= 12'h0AF;
        8'h7D: sinewave <= 12'h07D;
        8'h7E: sinewave <= 12'h04B;
        8'h7F: sinewave <= 12'h019;
        8'h80: sinewave <= 12'hFE7;
        8'h81: sinewave <= 12'hFB5;
        8'h82: sinewave <= 12'hF83;
        8'h83: sinewave <= 12'hF51;
        8'h84: sinewave <= 12'hF1F;
        8'h85: sinewave <= 12'hEED;
        8'h86: sinewave <= 12'hEBB;
        8'h87: sinewave <= 12'hE8A;
        8'h88: sinewave <= 12'hE59;
        8'h89: sinewave <= 12'hE28;
        8'h8A: sinewave <= 12'hDF7;
        8'h8B: sinewave <= 12'hDC6;
        8'h8C: sinewave <= 12'hD96;
        8'h8D: sinewave <= 12'hD67;
        8'h8E: sinewave <= 12'hD37;
        8'h8F: sinewave <= 12'hD08;
        8'h90: sinewave <= 12'hCDA;
        8'h91: sinewave <= 12'hCAC;
        8'h92: sinewave <= 12'hC7F;
        8'h93: sinewave <= 12'hC52;
        8'h94: sinewave <= 12'hC25;
        8'h95: sinewave <= 12'hBFA;
        8'h96: sinewave <= 12'hBCF;
        8'h97: sinewave <= 12'hBA4;
        8'h98: sinewave <= 12'hB7A;
        8'h99: sinewave <= 12'hB51;
        8'h9A: sinewave <= 12'hB29;
        8'h9B: sinewave <= 12'hB01;
        8'h9C: sinewave <= 12'hADB;
        8'h9D: sinewave <= 12'hAB5;
        8'h9E: sinewave <= 12'hA8F;
        8'h9F: sinewave <= 12'hA6B;
        8'hA0: sinewave <= 12'hA47;
        8'hA1: sinewave <= 12'hA25;
        8'hA2: sinewave <= 12'hA03;
        8'hA3: sinewave <= 12'h9E2;
        8'hA4: sinewave <= 12'h9C2;
        8'hA5: sinewave <= 12'h9A3;
        8'hA6: sinewave <= 12'h985;
        8'hA7: sinewave <= 12'h969;
        8'hA8: sinewave <= 12'h94D;
        8'hA9: sinewave <= 12'h932;
        8'hAA: sinewave <= 12'h918;
        8'hAB: sinewave <= 12'h8FF;
        8'hAC: sinewave <= 12'h8E8;
        8'hAD: sinewave <= 12'h8D1;
        8'hAE: sinewave <= 12'h8BB;
        8'hAF: sinewave <= 12'h8A7;
        8'hB0: sinewave <= 12'h894;
        8'hB1: sinewave <= 12'h882;
        8'hB2: sinewave <= 12'h871;
        8'hB3: sinewave <= 12'h861;
        8'hB4: sinewave <= 12'h852;
        8'hB5: sinewave <= 12'h845;
        8'hB6: sinewave <= 12'h839;
        8'hB7: sinewave <= 12'h82E;
        8'hB8: sinewave <= 12'h824;
        8'hB9: sinewave <= 12'h81B;
        8'hBA: sinewave <= 12'h814;
        8'hBB: sinewave <= 12'h80E;
        8'hBC: sinewave <= 12'h809;
        8'hBD: sinewave <= 12'h805;
        8'hBE: sinewave <= 12'h803;
        8'hBF: sinewave <= 12'h802;
        8'hC0: sinewave <= 12'h802;
        8'hC1: sinewave <= 12'h803;
        8'hC2: sinewave <= 12'h805;
        8'hC3: sinewave <= 12'h809;
        8'hC4: sinewave <= 12'h80E;
        8'hC5: sinewave <= 12'h814;
        8'hC6: sinewave <= 12'h81B;
        8'hC7: sinewave <= 12'h824;
        8'hC8: sinewave <= 12'h82E;
        8'hC9: sinewave <= 12'h839;
        8'hCA: sinewave <= 12'h845;
        8'hCB: sinewave <= 12'h852;
        8'hCC: sinewave <= 12'h861;
        8'hCD: sinewave <= 12'h871;
        8'hCE: sinewave <= 12'h882;
        8'hCF: sinewave <= 12'h894;
        8'hD0: sinewave <= 12'h8A7;
        8'hD1: sinewave <= 12'h8BB;
        8'hD2: sinewave <= 12'h8D1;
        8'hD3: sinewave <= 12'h8E8;
        8'hD4: sinewave <= 12'h8FF;
        8'hD5: sinewave <= 12'h918;
        8'hD6: sinewave <= 12'h932;
        8'hD7: sinewave <= 12'h94D;
        8'hD8: sinewave <= 12'h969;
        8'hD9: sinewave <= 12'h985;
        8'hDA: sinewave <= 12'h9A3;
        8'hDB: sinewave <= 12'h9C2;
        8'hDC: sinewave <= 12'h9E2;
        8'hDD: sinewave <= 12'hA03;
        8'hDE: sinewave <= 12'hA25;
        8'hDF: sinewave <= 12'hA47;
        8'hE0: sinewave <= 12'hA6B;
        8'hE1: sinewave <= 12'hA8F;
        8'hE2: sinewave <= 12'hAB5;
        8'hE3: sinewave <= 12'hADB;
        8'hE4: sinewave <= 12'hB01;
        8'hE5: sinewave <= 12'hB29;
        8'hE6: sinewave <= 12'hB51;
        8'hE7: sinewave <= 12'hB7A;
        8'hE8: sinewave <= 12'hBA4;
        8'hE9: sinewave <= 12'hBCF;
        8'hEA: sinewave <= 12'hBFA;
        8'hEB: sinewave <= 12'hC25;
        8'hEC: sinewave <= 12'hC52;
        8'hED: sinewave <= 12'hC7F;
        8'hEE: sinewave <= 12'hCAC;
        8'hEF: sinewave <= 12'hCDA;
        8'hF0: sinewave <= 12'hD08;
        8'hF1: sinewave <= 12'hD37;
        8'hF2: sinewave <= 12'hD67;
        8'hF3: sinewave <= 12'hD96;
        8'hF4: sinewave <= 12'hDC6;
        8'hF5: sinewave <= 12'hDF7;
        8'hF6: sinewave <= 12'hE28;
        8'hF7: sinewave <= 12'hE59;
        8'hF8: sinewave <= 12'hE8A;
        8'hF9: sinewave <= 12'hEBB;
        8'hFA: sinewave <= 12'hEED;
        8'hFB: sinewave <= 12'hF1F;
        8'hFC: sinewave <= 12'hF51;
        8'hFD: sinewave <= 12'hF83;
        8'hFE: sinewave <= 12'hFB5;
        8'hFF: sinewave <= 12'hFE7;
        endcase
    end
end

initial begin
	$dumpfile("simpleSine_waves.vcd");
	$dumpvars;
end

endmodule